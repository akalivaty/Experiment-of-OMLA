//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 1 0 1 1 1 0 0 1 1 1 1 1 1 1 1 1 0 0 1 1 1 1 0 0 0 1 0 0 0 0 0 1 1 1 0 0 1 1 1 1 0 0 0 0 1 0 1 1 0 1 1 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:39 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1230,
    new_n1231, new_n1232, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(new_n204));
  XOR2_X1   g0004(.A(new_n204), .B(KEYINPUT64), .Z(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n211), .A2(G20), .ZN(new_n212));
  INV_X1    g0012(.A(G58), .ZN(new_n213));
  INV_X1    g0013(.A(G68), .ZN(new_n214));
  NAND3_X1  g0014(.A1(new_n213), .A2(new_n214), .A3(KEYINPUT65), .ZN(new_n215));
  INV_X1    g0015(.A(KEYINPUT65), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n216), .B1(G58), .B2(G68), .ZN(new_n217));
  NAND3_X1  g0017(.A1(new_n215), .A2(new_n217), .A3(G50), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT67), .Z(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n222));
  NAND3_X1  g0022(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT66), .Z(new_n225));
  OAI21_X1  g0025(.A(new_n206), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n209), .B1(new_n212), .B2(new_n218), .C1(new_n226), .C2(KEYINPUT1), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XOR2_X1   g0028(.A(G238), .B(G244), .Z(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT68), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT69), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n233), .B(new_n237), .Z(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT70), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G351));
  XNOR2_X1  g0046(.A(KEYINPUT3), .B(G33), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n247), .A2(G232), .A3(G1698), .ZN(new_n248));
  INV_X1    g0048(.A(G1698), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n247), .A2(G226), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G33), .A2(G97), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n248), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G33), .A2(G41), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n211), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT72), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n253), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(KEYINPUT72), .A2(G33), .A3(G41), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n258), .A2(new_n211), .A3(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G1), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n261), .B1(G41), .B2(G45), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT71), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n261), .B(KEYINPUT71), .C1(G41), .C2(G45), .ZN(new_n265));
  NAND4_X1  g0065(.A1(new_n260), .A2(new_n264), .A3(G274), .A4(new_n265), .ZN(new_n266));
  AND2_X1   g0066(.A1(new_n260), .A2(new_n262), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G238), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n256), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT13), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT13), .ZN(new_n271));
  NAND4_X1  g0071(.A1(new_n256), .A2(new_n271), .A3(new_n266), .A4(new_n268), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n270), .A2(KEYINPUT78), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT78), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n269), .A2(new_n274), .A3(KEYINPUT13), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n273), .A2(G169), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(KEYINPUT14), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT14), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n273), .A2(new_n278), .A3(G169), .A4(new_n275), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n270), .A2(G179), .A3(new_n272), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT80), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  OR2_X1    g0082(.A1(new_n280), .A2(new_n281), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n277), .A2(new_n279), .A3(new_n282), .A4(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G33), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n210), .B1(new_n206), .B2(new_n285), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n285), .A2(G20), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G20), .ZN(new_n289));
  OAI22_X1  g0089(.A1(new_n288), .A2(new_n202), .B1(new_n289), .B2(G68), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n285), .ZN(new_n291));
  INV_X1    g0091(.A(G50), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n286), .B1(new_n290), .B2(new_n293), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n294), .B(KEYINPUT11), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n261), .A2(G13), .A3(G20), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(KEYINPUT73), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT73), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n298), .A2(new_n261), .A3(G13), .A4(G20), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n261), .A2(G20), .ZN(new_n301));
  INV_X1    g0101(.A(new_n286), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G68), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n297), .A2(new_n299), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(new_n214), .ZN(new_n307));
  XNOR2_X1  g0107(.A(new_n307), .B(KEYINPUT12), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n295), .A2(new_n305), .A3(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT79), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n309), .B(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n284), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G190), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n270), .A2(new_n272), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n273), .A2(new_n275), .ZN(new_n316));
  INV_X1    g0116(.A(G200), .ZN(new_n317));
  OAI221_X1 g0117(.A(new_n311), .B1(new_n314), .B2(new_n315), .C1(new_n316), .C2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n313), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n247), .A2(G222), .A3(new_n249), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n247), .A2(G223), .A3(G1698), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n320), .B(new_n321), .C1(new_n202), .C2(new_n247), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n255), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n267), .A2(G226), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n323), .A2(new_n266), .A3(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G169), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g0127(.A(KEYINPUT8), .B(G58), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n328), .A2(new_n288), .ZN(new_n329));
  INV_X1    g0129(.A(G150), .ZN(new_n330));
  OAI22_X1  g0130(.A1(new_n201), .A2(new_n289), .B1(new_n291), .B2(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n286), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n306), .A2(new_n292), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n300), .A2(G50), .A3(new_n302), .A4(new_n301), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n327), .B(new_n335), .C1(G179), .C2(new_n325), .ZN(new_n336));
  AND2_X1   g0136(.A1(new_n322), .A2(new_n255), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n324), .A2(new_n266), .ZN(new_n338));
  OAI21_X1  g0138(.A(G200), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT9), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n335), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n323), .A2(G190), .A3(new_n266), .A4(new_n324), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n332), .A2(new_n333), .A3(new_n334), .A4(KEYINPUT9), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NOR3_X1   g0145(.A1(new_n342), .A2(KEYINPUT10), .A3(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT10), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n343), .A2(new_n344), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n325), .A2(G200), .B1(new_n340), .B2(new_n335), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n336), .B1(new_n346), .B2(new_n350), .ZN(new_n351));
  XOR2_X1   g0151(.A(KEYINPUT8), .B(G58), .Z(new_n352));
  NOR2_X1   g0152(.A1(G20), .A2(G33), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(KEYINPUT75), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT75), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n291), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n352), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n357), .B1(new_n289), .B2(new_n202), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT76), .ZN(new_n359));
  XNOR2_X1  g0159(.A(KEYINPUT15), .B(G87), .ZN(new_n360));
  OAI22_X1  g0160(.A1(new_n358), .A2(new_n359), .B1(new_n288), .B2(new_n360), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n358), .A2(new_n359), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n286), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n300), .A2(G77), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n364), .B1(new_n304), .B2(G77), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n267), .A2(G244), .ZN(new_n367));
  AND2_X1   g0167(.A1(new_n367), .A2(new_n266), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n247), .A2(G232), .A3(new_n249), .ZN(new_n369));
  INV_X1    g0169(.A(G107), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n247), .A2(G1698), .ZN(new_n371));
  INV_X1    g0171(.A(G238), .ZN(new_n372));
  OAI221_X1 g0172(.A(new_n369), .B1(new_n370), .B2(new_n247), .C1(new_n371), .C2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n255), .ZN(new_n374));
  AND2_X1   g0174(.A1(new_n368), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(G179), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(G169), .B1(new_n368), .B2(new_n374), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n366), .A2(new_n377), .A3(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n368), .A2(G190), .A3(new_n374), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(KEYINPUT74), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT74), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n368), .A2(new_n374), .A3(new_n383), .A4(G190), .ZN(new_n384));
  AND2_X1   g0184(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n368), .A2(new_n374), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(G200), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n387), .A2(new_n363), .A3(new_n365), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n380), .B1(new_n385), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(KEYINPUT77), .B1(new_n351), .B2(new_n389), .ZN(new_n390));
  AND3_X1   g0190(.A1(new_n387), .A2(new_n363), .A3(new_n365), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n382), .A2(new_n384), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n378), .B1(new_n376), .B2(new_n375), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n391), .A2(new_n392), .B1(new_n393), .B2(new_n366), .ZN(new_n394));
  OAI21_X1  g0194(.A(KEYINPUT10), .B1(new_n342), .B2(new_n345), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n348), .A2(new_n349), .A3(new_n347), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT77), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n394), .A2(new_n397), .A3(new_n398), .A4(new_n336), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n390), .A2(new_n399), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n306), .A2(new_n352), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n401), .B1(new_n303), .B2(new_n352), .ZN(new_n402));
  XNOR2_X1  g0202(.A(G58), .B(G68), .ZN(new_n403));
  AOI22_X1  g0203(.A1(new_n403), .A2(G20), .B1(G159), .B2(new_n353), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT7), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT3), .ZN(new_n406));
  NOR3_X1   g0206(.A1(new_n406), .A2(KEYINPUT81), .A3(G33), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n407), .B1(new_n247), .B2(KEYINPUT81), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n405), .B1(new_n408), .B2(new_n289), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n285), .A2(KEYINPUT3), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n406), .A2(G33), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n410), .A2(new_n411), .A3(KEYINPUT81), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT81), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n413), .A2(new_n285), .A3(KEYINPUT3), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n412), .A2(new_n405), .A3(new_n289), .A4(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(G68), .ZN(new_n416));
  OAI211_X1 g0216(.A(KEYINPUT16), .B(new_n404), .C1(new_n409), .C2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT82), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n412), .A2(new_n414), .ZN(new_n419));
  OAI21_X1  g0219(.A(KEYINPUT7), .B1(new_n419), .B2(G20), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n420), .A2(G68), .A3(new_n415), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT82), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n421), .A2(new_n422), .A3(KEYINPUT16), .A4(new_n404), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n418), .A2(new_n423), .ZN(new_n424));
  OR2_X1    g0224(.A1(new_n405), .A2(KEYINPUT83), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n405), .A2(KEYINPUT83), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n425), .B(new_n426), .C1(new_n247), .C2(G20), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n410), .A2(new_n411), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n428), .A2(KEYINPUT83), .A3(new_n405), .A4(new_n289), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n427), .A2(new_n429), .A3(G68), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n404), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT16), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n286), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n402), .B1(new_n424), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n260), .A2(G232), .A3(new_n262), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n266), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(G226), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(G1698), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n441), .B1(G223), .B2(G1698), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n442), .B1(new_n414), .B2(new_n412), .ZN(new_n443));
  INV_X1    g0243(.A(G87), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n285), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n255), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n439), .A2(new_n446), .A3(G190), .ZN(new_n447));
  OAI22_X1  g0247(.A1(new_n408), .A2(new_n442), .B1(new_n285), .B2(new_n444), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n438), .B1(new_n255), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n447), .B1(new_n449), .B2(new_n317), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n436), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT17), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n449), .A2(G179), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n439), .A2(new_n446), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(G169), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  OAI21_X1  g0259(.A(KEYINPUT18), .B1(new_n436), .B2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT18), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n434), .B1(new_n423), .B2(new_n418), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n458), .B(new_n461), .C1(new_n462), .C2(new_n402), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n436), .A2(KEYINPUT17), .A3(new_n451), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n454), .A2(new_n460), .A3(new_n463), .A4(new_n464), .ZN(new_n465));
  NOR3_X1   g0265(.A1(new_n319), .A2(new_n400), .A3(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n360), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n300), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n419), .A2(new_n289), .A3(G68), .ZN(new_n469));
  AOI21_X1  g0269(.A(KEYINPUT19), .B1(new_n287), .B2(G97), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT19), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n289), .B1(new_n251), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(G97), .A2(G107), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n444), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n470), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n302), .B1(new_n469), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n261), .A2(G33), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n300), .A2(new_n302), .A3(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  AOI211_X1 g0279(.A(new_n468), .B(new_n476), .C1(new_n467), .C2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(G45), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n260), .B(G250), .C1(G1), .C2(new_n481), .ZN(new_n482));
  OR2_X1    g0282(.A1(new_n482), .A2(KEYINPUT85), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(KEYINPUT85), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n481), .A2(G1), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n483), .A2(new_n484), .B1(G274), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(G116), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n285), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(G244), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n489), .B1(new_n412), .B2(new_n414), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n488), .B1(new_n490), .B2(G1698), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT87), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT86), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n249), .A2(G238), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n419), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  OAI21_X1  g0296(.A(KEYINPUT86), .B1(new_n408), .B2(new_n494), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n491), .A2(new_n492), .A3(new_n496), .A4(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n255), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n493), .B1(new_n419), .B2(new_n495), .ZN(new_n500));
  AOI211_X1 g0300(.A(KEYINPUT86), .B(new_n494), .C1(new_n412), .C2(new_n414), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n492), .B1(new_n502), .B2(new_n491), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n486), .B1(new_n499), .B2(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n480), .B1(new_n504), .B2(new_n326), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n376), .B(new_n486), .C1(new_n499), .C2(new_n503), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT88), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n491), .A2(new_n496), .A3(new_n497), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT87), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n510), .A2(new_n255), .A3(new_n498), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n511), .A2(KEYINPUT88), .A3(new_n376), .A4(new_n486), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n505), .A2(new_n508), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n504), .A2(G200), .ZN(new_n514));
  OAI211_X1 g0314(.A(G190), .B(new_n486), .C1(new_n499), .C2(new_n503), .ZN(new_n515));
  AOI211_X1 g0315(.A(new_n468), .B(new_n476), .C1(G87), .C2(new_n479), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(KEYINPUT4), .B1(new_n490), .B2(new_n249), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n247), .A2(KEYINPUT4), .A3(G244), .A4(new_n249), .ZN(new_n521));
  NAND2_X1  g0321(.A1(G33), .A2(G283), .ZN(new_n522));
  INV_X1    g0322(.A(G250), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n521), .B(new_n522), .C1(new_n523), .C2(new_n371), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n255), .B1(new_n520), .B2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(G274), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n210), .B1(new_n257), .B2(new_n253), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n526), .B1(new_n527), .B2(new_n259), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT84), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT5), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G41), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n529), .B1(new_n485), .B2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n485), .A2(new_n529), .A3(new_n531), .ZN(new_n534));
  INV_X1    g0334(.A(G41), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT5), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n528), .A2(new_n533), .A3(new_n534), .A4(new_n536), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n261), .B(G45), .C1(new_n535), .C2(KEYINPUT5), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n536), .B1(new_n538), .B2(KEYINPUT84), .ZN(new_n539));
  OAI211_X1 g0339(.A(G257), .B(new_n260), .C1(new_n539), .C2(new_n532), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n525), .A2(new_n541), .A3(G190), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n317), .B1(new_n525), .B2(new_n541), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n427), .A2(new_n429), .A3(G107), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT6), .ZN(new_n545));
  AND2_X1   g0345(.A1(G97), .A2(G107), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n545), .B1(new_n546), .B2(new_n473), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n370), .A2(KEYINPUT6), .A3(G97), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n549), .A2(G20), .B1(G77), .B2(new_n353), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n544), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n286), .ZN(new_n552));
  INV_X1    g0352(.A(G97), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n306), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n300), .A2(G97), .A3(new_n302), .A4(new_n477), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n552), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n543), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n556), .B1(new_n551), .B2(new_n286), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n525), .A2(new_n541), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n560), .B1(new_n561), .B2(new_n326), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n525), .A2(new_n541), .A3(new_n376), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n542), .A2(new_n559), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n306), .A2(KEYINPUT25), .A3(new_n370), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT25), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n566), .B1(new_n300), .B2(G107), .ZN(new_n567));
  AOI22_X1  g0367(.A1(G107), .A2(new_n479), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT91), .ZN(new_n569));
  NAND2_X1  g0369(.A1(KEYINPUT22), .A2(G87), .ZN(new_n570));
  AOI211_X1 g0370(.A(G20), .B(new_n570), .C1(new_n412), .C2(new_n414), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n444), .A2(G20), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n572), .A2(new_n410), .A3(new_n411), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT22), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT23), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(new_n289), .B2(G107), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n370), .A2(KEYINPUT23), .A3(G20), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n577), .A2(new_n578), .B1(new_n287), .B2(G116), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  OAI21_X1  g0380(.A(KEYINPUT24), .B1(new_n571), .B2(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(KEYINPUT22), .B1(new_n247), .B2(new_n572), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n289), .A2(G33), .A3(G116), .ZN(new_n583));
  AND3_X1   g0383(.A1(new_n370), .A2(KEYINPUT23), .A3(G20), .ZN(new_n584));
  AOI21_X1  g0384(.A(KEYINPUT23), .B1(new_n370), .B2(G20), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n570), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n419), .A2(new_n289), .A3(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT24), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n587), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n581), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n569), .B1(new_n592), .B2(new_n286), .ZN(new_n593));
  AOI211_X1 g0393(.A(KEYINPUT91), .B(new_n302), .C1(new_n581), .C2(new_n591), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n568), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  OAI211_X1 g0395(.A(G264), .B(new_n260), .C1(new_n539), .C2(new_n532), .ZN(new_n596));
  AND2_X1   g0396(.A1(new_n537), .A2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(G257), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(G1698), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n599), .B1(G250), .B2(G1698), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n600), .B1(new_n414), .B2(new_n412), .ZN(new_n601));
  INV_X1    g0401(.A(G294), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n285), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n255), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(KEYINPUT92), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT92), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n606), .B(new_n255), .C1(new_n601), .C2(new_n603), .ZN(new_n607));
  AND3_X1   g0407(.A1(new_n597), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n604), .A2(new_n537), .A3(new_n596), .ZN(new_n609));
  OAI22_X1  g0409(.A1(new_n608), .A2(new_n326), .B1(new_n376), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n595), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n597), .A2(new_n605), .A3(new_n314), .A4(new_n607), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n609), .A2(new_n317), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n614), .B(new_n568), .C1(new_n594), .C2(new_n593), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n564), .A2(new_n611), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n306), .A2(new_n487), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n300), .A2(G116), .A3(new_n302), .A4(new_n477), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n522), .B(new_n289), .C1(G33), .C2(new_n553), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n487), .A2(G20), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n286), .A2(KEYINPUT89), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(KEYINPUT89), .B1(new_n286), .B2(new_n621), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n620), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT20), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OAI211_X1 g0426(.A(KEYINPUT20), .B(new_n620), .C1(new_n622), .C2(new_n623), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n619), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n598), .A2(new_n249), .ZN(new_n629));
  INV_X1    g0429(.A(G264), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(G1698), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n632), .B1(new_n412), .B2(new_n414), .ZN(new_n633));
  INV_X1    g0433(.A(G303), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n247), .A2(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n255), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  OAI211_X1 g0436(.A(G270), .B(new_n260), .C1(new_n539), .C2(new_n532), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n636), .A2(new_n537), .A3(G179), .A4(new_n637), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n628), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n619), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n286), .A2(new_n621), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT89), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n286), .A2(KEYINPUT89), .A3(new_n621), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(KEYINPUT20), .B1(new_n645), .B2(new_n620), .ZN(new_n646));
  INV_X1    g0446(.A(new_n627), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n640), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n636), .A2(new_n537), .A3(new_n637), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(new_n649), .A3(G169), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT21), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n639), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n648), .A2(new_n649), .A3(KEYINPUT21), .A4(G169), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n649), .A2(G200), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n628), .A2(new_n654), .ZN(new_n655));
  OAI22_X1  g0455(.A1(new_n655), .A2(KEYINPUT90), .B1(new_n314), .B2(new_n649), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n655), .A2(KEYINPUT90), .ZN(new_n657));
  OAI211_X1 g0457(.A(new_n652), .B(new_n653), .C1(new_n656), .C2(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n616), .A2(new_n658), .ZN(new_n659));
  AND3_X1   g0459(.A1(new_n466), .A2(new_n519), .A3(new_n659), .ZN(G372));
  NAND2_X1  g0460(.A1(new_n562), .A2(new_n563), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n513), .A2(new_n517), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(KEYINPUT26), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n514), .A2(KEYINPUT93), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n515), .A2(new_n516), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT93), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n504), .A2(new_n667), .A3(G200), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n665), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT26), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n505), .A2(new_n506), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n669), .A2(new_n670), .A3(new_n662), .A4(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n559), .A2(new_n542), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n615), .A2(new_n661), .A3(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n611), .A2(new_n653), .A3(new_n652), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(new_n669), .A3(new_n675), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n664), .A2(new_n672), .A3(new_n676), .A4(new_n671), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n466), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n678), .B(KEYINPUT94), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n460), .A2(new_n463), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n316), .A2(new_n317), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n315), .A2(new_n314), .ZN(new_n682));
  NOR3_X1   g0482(.A1(new_n312), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n313), .B1(new_n683), .B2(new_n380), .ZN(new_n684));
  AOI21_X1  g0484(.A(KEYINPUT17), .B1(new_n436), .B2(new_n451), .ZN(new_n685));
  NOR4_X1   g0485(.A1(new_n462), .A2(new_n453), .A3(new_n402), .A4(new_n450), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n680), .B1(new_n684), .B2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n397), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n336), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  OR2_X1    g0490(.A1(new_n679), .A2(new_n690), .ZN(G369));
  NAND2_X1  g0491(.A1(new_n652), .A2(new_n653), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n261), .A2(new_n289), .A3(G13), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n693), .A2(KEYINPUT27), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(KEYINPUT27), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(G213), .A3(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(G343), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n628), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n692), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n701), .B1(new_n658), .B2(new_n700), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(G330), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n611), .A2(new_n615), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n595), .A2(new_n698), .ZN(new_n706));
  OAI22_X1  g0506(.A1(new_n705), .A2(new_n706), .B1(new_n611), .B2(new_n699), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n692), .A2(new_n699), .ZN(new_n709));
  OR2_X1    g0509(.A1(new_n709), .A2(new_n705), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n595), .A2(new_n610), .A3(new_n699), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n708), .A2(new_n713), .ZN(G399));
  INV_X1    g0514(.A(new_n207), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(G41), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n474), .A2(G116), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n717), .A2(G1), .A3(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n719), .B1(new_n218), .B2(new_n717), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n720), .B(KEYINPUT28), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT29), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n677), .A2(new_n722), .A3(new_n699), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n513), .A2(new_n517), .A3(new_n670), .A4(new_n662), .ZN(new_n724));
  AND3_X1   g0524(.A1(new_n676), .A2(new_n671), .A3(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n669), .A2(new_n662), .A3(new_n671), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(KEYINPUT26), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n698), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n723), .B1(new_n728), .B2(new_n722), .ZN(new_n729));
  NOR4_X1   g0529(.A1(new_n518), .A2(new_n616), .A3(new_n658), .A4(new_n698), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n604), .A2(new_n596), .ZN(new_n731));
  OAI211_X1 g0531(.A(new_n486), .B(new_n731), .C1(new_n499), .C2(new_n503), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(KEYINPUT95), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT95), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n511), .A2(new_n734), .A3(new_n486), .A4(new_n731), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n561), .A2(new_n638), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n733), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT30), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n561), .A2(new_n609), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT96), .ZN(new_n740));
  AND3_X1   g0540(.A1(new_n504), .A2(new_n376), .A3(new_n649), .ZN(new_n741));
  AOI22_X1  g0541(.A1(new_n737), .A2(new_n738), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n733), .A2(KEYINPUT30), .A3(new_n735), .A4(new_n736), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n699), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(KEYINPUT31), .B1(new_n730), .B2(new_n744), .ZN(new_n745));
  AND2_X1   g0545(.A1(new_n732), .A2(KEYINPUT95), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n736), .B1(new_n732), .B2(KEYINPUT95), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n738), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n740), .A2(new_n741), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n748), .A2(new_n743), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(new_n698), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT31), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n745), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n729), .B1(G330), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n721), .B1(new_n755), .B2(G1), .ZN(G364));
  INV_X1    g0556(.A(G13), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(G20), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n261), .B1(new_n758), .B2(G45), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n716), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n210), .B1(G20), .B2(new_n326), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n289), .A2(new_n314), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR3_X1   g0566(.A1(new_n766), .A2(new_n317), .A3(G179), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n289), .A2(G190), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR3_X1   g0570(.A1(new_n770), .A2(new_n376), .A3(G200), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(G311), .ZN(new_n773));
  OAI22_X1  g0573(.A1(new_n768), .A2(new_n634), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n376), .A2(new_n317), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n765), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  AOI211_X1 g0577(.A(new_n247), .B(new_n774), .C1(G326), .C2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(G179), .A2(G200), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G190), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G20), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G294), .ZN(new_n782));
  NOR3_X1   g0582(.A1(new_n770), .A2(G179), .A3(new_n317), .ZN(new_n783));
  XOR2_X1   g0583(.A(new_n783), .B(KEYINPUT97), .Z(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G283), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n775), .A2(new_n769), .ZN(new_n786));
  INV_X1    g0586(.A(G317), .ZN(new_n787));
  AND2_X1   g0587(.A1(new_n787), .A2(KEYINPUT33), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n787), .A2(KEYINPUT33), .ZN(new_n789));
  NOR3_X1   g0589(.A1(new_n786), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  NOR3_X1   g0590(.A1(new_n766), .A2(new_n376), .A3(G200), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(G322), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n769), .A2(new_n779), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n790), .B(new_n794), .C1(G329), .C2(new_n796), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n778), .A2(new_n782), .A3(new_n785), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n784), .A2(G107), .ZN(new_n799));
  INV_X1    g0599(.A(new_n781), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(new_n553), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n428), .B(new_n801), .C1(G58), .C2(new_n791), .ZN(new_n802));
  INV_X1    g0602(.A(G159), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n795), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n804), .B(KEYINPUT32), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n768), .A2(new_n444), .B1(new_n786), .B2(new_n214), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n772), .A2(new_n202), .B1(new_n292), .B2(new_n776), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n799), .A2(new_n802), .A3(new_n805), .A4(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n764), .B1(new_n798), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(G13), .A2(G33), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(G20), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(new_n763), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n419), .A2(new_n715), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n816), .B1(new_n245), .B2(G45), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(G45), .B2(new_n218), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n715), .A2(new_n428), .ZN(new_n819));
  AOI22_X1  g0619(.A1(G355), .A2(new_n819), .B1(new_n487), .B2(new_n715), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n762), .B(new_n810), .C1(new_n814), .C2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n813), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n822), .B1(new_n702), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n703), .A2(new_n762), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n702), .A2(G330), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n824), .B1(new_n825), .B2(new_n826), .ZN(G396));
  NOR2_X1   g0627(.A1(new_n380), .A2(new_n698), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n366), .A2(new_n698), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(new_n385), .B2(new_n388), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n828), .B1(new_n830), .B2(new_n380), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n677), .A2(new_n699), .A3(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n833), .A2(KEYINPUT99), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n831), .B1(new_n677), .B2(new_n699), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n834), .B(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n754), .A2(G330), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n761), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n837), .B2(new_n836), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n763), .A2(new_n811), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n761), .B1(G77), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(G283), .ZN(new_n843));
  OAI22_X1  g0643(.A1(new_n792), .A2(new_n602), .B1(new_n786), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(G107), .B2(new_n767), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n784), .A2(G87), .ZN(new_n846));
  INV_X1    g0646(.A(new_n801), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n776), .A2(new_n634), .B1(new_n795), .B2(new_n773), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n247), .B(new_n848), .C1(G116), .C2(new_n771), .ZN(new_n849));
  NAND4_X1  g0649(.A1(new_n845), .A2(new_n846), .A3(new_n847), .A4(new_n849), .ZN(new_n850));
  AOI22_X1  g0650(.A1(G143), .A2(new_n791), .B1(new_n771), .B2(G159), .ZN(new_n851));
  INV_X1    g0651(.A(new_n786), .ZN(new_n852));
  AOI22_X1  g0652(.A1(G137), .A2(new_n777), .B1(new_n852), .B2(G150), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  XOR2_X1   g0654(.A(new_n854), .B(KEYINPUT34), .Z(new_n855));
  NAND2_X1  g0655(.A1(new_n784), .A2(G68), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n781), .A2(G58), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n767), .A2(G50), .B1(G132), .B2(new_n796), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n856), .A2(new_n419), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n850), .B1(new_n855), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n842), .B1(new_n860), .B2(new_n763), .ZN(new_n861));
  XOR2_X1   g0661(.A(new_n861), .B(KEYINPUT98), .Z(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n812), .B2(new_n831), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n839), .A2(new_n863), .ZN(G384));
  AOI211_X1 g0664(.A(new_n487), .B(new_n212), .C1(new_n549), .C2(KEYINPUT35), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(KEYINPUT35), .B2(new_n549), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n866), .B(KEYINPUT36), .ZN(new_n867));
  OAI21_X1  g0667(.A(G77), .B1(new_n213), .B2(new_n214), .ZN(new_n868));
  OAI22_X1  g0668(.A1(new_n218), .A2(new_n868), .B1(G50), .B2(new_n214), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n869), .A2(G1), .A3(new_n757), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n871), .B(KEYINPUT100), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n284), .A2(new_n312), .A3(new_n698), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n873), .A2(KEYINPUT101), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(KEYINPUT101), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n312), .A2(new_n698), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n313), .A2(new_n318), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n874), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  AND3_X1   g0679(.A1(new_n754), .A2(new_n831), .A3(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n458), .B1(new_n462), .B2(new_n402), .ZN(new_n881));
  XOR2_X1   g0681(.A(new_n696), .B(KEYINPUT102), .Z(new_n882));
  OAI21_X1  g0682(.A(new_n882), .B1(new_n462), .B2(new_n402), .ZN(new_n883));
  XOR2_X1   g0683(.A(KEYINPUT103), .B(KEYINPUT37), .Z(new_n884));
  NAND4_X1  g0684(.A1(new_n452), .A2(new_n881), .A3(new_n883), .A4(new_n884), .ZN(new_n885));
  AOI211_X1 g0685(.A(new_n402), .B(new_n450), .C1(new_n424), .C2(new_n435), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n421), .A2(new_n404), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n302), .B1(new_n887), .B2(new_n432), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n424), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n402), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n459), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n696), .B1(new_n889), .B2(new_n890), .ZN(new_n892));
  NOR3_X1   g0692(.A1(new_n886), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT37), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n885), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n465), .A2(new_n892), .ZN(new_n896));
  AND3_X1   g0696(.A1(new_n895), .A2(new_n896), .A3(KEYINPUT38), .ZN(new_n897));
  INV_X1    g0697(.A(new_n883), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n465), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n452), .A2(new_n881), .A3(new_n883), .ZN(new_n900));
  INV_X1    g0700(.A(new_n884), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n885), .ZN(new_n903));
  AOI21_X1  g0703(.A(KEYINPUT38), .B1(new_n899), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n897), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n880), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(KEYINPUT40), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT40), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT38), .ZN(new_n910));
  INV_X1    g0710(.A(new_n892), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n889), .A2(new_n890), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n458), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n911), .A2(new_n913), .A3(new_n452), .ZN(new_n914));
  AND3_X1   g0714(.A1(new_n452), .A2(new_n881), .A3(new_n883), .ZN(new_n915));
  AOI22_X1  g0715(.A1(KEYINPUT37), .A2(new_n914), .B1(new_n915), .B2(new_n884), .ZN(new_n916));
  INV_X1    g0716(.A(new_n680), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n911), .B1(new_n917), .B2(new_n687), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n910), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n895), .A2(new_n896), .A3(KEYINPUT38), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n880), .A2(new_n909), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n908), .A2(new_n922), .ZN(new_n923));
  AND2_X1   g0723(.A1(new_n754), .A2(new_n466), .ZN(new_n924));
  AND2_X1   g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n923), .A2(new_n924), .ZN(new_n926));
  INV_X1    g0726(.A(G330), .ZN(new_n927));
  NOR3_X1   g0727(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT39), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n930), .B1(new_n897), .B2(new_n904), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n919), .A2(KEYINPUT39), .A3(new_n920), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n313), .A2(new_n698), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT104), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n933), .B(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n931), .A2(new_n932), .A3(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n828), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n832), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n938), .A2(new_n879), .A3(new_n921), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n917), .A2(new_n882), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n936), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(KEYINPUT105), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT105), .ZN(new_n943));
  NAND4_X1  g0743(.A1(new_n936), .A2(new_n939), .A3(new_n943), .A4(new_n940), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n690), .B1(new_n729), .B2(new_n466), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n945), .B(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n929), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n947), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n949), .A2(new_n928), .B1(new_n261), .B2(new_n758), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n872), .B1(new_n948), .B2(new_n950), .ZN(G367));
  NOR2_X1   g0751(.A1(new_n237), .A2(new_n816), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n814), .B1(new_n207), .B2(new_n360), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n761), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n783), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n792), .A2(new_n634), .B1(new_n955), .B2(new_n553), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n772), .A2(new_n843), .B1(new_n602), .B2(new_n786), .ZN(new_n957));
  OAI221_X1 g0757(.A(new_n408), .B1(new_n773), .B2(new_n776), .C1(new_n787), .C2(new_n795), .ZN(new_n958));
  NOR3_X1   g0758(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n768), .A2(new_n487), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n960), .A2(KEYINPUT46), .B1(G107), .B2(new_n781), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n959), .B(new_n961), .C1(KEYINPUT46), .C2(new_n960), .ZN(new_n962));
  XNOR2_X1  g0762(.A(KEYINPUT110), .B(G137), .ZN(new_n963));
  OAI22_X1  g0763(.A1(new_n955), .A2(new_n202), .B1(new_n795), .B2(new_n963), .ZN(new_n964));
  AOI211_X1 g0764(.A(new_n428), .B(new_n964), .C1(G58), .C2(new_n767), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n781), .A2(G68), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n792), .B2(new_n330), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(KEYINPUT109), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n772), .A2(new_n292), .B1(new_n803), .B2(new_n786), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(G143), .B2(new_n777), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n965), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n967), .A2(KEYINPUT109), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n962), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT47), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n954), .B1(new_n974), .B2(new_n763), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n516), .A2(new_n699), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n669), .A2(new_n671), .A3(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n671), .B2(new_n976), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n975), .B1(new_n978), .B2(new_n823), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n564), .B1(new_n560), .B2(new_n699), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n662), .A2(new_n698), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n713), .A2(new_n982), .ZN(new_n983));
  XOR2_X1   g0783(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n984));
  XNOR2_X1  g0784(.A(new_n983), .B(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n982), .ZN(new_n986));
  AOI21_X1  g0786(.A(KEYINPUT44), .B1(new_n712), .B2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT108), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n712), .A2(KEYINPUT44), .A3(new_n986), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n987), .A2(new_n988), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n985), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n993), .B(new_n708), .Z(new_n994));
  INV_X1    g0794(.A(new_n709), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n710), .B1(new_n707), .B2(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n704), .B(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n755), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n755), .B1(new_n994), .B2(new_n998), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n716), .B(KEYINPUT41), .Z(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n760), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n986), .A2(new_n710), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT42), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n661), .B1(new_n980), .B2(new_n611), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(new_n699), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(KEYINPUT43), .B1(new_n978), .B2(KEYINPUT106), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1008), .B1(KEYINPUT106), .B2(new_n978), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n978), .A2(KEYINPUT43), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1007), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n1009), .B2(new_n1007), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n708), .A2(new_n986), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1012), .B(new_n1013), .Z(new_n1014));
  OAI21_X1  g0814(.A(new_n979), .B1(new_n1002), .B2(new_n1014), .ZN(G387));
  AOI21_X1  g0815(.A(new_n816), .B1(new_n233), .B2(G45), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n328), .A2(G50), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT50), .Z(new_n1018));
  OAI21_X1  g0818(.A(new_n481), .B1(new_n214), .B2(new_n202), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(new_n718), .B2(KEYINPUT111), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(KEYINPUT111), .B2(new_n718), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1016), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n718), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n1023), .A2(new_n819), .B1(new_n370), .B2(new_n715), .ZN(new_n1024));
  AOI211_X1 g0824(.A(new_n813), .B(new_n763), .C1(new_n1022), .C2(new_n1024), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n783), .A2(G116), .B1(G326), .B2(new_n796), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n792), .A2(new_n787), .B1(new_n772), .B2(new_n634), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n776), .A2(new_n793), .B1(new_n786), .B2(new_n773), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n767), .A2(G294), .B1(G283), .B2(new_n781), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n1029), .A2(KEYINPUT48), .B1(new_n1030), .B2(KEYINPUT113), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n1030), .A2(KEYINPUT113), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1031), .B(new_n1032), .C1(KEYINPUT48), .C2(new_n1029), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT49), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n408), .B(new_n1026), .C1(new_n1033), .C2(new_n1034), .ZN(new_n1035));
  AND2_X1   g0835(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n768), .A2(new_n202), .B1(new_n795), .B2(new_n330), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n408), .B(new_n1037), .C1(new_n784), .C2(G97), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT112), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n791), .A2(G50), .B1(new_n352), .B2(new_n852), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n771), .A2(G68), .B1(new_n777), .B2(G159), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1040), .B(new_n1041), .C1(new_n360), .C2(new_n800), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n1035), .A2(new_n1036), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT114), .ZN(new_n1044));
  OR2_X1    g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n764), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n762), .B(new_n1025), .C1(new_n1045), .C2(new_n1046), .ZN(new_n1047));
  OR2_X1    g0847(.A1(new_n707), .A2(new_n823), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n997), .A2(new_n760), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n998), .A2(KEYINPUT115), .A3(new_n716), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n755), .B2(new_n997), .ZN(new_n1051));
  AOI21_X1  g0851(.A(KEYINPUT115), .B1(new_n998), .B2(new_n716), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1049), .B1(new_n1051), .B2(new_n1052), .ZN(G393));
  OAI221_X1 g0853(.A(new_n814), .B1(new_n553), .B2(new_n207), .C1(new_n242), .C2(new_n816), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT116), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n762), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n1055), .B2(new_n1054), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n772), .A2(new_n602), .B1(new_n634), .B2(new_n786), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(G116), .B2(new_n781), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT118), .Z(new_n1060));
  AOI22_X1  g0860(.A1(new_n791), .A2(G311), .B1(new_n777), .B2(G317), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT52), .Z(new_n1062));
  OAI21_X1  g0862(.A(new_n428), .B1(new_n795), .B2(new_n793), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(new_n767), .B2(G283), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n1060), .A2(new_n799), .A3(new_n1062), .A4(new_n1064), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n791), .A2(G159), .B1(new_n777), .B2(G150), .ZN(new_n1066));
  XOR2_X1   g0866(.A(new_n1066), .B(KEYINPUT51), .Z(new_n1067));
  OAI22_X1  g0867(.A1(new_n772), .A2(new_n328), .B1(new_n292), .B2(new_n786), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n784), .A2(G87), .B1(KEYINPUT117), .B2(new_n1068), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n1068), .A2(KEYINPUT117), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n767), .A2(G68), .B1(G143), .B2(new_n796), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n781), .A2(G77), .ZN(new_n1072));
  AND3_X1   g0872(.A1(new_n1071), .A2(new_n419), .A3(new_n1072), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1067), .A2(new_n1069), .A3(new_n1070), .A4(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1065), .A2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1057), .B1(new_n1075), .B2(new_n763), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n982), .B2(new_n823), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(new_n994), .B2(new_n759), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n994), .A2(new_n998), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1079), .A2(new_n717), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n994), .A2(new_n998), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1078), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(G390));
  INV_X1    g0883(.A(new_n932), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n904), .ZN(new_n1085));
  AOI21_X1  g0885(.A(KEYINPUT39), .B1(new_n1085), .B2(new_n920), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n811), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n772), .A2(new_n553), .B1(new_n843), .B2(new_n776), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n247), .B(new_n1088), .C1(G87), .C2(new_n767), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n792), .A2(new_n487), .B1(new_n795), .B2(new_n602), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(G107), .B2(new_n852), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n1089), .A2(new_n856), .A3(new_n1072), .A4(new_n1091), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n791), .A2(G132), .B1(new_n777), .B2(G128), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT121), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n767), .A2(G150), .ZN(new_n1095));
  XOR2_X1   g0895(.A(new_n1095), .B(KEYINPUT53), .Z(new_n1096));
  INV_X1    g0896(.A(G125), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n786), .A2(new_n963), .B1(new_n795), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(G50), .B2(new_n783), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(KEYINPUT54), .B(G143), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n247), .B1(new_n772), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(G159), .B2(new_n781), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1096), .A2(new_n1099), .A3(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1092), .B1(new_n1094), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT122), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n764), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1106), .B1(new_n1105), .B2(new_n1104), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n762), .B1(new_n328), .B2(new_n840), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1087), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n754), .A2(G330), .A3(new_n831), .A4(new_n879), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n938), .A2(new_n879), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n935), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n1112), .A2(new_n1113), .B1(new_n931), .B2(new_n932), .ZN(new_n1114));
  OR2_X1    g0914(.A1(new_n873), .A2(KEYINPUT101), .ZN(new_n1115));
  AND3_X1   g0915(.A1(new_n313), .A2(new_n318), .A3(new_n877), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1115), .B1(new_n1116), .B2(new_n875), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n830), .A2(new_n380), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n727), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n676), .A2(new_n671), .A3(new_n724), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n699), .B(new_n1118), .C1(new_n1119), .C2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1117), .B1(new_n1121), .B2(new_n937), .ZN(new_n1122));
  NOR3_X1   g0922(.A1(new_n1122), .A2(new_n905), .A3(new_n935), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1111), .B1(new_n1114), .B2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1117), .B1(new_n937), .B2(new_n832), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n1125), .A2(new_n935), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n828), .B1(new_n728), .B2(new_n1118), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n906), .B(new_n1113), .C1(new_n1127), .C2(new_n1117), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1126), .A2(new_n1128), .A3(new_n1110), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1124), .A2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1109), .B1(new_n1130), .B2(new_n759), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n659), .A2(new_n519), .A3(new_n699), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n752), .B1(new_n1132), .B2(new_n751), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n744), .A2(KEYINPUT31), .ZN(new_n1134));
  OAI211_X1 g0934(.A(G330), .B(new_n831), .C1(new_n1133), .C2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n1117), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n1110), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n938), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1136), .A2(new_n1110), .A3(new_n1127), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  OAI211_X1 g0940(.A(G330), .B(new_n466), .C1(new_n1133), .C2(new_n1134), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(KEYINPUT119), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT119), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n754), .A2(new_n1143), .A3(G330), .A4(new_n466), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n946), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(KEYINPUT120), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT120), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1145), .A2(new_n946), .A3(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1140), .A2(new_n1147), .A3(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n717), .B1(new_n1150), .B2(new_n1130), .ZN(new_n1151));
  AND3_X1   g0951(.A1(new_n1145), .A2(new_n946), .A3(new_n1148), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1148), .B1(new_n1145), .B2(new_n946), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1154), .A2(new_n1124), .A3(new_n1129), .A4(new_n1140), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1131), .B1(new_n1151), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(G378));
  AOI21_X1  g0957(.A(new_n927), .B1(new_n908), .B2(new_n922), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n351), .B(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n696), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n335), .A2(new_n1162), .ZN(new_n1163));
  XOR2_X1   g0963(.A(new_n1163), .B(KEYINPUT123), .Z(new_n1164));
  XOR2_X1   g0964(.A(new_n1161), .B(new_n1164), .Z(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  AND3_X1   g0966(.A1(new_n942), .A2(new_n944), .A3(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1166), .B1(new_n942), .B2(new_n944), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1159), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n945), .A2(new_n1165), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n942), .A2(new_n944), .A3(new_n1166), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1170), .A2(new_n1158), .A3(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1169), .A2(new_n1172), .A3(new_n760), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n762), .B1(new_n292), .B2(new_n840), .ZN(new_n1174));
  INV_X1    g0974(.A(G132), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n776), .A2(new_n1097), .B1(new_n786), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n771), .A2(G137), .ZN(new_n1177));
  INV_X1    g0977(.A(G128), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n1177), .B1(new_n768), .B2(new_n1100), .C1(new_n1178), .C2(new_n792), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n1176), .B(new_n1179), .C1(G150), .C2(new_n781), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  OR2_X1    g0981(.A1(new_n1181), .A2(KEYINPUT59), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(KEYINPUT59), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n783), .A2(G159), .ZN(new_n1184));
  AOI211_X1 g0984(.A(G33), .B(G41), .C1(new_n796), .C2(G124), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .A4(new_n1185), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(G77), .A2(new_n767), .B1(new_n771), .B2(new_n467), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(G107), .A2(new_n791), .B1(new_n783), .B2(G58), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1187), .A2(new_n1188), .A3(new_n966), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n408), .A2(new_n535), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(G97), .A2(new_n852), .B1(new_n796), .B2(G283), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(new_n487), .B2(new_n776), .ZN(new_n1192));
  NOR3_X1   g0992(.A1(new_n1189), .A2(new_n1190), .A3(new_n1192), .ZN(new_n1193));
  OR2_X1    g0993(.A1(new_n1193), .A2(KEYINPUT58), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(KEYINPUT58), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1190), .B(new_n292), .C1(G33), .C2(G41), .ZN(new_n1196));
  AND4_X1   g0996(.A1(new_n1186), .A2(new_n1194), .A3(new_n1195), .A4(new_n1196), .ZN(new_n1197));
  OAI221_X1 g0997(.A(new_n1174), .B1(new_n764), .B2(new_n1197), .C1(new_n1166), .C2(new_n812), .ZN(new_n1198));
  AND2_X1   g0998(.A1(new_n1173), .A2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1140), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1154), .B1(new_n1130), .B2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1169), .A2(new_n1172), .A3(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT57), .ZN(new_n1203));
  AND2_X1   g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1169), .A2(new_n1172), .A3(new_n1201), .A4(KEYINPUT57), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(new_n716), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1199), .B1(new_n1204), .B2(new_n1206), .ZN(G375));
  OAI21_X1  g1007(.A(new_n428), .B1(new_n776), .B2(new_n602), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n772), .A2(new_n370), .B1(new_n487), .B2(new_n786), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n1208), .B(new_n1209), .C1(new_n467), .C2(new_n781), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n767), .A2(G97), .B1(G303), .B2(new_n796), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1211), .B1(new_n843), .B2(new_n792), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(G77), .B2(new_n784), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n419), .B1(new_n1175), .B2(new_n776), .C1(new_n955), .C2(new_n213), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n768), .A2(new_n803), .B1(new_n795), .B2(new_n1178), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n792), .A2(new_n963), .B1(new_n786), .B2(new_n1100), .ZN(new_n1216));
  NOR3_X1   g1016(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n771), .A2(G150), .B1(G50), .B2(new_n781), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1218), .B(KEYINPUT124), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n1210), .A2(new_n1213), .B1(new_n1217), .B2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT125), .ZN(new_n1221));
  AND2_X1   g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n763), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n761), .B1(G68), .B2(new_n841), .C1(new_n1222), .C2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(new_n1117), .B2(new_n811), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(new_n1140), .B2(new_n760), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1150), .A2(new_n1001), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1140), .B1(new_n1149), .B2(new_n1147), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1226), .B1(new_n1227), .B2(new_n1228), .ZN(G381));
  OR2_X1    g1029(.A1(G393), .A2(G396), .ZN(new_n1230));
  OR4_X1    g1030(.A1(G384), .A2(G390), .A3(G387), .A4(new_n1230), .ZN(new_n1231));
  OR2_X1    g1031(.A1(G375), .A2(G378), .ZN(new_n1232));
  OR3_X1    g1032(.A1(new_n1231), .A2(G381), .A3(new_n1232), .ZN(G407));
  OAI211_X1 g1033(.A(G407), .B(G213), .C1(G343), .C2(new_n1232), .ZN(G409));
  NAND2_X1  g1034(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1235));
  AOI21_X1  g1035(.A(KEYINPUT60), .B1(new_n1235), .B2(new_n1200), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1150), .ZN(new_n1237));
  OAI21_X1  g1037(.A(KEYINPUT126), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT126), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1239), .B(new_n1150), .C1(new_n1228), .C2(KEYINPUT60), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n717), .B1(new_n1228), .B2(KEYINPUT60), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1238), .A2(new_n1240), .A3(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(new_n1226), .ZN(new_n1243));
  INV_X1    g1043(.A(G384), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1242), .A2(G384), .A3(new_n1226), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n697), .A2(G213), .A3(G2897), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(G375), .A2(G378), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1169), .A2(new_n1172), .A3(new_n1201), .A4(new_n1001), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1156), .A2(new_n1251), .A3(new_n1173), .A4(new_n1198), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n697), .A2(G213), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n1247), .A2(new_n1249), .B1(new_n1250), .B2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT127), .ZN(new_n1257));
  AND3_X1   g1057(.A1(new_n1242), .A2(G384), .A3(new_n1226), .ZN(new_n1258));
  AOI21_X1  g1058(.A(G384), .B1(new_n1242), .B2(new_n1226), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1257), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1245), .A2(KEYINPUT127), .A3(new_n1246), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1260), .A2(new_n1261), .A3(new_n1248), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1256), .A2(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1254), .B1(G375), .B2(G378), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1264), .A2(new_n1260), .A3(new_n1261), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(KEYINPUT62), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT61), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT62), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1264), .A2(new_n1260), .A3(new_n1261), .A4(new_n1268), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1263), .A2(new_n1266), .A3(new_n1267), .A4(new_n1269), .ZN(new_n1270));
  OR2_X1    g1070(.A1(G387), .A2(new_n1082), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(G393), .A2(G396), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1230), .A2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(G387), .A2(new_n1082), .ZN(new_n1275));
  AND3_X1   g1075(.A1(new_n1271), .A2(new_n1274), .A3(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1274), .B1(new_n1271), .B2(new_n1275), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1270), .A2(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(KEYINPUT61), .B1(new_n1256), .B2(new_n1262), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT63), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1265), .A2(new_n1282), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1264), .A2(new_n1260), .A3(new_n1261), .A4(KEYINPUT63), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1281), .A2(new_n1278), .A3(new_n1283), .A4(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1280), .A2(new_n1285), .ZN(G405));
  NAND2_X1  g1086(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1287), .A2(new_n1232), .A3(new_n1250), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1232), .A2(new_n1250), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1247), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1288), .A2(new_n1291), .ZN(new_n1292));
  XNOR2_X1  g1092(.A(new_n1292), .B(new_n1278), .ZN(G402));
endmodule


