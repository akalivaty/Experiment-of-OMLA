//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 0 1 1 0 0 0 1 1 0 1 0 1 0 0 0 0 1 0 0 1 1 0 0 0 1 0 0 1 1 1 1 1 1 0 0 1 1 1 1 0 1 0 0 0 1 0 0 1 1 0 1 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:12 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n562, new_n563, new_n564, new_n565,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n624, new_n625, new_n628, new_n630, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1238, new_n1239;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  XOR2_X1   g015(.A(KEYINPUT65), .B(G120), .Z(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  XNOR2_X1  g017(.A(KEYINPUT66), .B(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G236), .A2(G238), .A3(G237), .A4(G235), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n454), .A2(new_n459), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT67), .Z(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G125), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n463), .A2(G137), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n463), .A2(KEYINPUT68), .A3(G101), .A4(G2104), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n463), .A2(G101), .A3(G2104), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT68), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n469), .A2(new_n470), .A3(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n467), .A2(new_n474), .ZN(G160));
  AND2_X1   g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  OR3_X1    g052(.A1(new_n476), .A2(new_n477), .A3(KEYINPUT69), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n464), .A2(KEYINPUT69), .ZN(new_n479));
  AOI21_X1  g054(.A(G2105), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n463), .B1(new_n478), .B2(new_n479), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  NOR2_X1   g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(new_n463), .B2(G112), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n481), .B(new_n483), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  INV_X1    g062(.A(G138), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n489), .B1(new_n476), .B2(new_n477), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT70), .ZN(new_n495));
  AND2_X1   g070(.A1(new_n495), .A2(G114), .ZN(new_n496));
  OAI21_X1  g071(.A(G2105), .B1(new_n495), .B2(G114), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n494), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n463), .A2(KEYINPUT4), .A3(G138), .ZN(new_n499));
  NAND2_X1  g074(.A1(G126), .A2(G2105), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(new_n464), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n492), .A2(new_n498), .A3(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  NAND2_X1  g079(.A1(G75), .A2(G543), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT72), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  OAI21_X1  g082(.A(KEYINPUT71), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  OAI21_X1  g083(.A(KEYINPUT5), .B1(new_n507), .B2(KEYINPUT71), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OAI211_X1 g085(.A(KEYINPUT71), .B(KEYINPUT5), .C1(new_n506), .C2(new_n507), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G62), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n505), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G651), .ZN(new_n515));
  INV_X1    g090(.A(G50), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(KEYINPUT6), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT6), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n521), .A2(new_n507), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G88), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n510), .A2(new_n511), .ZN(new_n525));
  INV_X1    g100(.A(new_n521), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OAI221_X1 g102(.A(new_n515), .B1(new_n516), .B2(new_n523), .C1(new_n524), .C2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(KEYINPUT73), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n512), .A2(new_n521), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n530), .A2(G88), .B1(G50), .B2(new_n522), .ZN(new_n531));
  AND2_X1   g106(.A1(new_n531), .A2(new_n515), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT73), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n529), .A2(new_n534), .ZN(G166));
  NAND2_X1  g110(.A1(new_n530), .A2(G89), .ZN(new_n536));
  XOR2_X1   g111(.A(KEYINPUT74), .B(KEYINPUT7), .Z(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n537), .A2(new_n538), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n539), .A2(new_n540), .B1(G51), .B2(new_n522), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n525), .A2(G63), .A3(G651), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n536), .A2(new_n541), .A3(new_n542), .ZN(G286));
  INV_X1    g118(.A(G286), .ZN(G168));
  NAND2_X1  g119(.A1(new_n522), .A2(G52), .ZN(new_n545));
  INV_X1    g120(.A(G90), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n527), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n525), .A2(G64), .ZN(new_n548));
  NAND2_X1  g123(.A1(G77), .A2(G543), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n517), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n547), .A2(new_n550), .ZN(G171));
  AOI22_X1  g126(.A1(new_n530), .A2(G81), .B1(G43), .B2(new_n522), .ZN(new_n552));
  NAND2_X1  g127(.A1(G68), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(G56), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n512), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G651), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(G860), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT75), .ZN(G153));
  NAND4_X1  g135(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT76), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND4_X1  g139(.A1(G319), .A2(G483), .A3(G661), .A4(new_n564), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT77), .ZN(G188));
  XNOR2_X1  g141(.A(KEYINPUT78), .B(KEYINPUT9), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n526), .A2(G53), .A3(G543), .A4(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT79), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(G53), .ZN(new_n571));
  NOR3_X1   g146(.A1(new_n521), .A2(new_n571), .A3(new_n507), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n572), .A2(KEYINPUT79), .A3(new_n567), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT9), .ZN(new_n574));
  OAI211_X1 g149(.A(new_n570), .B(new_n573), .C1(new_n574), .C2(new_n572), .ZN(new_n575));
  NAND2_X1  g150(.A1(G78), .A2(G543), .ZN(new_n576));
  INV_X1    g151(.A(G65), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n512), .B2(new_n577), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n578), .A2(G651), .B1(new_n530), .B2(G91), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT80), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n575), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n580), .B1(new_n575), .B2(new_n579), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n582), .A2(new_n583), .ZN(G299));
  INV_X1    g159(.A(G171), .ZN(G301));
  INV_X1    g160(.A(G166), .ZN(G303));
  AOI22_X1  g161(.A1(new_n530), .A2(G87), .B1(G49), .B2(new_n522), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n525), .B2(G74), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(G288));
  NAND2_X1  g164(.A1(new_n522), .A2(G48), .ZN(new_n590));
  INV_X1    g165(.A(G86), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n527), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n525), .A2(G61), .ZN(new_n593));
  NAND2_X1  g168(.A1(G73), .A2(G543), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n517), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(G305));
  NAND2_X1  g172(.A1(new_n522), .A2(G47), .ZN(new_n598));
  INV_X1    g173(.A(G85), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n527), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n525), .A2(G60), .ZN(new_n601));
  NAND2_X1  g176(.A1(G72), .A2(G543), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n517), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT81), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT10), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT82), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n530), .A2(new_n609), .A3(G92), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n609), .B1(new_n530), .B2(G92), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n608), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(G92), .ZN(new_n614));
  OAI21_X1  g189(.A(KEYINPUT82), .B1(new_n527), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n615), .A2(KEYINPUT10), .A3(new_n610), .ZN(new_n616));
  NAND2_X1  g191(.A1(G79), .A2(G543), .ZN(new_n617));
  INV_X1    g192(.A(G66), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n512), .B2(new_n618), .ZN(new_n619));
  AOI22_X1  g194(.A1(new_n619), .A2(G651), .B1(G54), .B2(new_n522), .ZN(new_n620));
  AND3_X1   g195(.A1(new_n613), .A2(new_n616), .A3(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n607), .B1(G868), .B2(new_n621), .ZN(G284));
  XOR2_X1   g197(.A(G284), .B(KEYINPUT83), .Z(G321));
  NAND2_X1  g198(.A1(G286), .A2(G868), .ZN(new_n624));
  INV_X1    g199(.A(G299), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(G868), .ZN(G280));
  XOR2_X1   g201(.A(G280), .B(KEYINPUT84), .Z(G297));
  INV_X1    g202(.A(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n621), .B1(new_n628), .B2(G860), .ZN(G148));
  NAND2_X1  g204(.A1(new_n621), .A2(new_n628), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(G868), .ZN(new_n631));
  INV_X1    g206(.A(new_n557), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n631), .B1(G868), .B2(new_n632), .ZN(G323));
  XNOR2_X1  g208(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g209(.A(KEYINPUT85), .B(KEYINPUT12), .ZN(new_n635));
  INV_X1    g210(.A(KEYINPUT3), .ZN(new_n636));
  INV_X1    g211(.A(G2104), .ZN(new_n637));
  NOR3_X1   g212(.A1(new_n636), .A2(new_n637), .A3(G2105), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n635), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT13), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2100), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n480), .A2(G135), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n482), .A2(G123), .ZN(new_n643));
  NOR2_X1   g218(.A1(G99), .A2(G2105), .ZN(new_n644));
  OAI21_X1  g219(.A(G2104), .B1(new_n463), .B2(G111), .ZN(new_n645));
  OAI211_X1 g220(.A(new_n642), .B(new_n643), .C1(new_n644), .C2(new_n645), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n646), .A2(G2096), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(G2096), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n641), .A2(new_n647), .A3(new_n648), .ZN(G156));
  XNOR2_X1  g224(.A(G2427), .B(G2438), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2430), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT15), .B(G2435), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n652), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n653), .A2(KEYINPUT14), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2443), .B(G2446), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n655), .B(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2451), .B(G2454), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  OAI21_X1  g239(.A(G14), .B1(new_n660), .B2(new_n664), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n665), .B1(new_n664), .B2(new_n660), .ZN(G401));
  XOR2_X1   g241(.A(G2072), .B(G2078), .Z(new_n667));
  XOR2_X1   g242(.A(G2084), .B(G2090), .Z(new_n668));
  XNOR2_X1  g243(.A(G2067), .B(G2678), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(KEYINPUT87), .B(KEYINPUT18), .Z(new_n671));
  AOI21_X1  g246(.A(new_n667), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  AND2_X1   g247(.A1(new_n670), .A2(KEYINPUT17), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n668), .A2(new_n669), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n671), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  MUX2_X1   g250(.A(new_n672), .B(new_n667), .S(new_n675), .Z(new_n676));
  XOR2_X1   g251(.A(G2096), .B(G2100), .Z(new_n677));
  XOR2_X1   g252(.A(new_n676), .B(new_n677), .Z(G227));
  XNOR2_X1  g253(.A(G1991), .B(G1996), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1971), .B(G1976), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT19), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G1956), .B(G2474), .Z(new_n686));
  XOR2_X1   g261(.A(G1961), .B(G1966), .Z(new_n687));
  AND2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(KEYINPUT20), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n686), .A2(new_n687), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  MUX2_X1   g268(.A(new_n693), .B(new_n692), .S(new_n685), .Z(new_n694));
  NOR2_X1   g269(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(KEYINPUT88), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT89), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n695), .B(KEYINPUT88), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n700), .A2(KEYINPUT89), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n682), .B1(new_n699), .B2(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1981), .B(G1986), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n700), .A2(KEYINPUT89), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n697), .A2(new_n698), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n705), .A2(new_n706), .A3(new_n681), .ZN(new_n707));
  AND3_X1   g282(.A1(new_n702), .A2(new_n704), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n704), .B1(new_n702), .B2(new_n707), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n680), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(new_n707), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n681), .B1(new_n705), .B2(new_n706), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n703), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n702), .A2(new_n704), .A3(new_n707), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n713), .A2(new_n714), .A3(new_n679), .ZN(new_n715));
  AND2_X1   g290(.A1(new_n710), .A2(new_n715), .ZN(G229));
  NOR2_X1   g291(.A1(G16), .A2(G22), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(G166), .B2(G16), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(G1971), .ZN(new_n719));
  INV_X1    g294(.A(G16), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(G6), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(new_n596), .B2(new_n720), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT32), .B(G1981), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n720), .A2(G23), .ZN(new_n725));
  INV_X1    g300(.A(G288), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n725), .B1(new_n726), .B2(new_n720), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT33), .B(G1976), .Z(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NOR3_X1   g304(.A1(new_n719), .A2(new_n724), .A3(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT34), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(G29), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G25), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n480), .A2(G131), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n482), .A2(G119), .ZN(new_n736));
  OR2_X1    g311(.A1(G95), .A2(G2105), .ZN(new_n737));
  OAI211_X1 g312(.A(new_n737), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n738));
  AND3_X1   g313(.A1(new_n735), .A2(new_n736), .A3(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n734), .B1(new_n739), .B2(new_n733), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT35), .B(G1991), .Z(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n720), .A2(G24), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n604), .A2(KEYINPUT90), .ZN(new_n744));
  OAI21_X1  g319(.A(G16), .B1(new_n604), .B2(KEYINPUT90), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n743), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n742), .B1(new_n746), .B2(G1986), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G1986), .B2(new_n746), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n730), .B2(new_n731), .ZN(new_n749));
  OR3_X1    g324(.A1(new_n732), .A2(new_n749), .A3(KEYINPUT36), .ZN(new_n750));
  OAI21_X1  g325(.A(KEYINPUT36), .B1(new_n732), .B2(new_n749), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n733), .A2(G35), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G162), .B2(new_n733), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT99), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT29), .B(G2090), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n720), .A2(G4), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(new_n621), .B2(new_n720), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n759), .A2(G1348), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n759), .A2(G1348), .ZN(new_n761));
  NOR3_X1   g336(.A1(new_n757), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n733), .A2(G26), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT28), .Z(new_n764));
  NAND2_X1  g339(.A1(new_n482), .A2(G128), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT93), .Z(new_n766));
  OAI21_X1  g341(.A(G2104), .B1(new_n463), .B2(G116), .ZN(new_n767));
  INV_X1    g342(.A(G104), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n767), .B1(new_n768), .B2(new_n463), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n480), .B2(G140), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n766), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n764), .B1(new_n771), .B2(G29), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G2067), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n720), .A2(G5), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G171), .B2(new_n720), .ZN(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(G1961), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n720), .A2(G19), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT91), .Z(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n632), .B2(new_n720), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT92), .B(G1341), .Z(new_n781));
  AOI22_X1  g356(.A1(new_n776), .A2(new_n777), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  OAI211_X1 g357(.A(new_n773), .B(new_n782), .C1(new_n777), .C2(new_n776), .ZN(new_n783));
  XOR2_X1   g358(.A(KEYINPUT31), .B(G11), .Z(new_n784));
  NOR2_X1   g359(.A1(new_n646), .A2(new_n733), .ZN(new_n785));
  INV_X1    g360(.A(G28), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n786), .A2(KEYINPUT30), .ZN(new_n787));
  AOI21_X1  g362(.A(G29), .B1(new_n786), .B2(KEYINPUT30), .ZN(new_n788));
  AOI211_X1 g363(.A(new_n784), .B(new_n785), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  AND2_X1   g364(.A1(KEYINPUT24), .A2(G34), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n733), .B1(KEYINPUT24), .B2(G34), .ZN(new_n791));
  OAI22_X1  g366(.A1(G160), .A2(new_n733), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(G2084), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  OAI211_X1 g369(.A(new_n789), .B(new_n794), .C1(new_n780), .C2(new_n781), .ZN(new_n795));
  NOR2_X1   g370(.A1(G168), .A2(new_n720), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(new_n720), .B2(G21), .ZN(new_n797));
  INV_X1    g372(.A(G1966), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n733), .A2(G33), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n480), .A2(G139), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT94), .B(KEYINPUT25), .Z(new_n802));
  NAND3_X1  g377(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  AOI22_X1  g379(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n805));
  OAI211_X1 g380(.A(new_n801), .B(new_n804), .C1(new_n463), .C2(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n800), .B1(new_n807), .B2(new_n733), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(G2072), .ZN(new_n809));
  OR3_X1    g384(.A1(new_n795), .A2(new_n799), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n797), .A2(new_n798), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT97), .Z(new_n812));
  NAND2_X1  g387(.A1(new_n733), .A2(G27), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(G164), .B2(new_n733), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(G2078), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT98), .ZN(new_n816));
  NOR4_X1   g391(.A1(new_n783), .A2(new_n810), .A3(new_n812), .A4(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n720), .A2(G20), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT23), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(new_n625), .B2(new_n720), .ZN(new_n820));
  INV_X1    g395(.A(G1956), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n733), .A2(G32), .ZN(new_n823));
  NAND3_X1  g398(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT26), .Z(new_n825));
  NAND3_X1  g400(.A1(new_n463), .A2(G105), .A3(G2104), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(new_n482), .B2(G129), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n480), .A2(KEYINPUT95), .A3(G141), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(KEYINPUT95), .B1(new_n480), .B2(G141), .ZN(new_n831));
  OAI211_X1 g406(.A(KEYINPUT96), .B(new_n828), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT95), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n478), .A2(new_n479), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(new_n463), .ZN(new_n836));
  INV_X1    g411(.A(G141), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n834), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(new_n829), .ZN(new_n839));
  AOI21_X1  g414(.A(KEYINPUT96), .B1(new_n839), .B2(new_n828), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n833), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n823), .B1(new_n841), .B2(new_n733), .ZN(new_n842));
  XNOR2_X1  g417(.A(KEYINPUT27), .B(G1996), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  AND3_X1   g419(.A1(new_n817), .A2(new_n822), .A3(new_n844), .ZN(new_n845));
  AND3_X1   g420(.A1(new_n752), .A2(new_n762), .A3(new_n845), .ZN(G311));
  NAND3_X1  g421(.A1(new_n752), .A2(new_n762), .A3(new_n845), .ZN(G150));
  NAND3_X1  g422(.A1(new_n613), .A2(new_n616), .A3(new_n620), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n848), .A2(new_n628), .ZN(new_n849));
  XOR2_X1   g424(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n522), .A2(G43), .ZN(new_n852));
  INV_X1    g427(.A(G81), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n852), .B1(new_n527), .B2(new_n853), .ZN(new_n854));
  AND2_X1   g429(.A1(new_n555), .A2(G651), .ZN(new_n855));
  NAND2_X1  g430(.A1(G80), .A2(G543), .ZN(new_n856));
  INV_X1    g431(.A(G67), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n856), .B1(new_n512), .B2(new_n857), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n858), .A2(G651), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n525), .A2(G93), .A3(new_n526), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n522), .A2(G55), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  OAI22_X1  g437(.A1(new_n854), .A2(new_n855), .B1(new_n859), .B2(new_n862), .ZN(new_n863));
  AOI22_X1  g438(.A1(new_n530), .A2(G93), .B1(G55), .B2(new_n522), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n858), .A2(G651), .ZN(new_n865));
  NAND4_X1  g440(.A1(new_n552), .A2(new_n864), .A3(new_n556), .A4(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n851), .B(new_n868), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n869), .A2(KEYINPUT39), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(KEYINPUT39), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n870), .A2(new_n558), .A3(new_n871), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n859), .A2(new_n862), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n873), .A2(new_n558), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT37), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n872), .A2(new_n875), .ZN(G145));
  INV_X1    g451(.A(KEYINPUT103), .ZN(new_n877));
  XOR2_X1   g452(.A(KEYINPUT101), .B(G37), .Z(new_n878));
  NAND2_X1  g453(.A1(new_n839), .A2(new_n828), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT96), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n881), .A2(new_n503), .A3(new_n832), .ZN(new_n882));
  OAI21_X1  g457(.A(G164), .B1(new_n833), .B2(new_n840), .ZN(new_n883));
  AND3_X1   g458(.A1(new_n882), .A2(new_n883), .A3(new_n806), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n806), .B1(new_n882), .B2(new_n883), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n771), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n882), .A2(new_n883), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(new_n807), .ZN(new_n888));
  INV_X1    g463(.A(new_n771), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n882), .A2(new_n883), .A3(new_n806), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n735), .A2(new_n736), .A3(new_n738), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n480), .A2(G142), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n482), .A2(G130), .ZN(new_n894));
  NOR2_X1   g469(.A1(G106), .A2(G2105), .ZN(new_n895));
  OAI21_X1  g470(.A(G2104), .B1(new_n463), .B2(G118), .ZN(new_n896));
  OAI211_X1 g471(.A(new_n893), .B(new_n894), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n892), .B(new_n897), .ZN(new_n898));
  AND2_X1   g473(.A1(new_n898), .A2(new_n639), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n898), .A2(new_n639), .ZN(new_n900));
  OAI21_X1  g475(.A(KEYINPUT102), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n886), .A2(new_n891), .A3(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n646), .B(G160), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(G162), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n901), .B1(new_n886), .B2(new_n891), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n878), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n899), .A2(new_n900), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n891), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n889), .B1(new_n888), .B2(new_n890), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n910), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n886), .A2(new_n891), .A3(new_n909), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n905), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n877), .B1(new_n908), .B2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n907), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n917), .A2(new_n905), .A3(new_n902), .ZN(new_n918));
  INV_X1    g493(.A(new_n914), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n909), .B1(new_n886), .B2(new_n891), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n904), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n918), .A2(new_n921), .A3(KEYINPUT103), .A4(new_n878), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n916), .A2(new_n922), .A3(KEYINPUT40), .ZN(new_n923));
  AOI21_X1  g498(.A(KEYINPUT40), .B1(new_n916), .B2(new_n922), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n923), .A2(new_n924), .ZN(G395));
  XNOR2_X1  g500(.A(new_n630), .B(new_n868), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n616), .A2(new_n620), .ZN(new_n927));
  INV_X1    g502(.A(new_n583), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n927), .A2(new_n928), .A3(new_n581), .A4(new_n613), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n848), .B1(new_n583), .B2(new_n582), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  OR3_X1    g507(.A1(new_n926), .A2(KEYINPUT104), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(KEYINPUT41), .B1(new_n929), .B2(new_n930), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n929), .A2(new_n930), .A3(KEYINPUT41), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n926), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(KEYINPUT104), .B1(new_n926), .B2(new_n932), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n933), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n596), .B(new_n604), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n529), .A2(new_n534), .A3(G288), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(G288), .B1(new_n529), .B2(new_n534), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n940), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n943), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n945), .A2(new_n941), .A3(new_n939), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n947), .B(KEYINPUT42), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n938), .B(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(G868), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n950), .B1(G868), .B2(new_n873), .ZN(G295));
  OAI21_X1  g526(.A(new_n950), .B1(G868), .B2(new_n873), .ZN(G331));
  INV_X1    g527(.A(KEYINPUT43), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n944), .A2(new_n946), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT106), .ZN(new_n955));
  AOI21_X1  g530(.A(G171), .B1(new_n955), .B2(G286), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n536), .A2(new_n541), .A3(KEYINPUT106), .A4(new_n542), .ZN(new_n958));
  AND3_X1   g533(.A1(new_n863), .A2(new_n866), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n958), .B1(new_n863), .B2(new_n866), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n957), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n958), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n867), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n863), .A2(new_n866), .A3(new_n958), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n963), .A2(new_n956), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n961), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n966), .B1(new_n935), .B2(new_n934), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n931), .A2(new_n961), .A3(new_n965), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n954), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  AND2_X1   g544(.A1(new_n969), .A2(new_n878), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT108), .ZN(new_n971));
  NOR3_X1   g546(.A1(new_n935), .A2(new_n934), .A3(new_n971), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n929), .A2(new_n930), .A3(new_n971), .A4(KEYINPUT41), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n966), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n968), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(new_n947), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n953), .B1(new_n970), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT41), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n931), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n929), .A2(new_n930), .A3(KEYINPUT41), .ZN(new_n980));
  AOI22_X1  g555(.A1(new_n979), .A2(new_n980), .B1(new_n965), .B2(new_n961), .ZN(new_n981));
  INV_X1    g556(.A(new_n968), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n947), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G37), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n983), .A2(new_n953), .A3(new_n969), .A4(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(KEYINPUT44), .ZN(new_n986));
  OAI21_X1  g561(.A(KEYINPUT110), .B1(new_n977), .B2(new_n986), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n966), .A2(new_n973), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n979), .A2(KEYINPUT108), .A3(new_n980), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n982), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  OAI211_X1 g565(.A(new_n878), .B(new_n969), .C1(new_n990), .C2(new_n954), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(KEYINPUT43), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT110), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n992), .A2(new_n993), .A3(KEYINPUT44), .A4(new_n985), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n987), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n969), .A2(new_n984), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n954), .B1(new_n968), .B2(new_n967), .ZN(new_n997));
  OAI21_X1  g572(.A(KEYINPUT43), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(KEYINPUT107), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT107), .ZN(new_n1000));
  OAI211_X1 g575(.A(new_n1000), .B(KEYINPUT43), .C1(new_n996), .C2(new_n997), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT109), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n1002), .B1(new_n991), .B2(KEYINPUT43), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n970), .A2(new_n976), .A3(KEYINPUT109), .A4(new_n953), .ZN(new_n1004));
  AOI22_X1  g579(.A1(new_n999), .A2(new_n1001), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g580(.A(KEYINPUT105), .B(KEYINPUT44), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n995), .B1(new_n1005), .B2(new_n1006), .ZN(G397));
  INV_X1    g582(.A(KEYINPUT127), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n771), .A2(G2067), .ZN(new_n1009));
  INV_X1    g584(.A(G2067), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n766), .A2(new_n1010), .A3(new_n770), .ZN(new_n1011));
  AND3_X1   g586(.A1(new_n1009), .A2(KEYINPUT114), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(KEYINPUT114), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n841), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G1996), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1015), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1016));
  XNOR2_X1  g591(.A(KEYINPUT111), .B(G1384), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n503), .A2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT45), .B1(new_n1018), .B2(KEYINPUT112), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1019), .B1(KEYINPUT112), .B2(new_n1018), .ZN(new_n1020));
  INV_X1    g595(.A(G125), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n636), .A2(new_n637), .ZN(new_n1022));
  NAND2_X1  g597(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1021), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n466), .ZN(new_n1025));
  OAI21_X1  g600(.A(G2105), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  AOI22_X1  g601(.A1(new_n464), .A2(new_n468), .B1(new_n472), .B2(new_n471), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1026), .A2(G40), .A3(new_n470), .A4(new_n1027), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1020), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1014), .A2(new_n1016), .A3(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n841), .A2(new_n1015), .A3(new_n1029), .ZN(new_n1031));
  XOR2_X1   g606(.A(new_n1031), .B(KEYINPUT113), .Z(new_n1032));
  NAND4_X1  g607(.A1(new_n1030), .A2(new_n741), .A3(new_n739), .A4(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n1011), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1008), .B1(new_n1034), .B2(new_n1029), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1029), .ZN(new_n1036));
  AOI211_X1 g611(.A(KEYINPUT127), .B(new_n1036), .C1(new_n1033), .C2(new_n1011), .ZN(new_n1037));
  XNOR2_X1  g612(.A(new_n739), .B(new_n741), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n1029), .ZN(new_n1039));
  NOR2_X1   g614(.A1(G290), .A2(G1986), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(new_n1029), .ZN(new_n1041));
  XNOR2_X1  g616(.A(new_n1041), .B(KEYINPUT48), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1030), .A2(new_n1039), .A3(new_n1032), .A4(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1014), .A2(new_n1029), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT47), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1029), .A2(new_n1015), .ZN(new_n1046));
  XNOR2_X1  g621(.A(new_n1046), .B(KEYINPUT46), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1044), .A2(new_n1045), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1045), .B1(new_n1044), .B2(new_n1047), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1043), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NOR3_X1   g626(.A1(new_n1035), .A2(new_n1037), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(G305), .A2(G1981), .ZN(new_n1053));
  INV_X1    g628(.A(G1981), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n596), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT49), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1053), .A2(KEYINPUT49), .A3(new_n1055), .ZN(new_n1059));
  INV_X1    g634(.A(G8), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1028), .ZN(new_n1061));
  AOI22_X1  g636(.A1(new_n490), .A2(new_n491), .B1(new_n501), .B2(new_n464), .ZN(new_n1062));
  AOI21_X1  g637(.A(G1384), .B1(new_n1062), .B2(new_n498), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1060), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1058), .A2(new_n1059), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(G1976), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1064), .B1(G288), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(KEYINPUT52), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n726), .A2(G1976), .ZN(new_n1069));
  OR3_X1    g644(.A1(new_n1069), .A2(new_n1067), .A3(KEYINPUT52), .ZN(new_n1070));
  AND3_X1   g645(.A1(new_n1065), .A2(new_n1068), .A3(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n529), .A2(new_n534), .A3(G8), .ZN(new_n1072));
  OR2_X1    g647(.A1(new_n1072), .A2(KEYINPUT55), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(KEYINPUT55), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(G1384), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n503), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT45), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1028), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n503), .A2(KEYINPUT45), .A3(new_n1017), .ZN(new_n1080));
  AND2_X1   g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  OR2_X1    g656(.A1(new_n1081), .A2(G1971), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1028), .B1(new_n1077), .B2(KEYINPUT50), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT50), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n503), .A2(new_n1084), .A3(new_n1076), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1082), .B1(G2090), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(G8), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1075), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT115), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1085), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1063), .A2(KEYINPUT115), .A3(new_n1084), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(new_n1083), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1082), .B1(new_n1094), .B2(G2090), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1073), .A2(G8), .A3(new_n1074), .A4(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n503), .A2(KEYINPUT45), .A3(new_n1076), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT117), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n503), .A2(KEYINPUT117), .A3(KEYINPUT45), .A4(new_n1076), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1099), .A2(new_n1100), .A3(new_n1061), .A4(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(new_n798), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1085), .A2(new_n1090), .ZN(new_n1104));
  AOI21_X1  g679(.A(KEYINPUT115), .B1(new_n1063), .B2(new_n1084), .ZN(new_n1105));
  OAI211_X1 g680(.A(new_n793), .B(new_n1083), .C1(new_n1104), .C2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1060), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1107));
  AND2_X1   g682(.A1(new_n1107), .A2(G168), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1071), .A2(new_n1089), .A3(new_n1096), .A4(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT63), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  AND4_X1   g686(.A1(new_n1096), .A2(new_n1065), .A3(new_n1068), .A4(new_n1070), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1095), .A2(G8), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1075), .A2(new_n1113), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1112), .A2(KEYINPUT63), .A3(new_n1108), .A4(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1111), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1065), .A2(new_n1066), .A3(new_n726), .ZN(new_n1117));
  XOR2_X1   g692(.A(new_n1055), .B(KEYINPUT116), .Z(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1096), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n1119), .A2(new_n1064), .B1(new_n1071), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1116), .A2(new_n1121), .ZN(new_n1122));
  XOR2_X1   g697(.A(KEYINPUT122), .B(KEYINPUT51), .Z(new_n1123));
  NAND2_X1  g698(.A1(G286), .A2(G8), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1124), .B1(new_n1107), .B2(KEYINPUT123), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT123), .ZN(new_n1126));
  AOI211_X1 g701(.A(new_n1126), .B(new_n1060), .C1(new_n1103), .C2(new_n1106), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1123), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT124), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  OAI211_X1 g705(.A(KEYINPUT124), .B(new_n1123), .C1(new_n1125), .C2(new_n1127), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1124), .ZN(new_n1132));
  NOR3_X1   g707(.A1(new_n1107), .A2(KEYINPUT51), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1130), .A2(new_n1131), .A3(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(new_n1132), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(G1348), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1094), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT119), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1061), .A2(new_n1141), .A3(new_n1063), .ZN(new_n1142));
  OAI21_X1  g717(.A(KEYINPUT119), .B1(new_n1077), .B2(new_n1028), .ZN(new_n1143));
  AOI21_X1  g718(.A(G2067), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1140), .A2(KEYINPUT60), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT60), .ZN(new_n1147));
  AOI21_X1  g722(.A(G1348), .B1(new_n1093), .B2(new_n1083), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1147), .B1(new_n1148), .B2(new_n1144), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1146), .A2(new_n1149), .A3(new_n621), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1140), .A2(KEYINPUT60), .A3(new_n1145), .A4(new_n848), .ZN(new_n1151));
  XOR2_X1   g726(.A(KEYINPUT58), .B(G1341), .Z(new_n1152));
  NAND3_X1  g727(.A1(new_n1142), .A2(new_n1143), .A3(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1079), .A2(new_n1015), .A3(new_n1080), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n557), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  OR2_X1    g730(.A1(new_n1155), .A2(KEYINPUT59), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(KEYINPUT59), .ZN(new_n1157));
  AND4_X1   g732(.A1(new_n1150), .A2(new_n1151), .A3(new_n1156), .A4(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT57), .ZN(new_n1159));
  AND3_X1   g734(.A1(new_n575), .A2(new_n579), .A3(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1159), .B1(new_n575), .B2(new_n579), .ZN(new_n1161));
  OR2_X1    g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT120), .ZN(new_n1163));
  XNOR2_X1  g738(.A(KEYINPUT56), .B(G2072), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1079), .A2(new_n1080), .A3(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT118), .ZN(new_n1166));
  AOI22_X1  g741(.A1(new_n1165), .A2(new_n1166), .B1(new_n1086), .B2(new_n821), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1079), .A2(KEYINPUT118), .A3(new_n1080), .A4(new_n1164), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1163), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1086), .A2(new_n821), .ZN(new_n1171));
  AND4_X1   g746(.A1(new_n1163), .A2(new_n1170), .A3(new_n1168), .A4(new_n1171), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1162), .B1(new_n1169), .B2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1170), .A2(new_n1168), .A3(new_n1171), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1174), .A2(new_n1162), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT61), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1173), .A2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1179), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1176), .B1(new_n1175), .B2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1158), .A2(new_n1178), .A3(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(new_n1175), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1174), .A2(KEYINPUT120), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1167), .A2(new_n1163), .A3(new_n1168), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1179), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n848), .B1(new_n1140), .B2(new_n1145), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1183), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1188), .A2(KEYINPUT121), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT121), .ZN(new_n1190));
  OAI211_X1 g765(.A(new_n1190), .B(new_n1183), .C1(new_n1186), .C2(new_n1187), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1182), .A2(new_n1189), .A3(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(G2078), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1081), .A2(new_n1193), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT53), .ZN(new_n1195));
  AOI22_X1  g770(.A1(new_n1194), .A2(new_n1195), .B1(new_n777), .B2(new_n1094), .ZN(new_n1196));
  XNOR2_X1  g771(.A(new_n474), .B(KEYINPUT125), .ZN(new_n1197));
  INV_X1    g772(.A(G40), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1193), .A2(KEYINPUT53), .ZN(new_n1199));
  NOR3_X1   g774(.A1(new_n467), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  NAND4_X1  g775(.A1(new_n1020), .A2(new_n1080), .A3(new_n1197), .A4(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1196), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1202), .A2(G171), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1203), .A2(KEYINPUT126), .ZN(new_n1204));
  INV_X1    g779(.A(KEYINPUT126), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n1202), .A2(new_n1205), .A3(G171), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1204), .A2(new_n1206), .ZN(new_n1207));
  OR2_X1    g782(.A1(new_n1102), .A2(new_n1199), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1196), .A2(new_n1208), .ZN(new_n1209));
  NOR2_X1   g784(.A1(new_n1209), .A2(G171), .ZN(new_n1210));
  INV_X1    g785(.A(KEYINPUT54), .ZN(new_n1211));
  NOR2_X1   g786(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1209), .A2(G171), .ZN(new_n1213));
  OAI21_X1  g788(.A(new_n1213), .B1(G171), .B2(new_n1202), .ZN(new_n1214));
  AOI22_X1  g789(.A1(new_n1207), .A2(new_n1212), .B1(new_n1211), .B2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g790(.A1(new_n1138), .A2(new_n1192), .A3(new_n1215), .ZN(new_n1216));
  INV_X1    g791(.A(new_n1213), .ZN(new_n1217));
  INV_X1    g792(.A(new_n1137), .ZN(new_n1218));
  AOI21_X1  g793(.A(new_n1133), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1219));
  AOI21_X1  g794(.A(new_n1218), .B1(new_n1219), .B2(new_n1131), .ZN(new_n1220));
  INV_X1    g795(.A(KEYINPUT62), .ZN(new_n1221));
  OAI21_X1  g796(.A(new_n1217), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  AOI211_X1 g797(.A(KEYINPUT62), .B(new_n1218), .C1(new_n1219), .C2(new_n1131), .ZN(new_n1223));
  OAI21_X1  g798(.A(new_n1216), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  AND2_X1   g799(.A1(new_n1112), .A2(new_n1089), .ZN(new_n1225));
  AOI21_X1  g800(.A(new_n1122), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  AND2_X1   g801(.A1(G290), .A2(G1986), .ZN(new_n1227));
  OAI21_X1  g802(.A(new_n1029), .B1(new_n1227), .B2(new_n1040), .ZN(new_n1228));
  NAND4_X1  g803(.A1(new_n1030), .A2(new_n1039), .A3(new_n1032), .A4(new_n1228), .ZN(new_n1229));
  OAI21_X1  g804(.A(new_n1052), .B1(new_n1226), .B2(new_n1229), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g805(.A1(new_n916), .A2(new_n922), .ZN(new_n1232));
  INV_X1    g806(.A(G227), .ZN(new_n1233));
  NAND2_X1  g807(.A1(G319), .A2(new_n1233), .ZN(new_n1234));
  AOI211_X1 g808(.A(G401), .B(new_n1234), .C1(new_n710), .C2(new_n715), .ZN(new_n1235));
  NAND2_X1  g809(.A1(new_n1232), .A2(new_n1235), .ZN(new_n1236));
  NOR2_X1   g810(.A1(new_n1236), .A2(new_n1005), .ZN(G308));
  AND2_X1   g811(.A1(new_n999), .A2(new_n1001), .ZN(new_n1238));
  AND2_X1   g812(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1239));
  OAI211_X1 g813(.A(new_n1232), .B(new_n1235), .C1(new_n1238), .C2(new_n1239), .ZN(G225));
endmodule


