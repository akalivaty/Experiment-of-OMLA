//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 1 0 1 1 1 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 0 0 1 1 0 1 0 1 0 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:01 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n783, new_n784, new_n785,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n993, new_n994, new_n995, new_n996, new_n997, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040;
  INV_X1    g000(.A(G953), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G227), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT78), .ZN(new_n189));
  XNOR2_X1  g003(.A(G110), .B(G140), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G104), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT3), .B1(new_n193), .B2(G107), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT3), .ZN(new_n195));
  INV_X1    g009(.A(G107), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n195), .A2(new_n196), .A3(G104), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n193), .A2(G107), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n194), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G101), .ZN(new_n200));
  INV_X1    g014(.A(G101), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n194), .A2(new_n197), .A3(new_n201), .A4(new_n198), .ZN(new_n202));
  AND3_X1   g016(.A1(new_n200), .A2(KEYINPUT4), .A3(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT4), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n199), .A2(new_n204), .A3(G101), .ZN(new_n205));
  XNOR2_X1  g019(.A(G143), .B(G146), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT0), .B(G128), .ZN(new_n207));
  OR2_X1    g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n206), .A2(KEYINPUT0), .A3(G128), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n205), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n203), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT80), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n212), .B1(new_n196), .B2(G104), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT79), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n214), .B1(new_n193), .B2(G107), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n193), .A2(KEYINPUT80), .A3(G107), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n196), .A2(KEYINPUT79), .A3(G104), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n213), .A2(new_n215), .A3(new_n216), .A4(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G101), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(new_n202), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(KEYINPUT82), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT82), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n219), .A2(new_n222), .A3(new_n202), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G128), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n226));
  INV_X1    g040(.A(G146), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G143), .ZN(new_n228));
  INV_X1    g042(.A(G143), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G146), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n226), .A2(new_n228), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT1), .B1(new_n229), .B2(G146), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT66), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT66), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n228), .A2(new_n235), .A3(KEYINPUT1), .ZN(new_n236));
  XNOR2_X1  g050(.A(KEYINPUT67), .B(G128), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n234), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n206), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n232), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT10), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n211), .B1(new_n224), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT68), .ZN(new_n244));
  INV_X1    g058(.A(G134), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G137), .ZN(new_n246));
  AND2_X1   g060(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n247));
  NOR2_X1   g061(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n245), .A2(G137), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G131), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT65), .ZN(new_n254));
  NAND2_X1  g068(.A1(KEYINPUT11), .A2(G134), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n254), .B1(new_n255), .B2(G137), .ZN(new_n256));
  INV_X1    g070(.A(G137), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n257), .A2(KEYINPUT65), .A3(KEYINPUT11), .A4(G134), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  AND3_X1   g073(.A1(new_n252), .A2(new_n253), .A3(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n253), .B1(new_n252), .B2(new_n259), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n244), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT64), .B(KEYINPUT11), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n250), .B1(new_n263), .B2(new_n246), .ZN(new_n264));
  AND2_X1   g078(.A1(new_n256), .A2(new_n258), .ZN(new_n265));
  OAI21_X1  g079(.A(G131), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  AOI22_X1  g080(.A1(new_n249), .A2(new_n251), .B1(new_n256), .B2(new_n258), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(new_n253), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n266), .A2(new_n268), .A3(KEYINPUT68), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n262), .A2(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n225), .B1(new_n228), .B2(KEYINPUT1), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n231), .B1(new_n271), .B2(new_n206), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n219), .A2(new_n272), .A3(new_n202), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(new_n241), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT81), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT81), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n273), .A2(new_n276), .A3(new_n241), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  AND3_X1   g092(.A1(new_n243), .A2(new_n270), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n240), .A2(new_n220), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n273), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n281), .A2(new_n269), .A3(new_n262), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT12), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n283), .B1(new_n266), .B2(new_n268), .ZN(new_n284));
  AOI22_X1  g098(.A1(new_n282), .A2(new_n283), .B1(new_n281), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n192), .B1(new_n279), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n238), .A2(new_n239), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n231), .ZN(new_n288));
  AND3_X1   g102(.A1(new_n219), .A2(new_n222), .A3(new_n202), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n222), .B1(new_n219), .B2(new_n202), .ZN(new_n290));
  OAI211_X1 g104(.A(KEYINPUT10), .B(new_n288), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n211), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n276), .B1(new_n273), .B2(new_n241), .ZN(new_n293));
  AND3_X1   g107(.A1(new_n273), .A2(new_n276), .A3(new_n241), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n291), .B(new_n292), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n270), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n243), .A2(new_n270), .A3(new_n278), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n297), .A2(new_n298), .A3(new_n191), .ZN(new_n299));
  AOI21_X1  g113(.A(G902), .B1(new_n286), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G469), .ZN(new_n301));
  OAI21_X1  g115(.A(KEYINPUT83), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n286), .A2(new_n299), .ZN(new_n303));
  INV_X1    g117(.A(G902), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT83), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n305), .A2(new_n306), .A3(G469), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n298), .A2(new_n191), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n308), .A2(new_n285), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n191), .B1(new_n297), .B2(new_n298), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n301), .B(new_n304), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n311), .A2(KEYINPUT84), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT84), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n270), .B1(new_n243), .B2(new_n278), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n192), .B1(new_n279), .B2(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(KEYINPUT12), .B1(new_n296), .B2(new_n281), .ZN(new_n316));
  AND2_X1   g130(.A1(new_n281), .A2(new_n284), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n298), .B(new_n191), .C1(new_n316), .C2(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(G902), .B1(new_n315), .B2(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n313), .B1(new_n319), .B2(new_n301), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n302), .B(new_n307), .C1(new_n312), .C2(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(G214), .B1(G237), .B2(G902), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G119), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G116), .ZN(new_n325));
  INV_X1    g139(.A(G116), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G119), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n325), .A2(new_n327), .A3(KEYINPUT5), .ZN(new_n328));
  OAI211_X1 g142(.A(new_n328), .B(G113), .C1(KEYINPUT5), .C2(new_n325), .ZN(new_n329));
  INV_X1    g143(.A(G113), .ZN(new_n330));
  AND2_X1   g144(.A1(new_n330), .A2(KEYINPUT2), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n330), .A2(KEYINPUT2), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n325), .B(new_n327), .C1(new_n331), .C2(new_n332), .ZN(new_n333));
  AND2_X1   g147(.A1(new_n329), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n334), .B1(new_n289), .B2(new_n290), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT85), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n325), .A2(new_n327), .ZN(new_n337));
  XNOR2_X1  g151(.A(KEYINPUT2), .B(G113), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n333), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(new_n205), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n336), .B1(new_n203), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n200), .A2(KEYINPUT4), .A3(new_n202), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n343), .A2(KEYINPUT85), .A3(new_n340), .A4(new_n205), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n335), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT86), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n335), .A2(new_n342), .A3(KEYINPUT86), .A4(new_n344), .ZN(new_n348));
  XNOR2_X1  g162(.A(G110), .B(G122), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n347), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n335), .A2(new_n342), .A3(new_n344), .A4(new_n349), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n352), .A2(KEYINPUT6), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n209), .B1(new_n206), .B2(new_n207), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(G125), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n357), .B1(G125), .B2(new_n240), .ZN(new_n358));
  INV_X1    g172(.A(G224), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n359), .A2(G953), .ZN(new_n360));
  XOR2_X1   g174(.A(new_n358), .B(new_n360), .Z(new_n361));
  INV_X1    g175(.A(KEYINPUT6), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n347), .A2(new_n362), .A3(new_n348), .A4(new_n350), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n354), .A2(new_n361), .A3(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n358), .B1(new_n359), .B2(G953), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n365), .B1(KEYINPUT87), .B2(new_n358), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(KEYINPUT7), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT7), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n360), .B1(KEYINPUT87), .B2(new_n368), .ZN(new_n369));
  OR2_X1    g183(.A1(new_n358), .A2(new_n369), .ZN(new_n370));
  OR2_X1    g184(.A1(new_n334), .A2(new_n220), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n334), .A2(new_n220), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n349), .B(KEYINPUT8), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  AND3_X1   g188(.A1(new_n370), .A2(new_n352), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(G902), .B1(new_n367), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n364), .A2(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(G210), .B1(G237), .B2(G902), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n364), .A2(new_n378), .A3(new_n376), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n323), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G221), .ZN(new_n383));
  XNOR2_X1  g197(.A(KEYINPUT9), .B(G234), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n383), .B1(new_n385), .B2(new_n304), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(G122), .ZN(new_n388));
  NOR3_X1   g202(.A1(new_n388), .A2(KEYINPUT14), .A3(G116), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT93), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n196), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(KEYINPUT14), .B1(new_n388), .B2(G116), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT14), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(new_n326), .A3(G122), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n388), .A2(G116), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n392), .A2(new_n394), .A3(KEYINPUT93), .A4(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT94), .ZN(new_n397));
  AND3_X1   g211(.A1(new_n391), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n397), .B1(new_n391), .B2(new_n396), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(G116), .B(G122), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n196), .ZN(new_n402));
  OR2_X1    g216(.A1(KEYINPUT67), .A2(G128), .ZN(new_n403));
  NAND2_X1  g217(.A1(KEYINPUT67), .A2(G128), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n403), .A2(G143), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n229), .A2(G128), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(new_n245), .A3(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n245), .B1(new_n405), .B2(new_n406), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n402), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(KEYINPUT95), .B1(new_n400), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n391), .A2(new_n396), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(KEYINPUT94), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n391), .A2(new_n396), .A3(new_n397), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT95), .ZN(new_n416));
  INV_X1    g230(.A(new_n409), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(new_n407), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n415), .A2(new_n416), .A3(new_n402), .A4(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n411), .A2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n405), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT13), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n406), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n229), .A2(KEYINPUT13), .A3(G128), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(G134), .B1(new_n421), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT92), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  OAI211_X1 g242(.A(KEYINPUT92), .B(G134), .C1(new_n421), .C2(new_n425), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n401), .B(new_n196), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT91), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n408), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n430), .B(new_n433), .C1(new_n432), .C2(new_n431), .ZN(new_n434));
  INV_X1    g248(.A(G217), .ZN(new_n435));
  NOR3_X1   g249(.A1(new_n384), .A2(new_n435), .A3(G953), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n420), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n436), .B1(new_n420), .B2(new_n434), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n304), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(G478), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT96), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n441), .A2(KEYINPUT15), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(KEYINPUT15), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n440), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n439), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n445), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n304), .B(new_n447), .C1(new_n437), .C2(new_n438), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT20), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT89), .ZN(new_n451));
  INV_X1    g265(.A(G140), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(G125), .ZN(new_n453));
  INV_X1    g267(.A(G125), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(G140), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n453), .A2(new_n455), .A3(KEYINPUT16), .ZN(new_n456));
  OR3_X1    g270(.A1(new_n454), .A2(KEYINPUT16), .A3(G140), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n227), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n456), .A2(new_n457), .A3(G146), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT17), .ZN(new_n462));
  INV_X1    g276(.A(G237), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n463), .A2(new_n187), .A3(G214), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT88), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n465), .A2(new_n229), .ZN(new_n466));
  NOR2_X1   g280(.A1(KEYINPUT88), .A2(G143), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g282(.A1(G237), .A2(G953), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n469), .B(G214), .C1(KEYINPUT88), .C2(G143), .ZN(new_n470));
  AOI211_X1 g284(.A(new_n462), .B(new_n253), .C1(new_n468), .C2(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n451), .B1(new_n461), .B2(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n253), .B1(new_n468), .B2(new_n470), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n468), .A2(new_n253), .A3(new_n470), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n474), .A2(new_n462), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n468), .A2(new_n470), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n477), .A2(KEYINPUT17), .A3(G131), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n478), .A2(KEYINPUT89), .A3(new_n459), .A4(new_n460), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n472), .A2(new_n476), .A3(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(G113), .B(G122), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n481), .B(new_n193), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n473), .A2(KEYINPUT18), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n453), .A2(new_n455), .ZN(new_n484));
  NOR3_X1   g298(.A1(new_n484), .A2(KEYINPUT76), .A3(G146), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT76), .ZN(new_n486));
  XNOR2_X1  g300(.A(G125), .B(G140), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n486), .B1(new_n487), .B2(new_n227), .ZN(new_n488));
  OAI22_X1  g302(.A1(new_n485), .A2(new_n488), .B1(new_n227), .B2(new_n487), .ZN(new_n489));
  AND2_X1   g303(.A1(KEYINPUT18), .A2(G131), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n483), .B(new_n489), .C1(new_n477), .C2(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n480), .A2(new_n482), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n474), .A2(new_n475), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n487), .A2(KEYINPUT19), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n487), .A2(KEYINPUT19), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n227), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n493), .A2(new_n460), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(new_n491), .ZN(new_n498));
  INV_X1    g312(.A(new_n482), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n492), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g315(.A1(G475), .A2(G902), .ZN(new_n502));
  XOR2_X1   g316(.A(new_n502), .B(KEYINPUT90), .Z(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n450), .B1(new_n501), .B2(new_n504), .ZN(new_n505));
  AOI211_X1 g319(.A(KEYINPUT20), .B(new_n503), .C1(new_n492), .C2(new_n500), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n480), .A2(new_n491), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n499), .ZN(new_n508));
  AOI21_X1  g322(.A(G902), .B1(new_n508), .B2(new_n492), .ZN(new_n509));
  INV_X1    g323(.A(G475), .ZN(new_n510));
  OAI22_X1  g324(.A1(new_n505), .A2(new_n506), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(G234), .A2(G237), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n512), .A2(G952), .A3(new_n187), .ZN(new_n513));
  XOR2_X1   g327(.A(new_n513), .B(KEYINPUT97), .Z(new_n514));
  AND3_X1   g328(.A1(new_n512), .A2(G902), .A3(G953), .ZN(new_n515));
  XNOR2_X1  g329(.A(KEYINPUT21), .B(G898), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n518), .B(KEYINPUT98), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NOR3_X1   g334(.A1(new_n449), .A2(new_n511), .A3(new_n520), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n321), .A2(new_n382), .A3(new_n387), .A4(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(KEYINPUT73), .B1(new_n324), .B2(G128), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT73), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n524), .A2(new_n225), .A3(G119), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n225), .A2(G119), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT23), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n523), .B(new_n525), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n403), .A2(KEYINPUT23), .A3(G119), .A4(new_n404), .ZN(new_n529));
  AND2_X1   g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(G110), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n237), .A2(new_n324), .ZN(new_n532));
  OR2_X1    g346(.A1(new_n532), .A2(new_n526), .ZN(new_n533));
  XNOR2_X1  g347(.A(KEYINPUT24), .B(G110), .ZN(new_n534));
  OAI221_X1 g348(.A(new_n461), .B1(new_n530), .B2(new_n531), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n485), .A2(new_n488), .ZN(new_n536));
  INV_X1    g350(.A(new_n460), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n528), .A2(new_n531), .A3(new_n529), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT74), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n534), .B1(new_n532), .B2(new_n526), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n528), .A2(KEYINPUT74), .A3(new_n531), .A4(new_n529), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT75), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n538), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AND2_X1   g360(.A1(new_n542), .A2(new_n543), .ZN(new_n547));
  AOI21_X1  g361(.A(KEYINPUT75), .B1(new_n547), .B2(new_n541), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n535), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  XNOR2_X1  g363(.A(KEYINPUT22), .B(G137), .ZN(new_n550));
  AND3_X1   g364(.A1(new_n187), .A2(G221), .A3(G234), .ZN(new_n551));
  XOR2_X1   g365(.A(new_n550), .B(new_n551), .Z(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n535), .B(new_n552), .C1(new_n546), .C2(new_n548), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n554), .A2(new_n304), .A3(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT77), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT25), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n435), .B1(G234), .B2(new_n304), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n556), .A2(new_n558), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n554), .A2(KEYINPUT25), .A3(new_n304), .A4(new_n555), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(KEYINPUT77), .A3(new_n564), .ZN(new_n565));
  AND2_X1   g379(.A1(new_n554), .A2(new_n555), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n560), .A2(G902), .ZN(new_n567));
  AOI22_X1  g381(.A1(new_n562), .A2(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(G472), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n463), .A2(new_n187), .A3(G210), .ZN(new_n570));
  XOR2_X1   g384(.A(new_n570), .B(KEYINPUT27), .Z(new_n571));
  XNOR2_X1  g385(.A(KEYINPUT26), .B(G101), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n571), .B(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT28), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT69), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n340), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n333), .A2(new_n339), .A3(KEYINPUT69), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n253), .B1(new_n251), .B2(new_n246), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n580), .B1(new_n267), .B2(new_n253), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n579), .B1(new_n288), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n262), .A2(new_n269), .A3(new_n356), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n288), .A2(new_n581), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n356), .B1(new_n260), .B2(new_n261), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(new_n340), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n575), .B1(new_n584), .B2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(KEYINPUT28), .B1(new_n582), .B2(new_n583), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n574), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT30), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n592), .B1(new_n288), .B2(new_n581), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n583), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n587), .A2(new_n592), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n594), .A2(new_n595), .A3(new_n340), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n596), .A2(new_n584), .A3(new_n573), .ZN(new_n597));
  AOI21_X1  g411(.A(KEYINPUT29), .B1(new_n591), .B2(new_n597), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n582), .A2(new_n583), .ZN(new_n599));
  INV_X1    g413(.A(new_n579), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n600), .B1(new_n583), .B2(new_n585), .ZN(new_n601));
  OAI21_X1  g415(.A(KEYINPUT28), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n262), .A2(new_n269), .A3(new_n356), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n600), .A2(new_n585), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n575), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(KEYINPUT71), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT71), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n590), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT29), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n573), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n602), .A2(new_n606), .A3(new_n608), .A4(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(new_n304), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n598), .B1(new_n612), .B2(KEYINPUT72), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT72), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n611), .A2(new_n614), .A3(new_n304), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n569), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n573), .B1(new_n589), .B2(new_n590), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n573), .B1(new_n582), .B2(new_n583), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n583), .A2(new_n593), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n266), .A2(new_n268), .ZN(new_n620));
  AOI22_X1  g434(.A1(new_n620), .A2(new_n356), .B1(new_n288), .B2(new_n581), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n340), .B1(new_n621), .B2(KEYINPUT30), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n618), .B1(new_n619), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(KEYINPUT31), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT31), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n596), .A2(new_n625), .A3(new_n618), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n617), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n569), .A2(new_n304), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(KEYINPUT70), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT32), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n627), .A2(KEYINPUT32), .A3(new_n629), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n568), .B1(new_n616), .B2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n522), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(KEYINPUT99), .B(G101), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G3));
  NAND3_X1  g452(.A1(new_n321), .A2(new_n568), .A3(new_n387), .ZN(new_n639));
  MUX2_X1   g453(.A(new_n304), .B(new_n439), .S(new_n440), .Z(new_n640));
  INV_X1    g454(.A(new_n438), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n420), .A2(new_n434), .A3(new_n436), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n436), .A2(KEYINPUT101), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT33), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AND3_X1   g459(.A1(new_n641), .A2(new_n642), .A3(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n645), .B1(new_n641), .B2(new_n642), .ZN(new_n647));
  OAI21_X1  g461(.A(G478), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n640), .A2(new_n648), .A3(new_n511), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n382), .A2(new_n650), .A3(new_n519), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n627), .A2(new_n304), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT100), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  OAI21_X1  g469(.A(G472), .B1(new_n652), .B2(new_n653), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n630), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NOR3_X1   g471(.A1(new_n639), .A2(new_n651), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(KEYINPUT34), .B(G104), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G6));
  INV_X1    g474(.A(KEYINPUT102), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n501), .A2(new_n661), .A3(new_n450), .A4(new_n504), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n662), .B1(new_n509), .B2(new_n510), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n505), .A2(new_n506), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n663), .B1(KEYINPUT102), .B2(new_n664), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n665), .A2(KEYINPUT103), .A3(new_n519), .A4(new_n449), .ZN(new_n666));
  INV_X1    g480(.A(new_n492), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n482), .B1(new_n480), .B2(new_n491), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n304), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  AOI22_X1  g483(.A1(new_n661), .A2(new_n506), .B1(new_n669), .B2(G475), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n501), .A2(new_n504), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(KEYINPUT20), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n501), .A2(new_n450), .A3(new_n504), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n672), .A2(KEYINPUT102), .A3(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n449), .A2(new_n670), .A3(new_n674), .A4(new_n519), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT103), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AND3_X1   g491(.A1(new_n382), .A2(new_n666), .A3(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n679), .A2(new_n657), .A3(new_n639), .ZN(new_n680));
  XNOR2_X1  g494(.A(KEYINPUT35), .B(G107), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G9));
  XNOR2_X1  g496(.A(new_n549), .B(KEYINPUT104), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n553), .A2(KEYINPUT36), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  OR2_X1    g500(.A1(new_n549), .A2(KEYINPUT104), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n549), .A2(KEYINPUT104), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n687), .A2(new_n684), .A3(new_n688), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n567), .ZN(new_n691));
  AND3_X1   g505(.A1(new_n563), .A2(KEYINPUT77), .A3(new_n564), .ZN(new_n692));
  OAI22_X1  g506(.A1(new_n690), .A2(new_n691), .B1(new_n692), .B2(new_n561), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n321), .A2(new_n382), .A3(new_n693), .A4(new_n387), .ZN(new_n694));
  OAI211_X1 g508(.A(new_n630), .B(new_n521), .C1(new_n655), .C2(new_n656), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(KEYINPUT37), .B(G110), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G12));
  NAND2_X1  g512(.A1(new_n670), .A2(new_n674), .ZN(new_n699));
  INV_X1    g513(.A(new_n449), .ZN(new_n700));
  XOR2_X1   g514(.A(new_n514), .B(KEYINPUT105), .Z(new_n701));
  INV_X1    g515(.A(G900), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n515), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n699), .A2(new_n700), .A3(new_n704), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n705), .B1(new_n616), .B2(new_n634), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n694), .A2(new_n706), .ZN(new_n707));
  XOR2_X1   g521(.A(KEYINPUT106), .B(G128), .Z(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G30));
  NAND2_X1  g523(.A1(new_n321), .A2(new_n387), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n704), .B(KEYINPUT39), .ZN(new_n711));
  OR2_X1    g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT108), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n712), .B(new_n713), .ZN(new_n714));
  AND2_X1   g528(.A1(new_n714), .A2(KEYINPUT40), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n714), .A2(KEYINPUT40), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n380), .A2(new_n381), .ZN(new_n717));
  XOR2_X1   g531(.A(new_n717), .B(KEYINPUT38), .Z(new_n718));
  NAND2_X1  g532(.A1(new_n596), .A2(new_n584), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n574), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n304), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n599), .A2(new_n601), .A3(new_n574), .ZN(new_n722));
  OAI21_X1  g536(.A(G472), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n632), .A2(new_n633), .A3(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(KEYINPUT107), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n323), .B1(new_n446), .B2(new_n448), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n511), .ZN(new_n727));
  OR4_X1    g541(.A1(new_n693), .A2(new_n718), .A3(new_n725), .A4(new_n727), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n715), .A2(new_n716), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(new_n229), .ZN(G45));
  INV_X1    g544(.A(new_n704), .ZN(new_n731));
  AND4_X1   g545(.A1(new_n511), .A2(new_n640), .A3(new_n648), .A4(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n321), .A2(new_n382), .A3(new_n732), .A4(new_n387), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n693), .B1(new_n616), .B2(new_n634), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(new_n227), .ZN(G48));
  AND3_X1   g550(.A1(new_n364), .A2(new_n378), .A3(new_n376), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n378), .B1(new_n364), .B2(new_n376), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n322), .B(new_n519), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n739), .A2(new_n649), .ZN(new_n740));
  AND3_X1   g554(.A1(new_n627), .A2(KEYINPUT32), .A3(new_n629), .ZN(new_n741));
  AOI21_X1  g555(.A(KEYINPUT32), .B1(new_n627), .B2(new_n629), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(new_n615), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n614), .B1(new_n611), .B2(new_n304), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n744), .A2(new_n745), .A3(new_n598), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n743), .B1(new_n746), .B2(new_n569), .ZN(new_n747));
  OR2_X1    g561(.A1(new_n319), .A2(new_n301), .ZN(new_n748));
  OAI211_X1 g562(.A(new_n387), .B(new_n748), .C1(new_n312), .C2(new_n320), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n740), .A2(new_n747), .A3(new_n750), .A4(new_n568), .ZN(new_n751));
  XNOR2_X1  g565(.A(KEYINPUT41), .B(G113), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n751), .B(new_n752), .ZN(G15));
  INV_X1    g567(.A(new_n566), .ZN(new_n754));
  OAI22_X1  g568(.A1(new_n692), .A2(new_n561), .B1(new_n754), .B2(new_n691), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n612), .A2(KEYINPUT72), .ZN(new_n756));
  INV_X1    g570(.A(new_n598), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n756), .A2(new_n615), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(G472), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n755), .B1(new_n759), .B2(new_n743), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n678), .A2(new_n760), .A3(new_n750), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G116), .ZN(G18));
  OAI21_X1  g576(.A(new_n322), .B1(new_n737), .B2(new_n738), .ZN(new_n763));
  INV_X1    g577(.A(new_n511), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n700), .A2(new_n764), .A3(new_n519), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n749), .A2(new_n763), .A3(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n691), .B1(new_n686), .B2(new_n689), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n767), .B1(new_n562), .B2(new_n565), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n768), .B1(new_n759), .B2(new_n743), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G119), .ZN(G21));
  AND3_X1   g585(.A1(new_n602), .A2(new_n606), .A3(new_n608), .ZN(new_n772));
  OAI211_X1 g586(.A(new_n624), .B(new_n626), .C1(new_n772), .C2(new_n574), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n629), .B(KEYINPUT109), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n652), .A2(G472), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n777), .A2(new_n755), .ZN(new_n778));
  OAI211_X1 g592(.A(new_n511), .B(new_n726), .C1(new_n737), .C2(new_n738), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n778), .A2(new_n750), .A3(new_n519), .A4(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G122), .ZN(G24));
  NOR2_X1   g596(.A1(new_n749), .A2(new_n763), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n777), .A2(new_n768), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n783), .A2(new_n784), .A3(new_n732), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G125), .ZN(G27));
  NAND4_X1  g600(.A1(new_n380), .A2(new_n387), .A3(new_n322), .A4(new_n381), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n301), .B1(new_n303), .B2(new_n304), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n789), .B1(new_n312), .B2(new_n320), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(KEYINPUT110), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n311), .A2(KEYINPUT84), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n319), .A2(new_n313), .A3(new_n301), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT110), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n794), .A2(new_n795), .A3(new_n789), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n787), .B1(new_n791), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n797), .A2(KEYINPUT42), .A3(new_n732), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n742), .B1(KEYINPUT112), .B2(new_n633), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n799), .B1(KEYINPUT112), .B2(new_n633), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n568), .B1(new_n800), .B2(new_n616), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT111), .ZN(new_n803));
  INV_X1    g617(.A(new_n787), .ZN(new_n804));
  AOI211_X1 g618(.A(KEYINPUT110), .B(new_n788), .C1(new_n792), .C2(new_n793), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n795), .B1(new_n794), .B2(new_n789), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n732), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n807), .A2(new_n635), .A3(new_n808), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n803), .B1(new_n809), .B2(KEYINPUT42), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n797), .A2(new_n760), .A3(new_n732), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT42), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n811), .A2(KEYINPUT111), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n802), .B1(new_n810), .B2(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(new_n253), .ZN(G33));
  NAND2_X1  g629(.A1(new_n791), .A2(new_n796), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n816), .A2(new_n760), .A3(new_n705), .A4(new_n804), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT113), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n797), .A2(KEYINPUT113), .A3(new_n760), .A4(new_n705), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(G134), .ZN(G36));
  INV_X1    g636(.A(KEYINPUT45), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n301), .B1(new_n303), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n824), .B1(new_n823), .B2(new_n303), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT114), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n301), .A2(new_n304), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n829), .A2(KEYINPUT46), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n794), .B1(new_n829), .B2(KEYINPUT46), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n387), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  OR2_X1    g646(.A1(new_n832), .A2(new_n711), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n764), .A2(new_n640), .A3(new_n648), .ZN(new_n834));
  XOR2_X1   g648(.A(new_n834), .B(KEYINPUT43), .Z(new_n835));
  NAND3_X1  g649(.A1(new_n835), .A2(new_n657), .A3(new_n693), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT44), .ZN(new_n837));
  OR2_X1    g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n717), .A2(new_n323), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n836), .A2(new_n837), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n833), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(new_n257), .ZN(G39));
  XOR2_X1   g657(.A(new_n832), .B(KEYINPUT47), .Z(new_n844));
  INV_X1    g658(.A(new_n839), .ZN(new_n845));
  NOR4_X1   g659(.A1(new_n845), .A2(new_n747), .A3(new_n808), .A4(new_n568), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(G140), .ZN(G42));
  NOR3_X1   g662(.A1(new_n834), .A2(new_n386), .A3(new_n323), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n794), .A2(new_n748), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT49), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n849), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n853), .B1(new_n852), .B2(new_n851), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n854), .A2(new_n568), .A3(new_n718), .A4(new_n725), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n855), .B(KEYINPUT115), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n761), .A2(new_n770), .A3(new_n751), .A4(new_n781), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n857), .B(KEYINPUT116), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n784), .A2(new_n732), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n699), .A2(new_n449), .A3(new_n704), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n839), .A2(new_n387), .A3(new_n321), .A4(new_n861), .ZN(new_n862));
  OAI22_X1  g676(.A1(new_n807), .A2(new_n860), .B1(new_n862), .B2(new_n734), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n863), .B1(new_n819), .B2(new_n820), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n700), .A2(new_n511), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n382), .A2(new_n519), .A3(new_n865), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n639), .A2(new_n866), .A3(new_n657), .ZN(new_n867));
  OAI21_X1  g681(.A(KEYINPUT117), .B1(new_n867), .B2(new_n696), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n321), .A2(new_n387), .ZN(new_n869));
  INV_X1    g683(.A(new_n865), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n870), .A2(new_n739), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n627), .A2(new_n304), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n569), .B1(new_n872), .B2(KEYINPUT100), .ZN(new_n873));
  AOI22_X1  g687(.A1(new_n873), .A2(new_n654), .B1(new_n629), .B2(new_n627), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n869), .A2(new_n871), .A3(new_n568), .A4(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT117), .ZN(new_n876));
  OAI211_X1 g690(.A(new_n875), .B(new_n876), .C1(new_n694), .C2(new_n695), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n658), .A2(new_n636), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n864), .A2(new_n868), .A3(new_n877), .A4(new_n878), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n859), .A2(new_n879), .A3(new_n814), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT53), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OR2_X1    g696(.A1(new_n694), .A2(new_n706), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n869), .A2(new_n769), .A3(new_n382), .A4(new_n732), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n704), .A2(new_n386), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n724), .A2(new_n768), .A3(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n816), .A2(new_n886), .A3(new_n780), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n883), .A2(new_n884), .A3(new_n887), .A4(new_n785), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT52), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n707), .A2(new_n735), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n891), .A2(KEYINPUT52), .A3(new_n785), .A4(new_n887), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT118), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n890), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n893), .B1(new_n890), .B2(new_n892), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(new_n863), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n821), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n877), .A2(new_n868), .A3(new_n878), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(new_n813), .ZN(new_n901));
  AOI21_X1  g715(.A(KEYINPUT111), .B1(new_n811), .B2(new_n812), .ZN(new_n902));
  OAI22_X1  g716(.A1(new_n901), .A2(new_n902), .B1(new_n801), .B2(new_n798), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n890), .A2(new_n892), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n900), .A2(new_n903), .A3(new_n904), .A4(new_n858), .ZN(new_n905));
  AOI22_X1  g719(.A1(new_n882), .A2(new_n896), .B1(KEYINPUT53), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(KEYINPUT54), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n904), .A2(KEYINPUT118), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n890), .A2(new_n892), .A3(new_n893), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n857), .A2(KEYINPUT119), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n794), .A2(new_n387), .A3(new_n519), .A4(new_n748), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n912), .A2(new_n779), .ZN(new_n913));
  AOI22_X1  g727(.A1(new_n769), .A2(new_n766), .B1(new_n913), .B2(new_n778), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT119), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n914), .A2(new_n915), .A3(new_n751), .A4(new_n761), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n911), .A2(KEYINPUT53), .A3(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n900), .A2(new_n903), .A3(new_n917), .ZN(new_n918));
  OAI21_X1  g732(.A(KEYINPUT120), .B1(new_n910), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n911), .A2(KEYINPUT53), .A3(new_n916), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n879), .A2(new_n814), .A3(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT120), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n896), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT54), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n905), .A2(new_n881), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n919), .A2(new_n923), .A3(new_n924), .A4(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n907), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n725), .A2(new_n568), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n750), .A2(new_n839), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n928), .A2(new_n514), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n511), .B1(new_n640), .B2(new_n648), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(new_n784), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n835), .A2(new_n701), .ZN(new_n934));
  OR2_X1    g748(.A1(new_n934), .A2(new_n929), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n934), .A2(new_n755), .A3(new_n777), .ZN(new_n936));
  AND3_X1   g750(.A1(new_n718), .A2(new_n323), .A3(new_n750), .ZN(new_n937));
  AND3_X1   g751(.A1(new_n936), .A2(KEYINPUT50), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(KEYINPUT50), .B1(new_n936), .B2(new_n937), .ZN(new_n939));
  OAI221_X1 g753(.A(new_n932), .B1(new_n933), .B2(new_n935), .C1(new_n938), .C2(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n850), .A2(new_n387), .ZN(new_n941));
  OR2_X1    g755(.A1(new_n844), .A2(new_n941), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n936), .A2(new_n839), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n940), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n944), .A2(KEYINPUT51), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n936), .A2(new_n783), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n946), .A2(G952), .A3(new_n187), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n935), .A2(new_n801), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT48), .ZN(new_n949));
  AOI211_X1 g763(.A(new_n947), .B(new_n949), .C1(new_n650), .C2(new_n930), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n950), .B1(new_n944), .B2(KEYINPUT51), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n927), .A2(new_n945), .A3(new_n951), .ZN(new_n952));
  NOR2_X1   g766(.A1(G952), .A2(G953), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n856), .B1(new_n952), .B2(new_n953), .ZN(G75));
  NOR2_X1   g768(.A1(new_n187), .A2(G952), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n919), .A2(new_n923), .A3(new_n925), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n957), .A2(G902), .ZN(new_n958));
  AOI21_X1  g772(.A(KEYINPUT56), .B1(new_n958), .B2(G210), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n354), .A2(new_n363), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(new_n361), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT55), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n956), .B1(new_n959), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n964), .B1(new_n959), .B2(new_n963), .ZN(G51));
  NAND2_X1  g779(.A1(new_n957), .A2(KEYINPUT54), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT121), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n966), .A2(new_n967), .A3(new_n926), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n957), .A2(KEYINPUT121), .A3(KEYINPUT54), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n828), .B(KEYINPUT57), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n971), .B1(new_n310), .B2(new_n309), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n958), .A2(new_n827), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n955), .B1(new_n972), .B2(new_n973), .ZN(G54));
  NAND4_X1  g788(.A1(new_n958), .A2(KEYINPUT58), .A3(G475), .A4(new_n501), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT122), .ZN(new_n976));
  OR2_X1    g790(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n975), .A2(new_n976), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n958), .A2(KEYINPUT58), .A3(G475), .ZN(new_n979));
  INV_X1    g793(.A(new_n501), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n955), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  AND3_X1   g795(.A1(new_n977), .A2(new_n978), .A3(new_n981), .ZN(G60));
  NOR2_X1   g796(.A1(new_n646), .A2(new_n647), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n440), .A2(new_n304), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT59), .Z(new_n985));
  AND2_X1   g799(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n968), .A2(new_n969), .A3(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT123), .ZN(new_n988));
  AND3_X1   g802(.A1(new_n987), .A2(new_n988), .A3(new_n956), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n988), .B1(new_n987), .B2(new_n956), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n983), .B1(new_n927), .B2(new_n985), .ZN(new_n991));
  NOR3_X1   g805(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(G63));
  NAND2_X1  g806(.A1(G217), .A2(G902), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n993), .B(KEYINPUT60), .Z(new_n994));
  NAND2_X1  g808(.A1(new_n957), .A2(new_n994), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n955), .B1(new_n995), .B2(new_n754), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n996), .B1(new_n690), .B2(new_n995), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n997), .B(KEYINPUT61), .Z(G66));
  INV_X1    g812(.A(new_n516), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n187), .B1(new_n999), .B2(G224), .ZN(new_n1000));
  OR2_X1    g814(.A1(new_n859), .A2(new_n899), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n1000), .B1(new_n1001), .B2(new_n187), .ZN(new_n1002));
  INV_X1    g816(.A(G898), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n960), .B1(new_n1003), .B2(G953), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1002), .B(new_n1004), .ZN(G69));
  NAND2_X1  g819(.A1(new_n891), .A2(new_n785), .ZN(new_n1006));
  OR3_X1    g820(.A1(new_n729), .A2(KEYINPUT62), .A3(new_n1006), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n842), .B1(new_n844), .B2(new_n846), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n870), .A2(new_n649), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n1009), .B(KEYINPUT124), .ZN(new_n1010));
  OR4_X1    g824(.A1(new_n635), .A2(new_n714), .A3(new_n845), .A4(new_n1010), .ZN(new_n1011));
  OAI21_X1  g825(.A(KEYINPUT62), .B1(new_n729), .B2(new_n1006), .ZN(new_n1012));
  NAND4_X1  g826(.A1(new_n1007), .A2(new_n1008), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1013), .A2(new_n187), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n594), .A2(new_n595), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n494), .A2(new_n495), .ZN(new_n1016));
  XOR2_X1   g830(.A(new_n1015), .B(new_n1016), .Z(new_n1017));
  NAND2_X1  g831(.A1(new_n1014), .A2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1017), .B1(G900), .B2(G953), .ZN(new_n1019));
  NOR3_X1   g833(.A1(new_n833), .A2(new_n779), .A3(new_n801), .ZN(new_n1020));
  INV_X1    g834(.A(new_n821), .ZN(new_n1021));
  NOR3_X1   g835(.A1(new_n1020), .A2(new_n1021), .A3(new_n1006), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n1022), .A2(new_n903), .A3(new_n1008), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n1019), .B1(new_n1023), .B2(G953), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1018), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n187), .B1(G227), .B2(G900), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1026), .B1(new_n1024), .B2(KEYINPUT125), .ZN(new_n1027));
  XOR2_X1   g841(.A(new_n1025), .B(new_n1027), .Z(G72));
  XOR2_X1   g842(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n1029));
  NOR2_X1   g843(.A1(new_n569), .A2(new_n304), .ZN(new_n1030));
  XNOR2_X1  g844(.A(new_n1029), .B(new_n1030), .ZN(new_n1031));
  OAI21_X1  g845(.A(new_n1031), .B1(new_n1013), .B2(new_n1001), .ZN(new_n1032));
  NAND3_X1  g846(.A1(new_n1032), .A2(new_n574), .A3(new_n719), .ZN(new_n1033));
  OAI21_X1  g847(.A(new_n1031), .B1(new_n1023), .B2(new_n1001), .ZN(new_n1034));
  INV_X1    g848(.A(new_n597), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g850(.A1(new_n1033), .A2(new_n956), .A3(new_n1036), .ZN(new_n1037));
  NAND4_X1  g851(.A1(new_n906), .A2(new_n597), .A3(new_n720), .A4(new_n1031), .ZN(new_n1038));
  OR2_X1    g852(.A1(new_n1038), .A2(KEYINPUT127), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1038), .A2(KEYINPUT127), .ZN(new_n1040));
  AOI21_X1  g854(.A(new_n1037), .B1(new_n1039), .B2(new_n1040), .ZN(G57));
endmodule


