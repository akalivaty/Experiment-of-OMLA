//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 1 0 1 1 1 1 1 1 1 0 0 1 1 0 0 0 1 1 0 0 0 1 1 1 0 1 0 0 0 0 1 0 1 1 1 1 0 0 0 0 1 0 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:20 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  XOR2_X1   g001(.A(G125), .B(G140), .Z(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(G146), .ZN(new_n189));
  INV_X1    g003(.A(G140), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(KEYINPUT70), .A3(G125), .ZN(new_n191));
  AND3_X1   g005(.A1(KEYINPUT70), .A2(KEYINPUT71), .A3(G125), .ZN(new_n192));
  OAI21_X1  g006(.A(G140), .B1(KEYINPUT71), .B2(G125), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n191), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(KEYINPUT83), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT83), .ZN(new_n196));
  OAI211_X1 g010(.A(new_n196), .B(new_n191), .C1(new_n192), .C2(new_n193), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n189), .B1(new_n198), .B2(G146), .ZN(new_n199));
  INV_X1    g013(.A(G237), .ZN(new_n200));
  INV_X1    g014(.A(G953), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n200), .A2(new_n201), .A3(G214), .ZN(new_n202));
  INV_X1    g016(.A(G143), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NOR2_X1   g018(.A1(G237), .A2(G953), .ZN(new_n205));
  AOI21_X1  g019(.A(G143), .B1(new_n205), .B2(G214), .ZN(new_n206));
  OAI21_X1  g020(.A(G131), .B1(new_n204), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT18), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n202), .A2(new_n203), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n205), .A2(G143), .A3(G214), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(KEYINPUT18), .A2(G131), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  OAI22_X1  g027(.A1(new_n207), .A2(new_n208), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT84), .B1(new_n199), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G131), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n216), .B1(new_n209), .B2(new_n210), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n204), .A2(new_n206), .ZN(new_n218));
  AOI22_X1  g032(.A1(KEYINPUT18), .A2(new_n217), .B1(new_n218), .B2(new_n212), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT84), .ZN(new_n220));
  INV_X1    g034(.A(G146), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n221), .B1(new_n195), .B2(new_n197), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n219), .B(new_n220), .C1(new_n189), .C2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n215), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g038(.A(G113), .B(G122), .ZN(new_n225));
  INV_X1    g039(.A(G104), .ZN(new_n226));
  XNOR2_X1  g040(.A(new_n225), .B(new_n226), .ZN(new_n227));
  OAI211_X1 g041(.A(KEYINPUT16), .B(new_n191), .C1(new_n192), .C2(new_n193), .ZN(new_n228));
  NOR2_X1   g042(.A1(KEYINPUT16), .A2(G140), .ZN(new_n229));
  AND2_X1   g043(.A1(KEYINPUT71), .A2(G125), .ZN(new_n230));
  NOR2_X1   g044(.A1(KEYINPUT71), .A2(G125), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n229), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n228), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(new_n221), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n228), .A2(G146), .A3(new_n232), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n234), .A2(KEYINPUT72), .A3(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT72), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n228), .A2(new_n237), .A3(G146), .A4(new_n232), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n217), .A2(KEYINPUT17), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT17), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n209), .A2(new_n216), .A3(new_n210), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n207), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n239), .A2(new_n240), .A3(new_n243), .ZN(new_n244));
  AND3_X1   g058(.A1(new_n224), .A2(new_n227), .A3(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n227), .B1(new_n224), .B2(new_n244), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n187), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G475), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT20), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n224), .A2(new_n244), .A3(new_n227), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n195), .A2(KEYINPUT19), .A3(new_n197), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT19), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n188), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(KEYINPUT85), .B1(new_n254), .B2(new_n221), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n235), .A2(KEYINPUT73), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT73), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n228), .A2(new_n257), .A3(new_n232), .A4(G146), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n207), .A2(new_n242), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n255), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n254), .A2(KEYINPUT85), .A3(new_n221), .ZN(new_n263));
  AOI22_X1  g077(.A1(new_n262), .A2(new_n263), .B1(new_n223), .B2(new_n215), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n250), .B1(new_n264), .B2(new_n227), .ZN(new_n265));
  NOR2_X1   g079(.A1(G475), .A2(G902), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n249), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n254), .A2(new_n221), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT85), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  AND2_X1   g084(.A1(new_n259), .A2(new_n260), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n270), .A2(new_n271), .A3(new_n263), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n227), .B1(new_n272), .B2(new_n224), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n249), .B(new_n266), .C1(new_n273), .C2(new_n245), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n248), .B1(new_n267), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(G952), .ZN(new_n277));
  AOI211_X1 g091(.A(G953), .B(new_n277), .C1(G234), .C2(G237), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  AOI211_X1 g093(.A(new_n187), .B(new_n201), .C1(G234), .C2(G237), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  XOR2_X1   g095(.A(KEYINPUT21), .B(G898), .Z(new_n282));
  OAI21_X1  g096(.A(new_n279), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n283), .B(KEYINPUT87), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(G122), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(G116), .ZN(new_n287));
  INV_X1    g101(.A(G116), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G122), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(G107), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n287), .A2(new_n289), .A3(G107), .ZN(new_n293));
  AND2_X1   g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n203), .A2(G128), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT13), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G128), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(G143), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n295), .A2(new_n296), .ZN(new_n301));
  OAI21_X1  g115(.A(G134), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G134), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n295), .A2(new_n299), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(KEYINPUT86), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT86), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n294), .A2(new_n302), .A3(new_n306), .A4(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n287), .A2(KEYINPUT14), .A3(G107), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n292), .A2(new_n293), .A3(new_n310), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n287), .A2(new_n289), .A3(KEYINPUT14), .A4(G107), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n303), .B1(new_n295), .B2(new_n299), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n311), .B(new_n312), .C1(new_n305), .C2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n309), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(KEYINPUT9), .B(G234), .ZN(new_n316));
  INV_X1    g130(.A(G217), .ZN(new_n317));
  NOR3_X1   g131(.A1(new_n316), .A2(new_n317), .A3(G953), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n315), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n309), .A2(new_n314), .A3(new_n318), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(new_n187), .ZN(new_n323));
  INV_X1    g137(.A(G478), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n324), .A2(KEYINPUT15), .ZN(new_n325));
  XOR2_X1   g139(.A(new_n323), .B(new_n325), .Z(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  NOR3_X1   g141(.A1(new_n276), .A2(new_n285), .A3(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(G210), .B1(G237), .B2(G902), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n221), .A2(G143), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n203), .A2(G146), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NOR2_X1   g147(.A1(KEYINPUT0), .A2(G128), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT0), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n335), .A2(new_n298), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n333), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  XNOR2_X1  g151(.A(G143), .B(G146), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n338), .B1(new_n335), .B2(new_n298), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n230), .A2(new_n231), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n337), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT82), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(KEYINPUT1), .B1(new_n203), .B2(G146), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT67), .ZN(new_n346));
  OAI21_X1  g160(.A(G128), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(KEYINPUT67), .B1(new_n331), .B2(KEYINPUT1), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n333), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n298), .A2(KEYINPUT1), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n338), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n349), .A2(new_n351), .A3(new_n340), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n337), .A2(new_n339), .A3(KEYINPUT82), .A4(new_n341), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n344), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(G224), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n355), .A2(G953), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n356), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n344), .A2(new_n352), .A3(new_n358), .A4(new_n353), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  XNOR2_X1  g175(.A(G110), .B(G122), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT3), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n363), .A2(new_n291), .A3(G104), .ZN(new_n364));
  AOI21_X1  g178(.A(KEYINPUT3), .B1(new_n226), .B2(G107), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n226), .A2(G107), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G101), .ZN(new_n368));
  INV_X1    g182(.A(G101), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n369), .B(new_n364), .C1(new_n365), .C2(new_n366), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n368), .A2(KEYINPUT4), .A3(new_n370), .ZN(new_n371));
  XNOR2_X1  g185(.A(G116), .B(G119), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  OR2_X1    g187(.A1(KEYINPUT2), .A2(G113), .ZN(new_n374));
  AND3_X1   g188(.A1(KEYINPUT68), .A2(KEYINPUT2), .A3(G113), .ZN(new_n375));
  AOI21_X1  g189(.A(KEYINPUT68), .B1(KEYINPUT2), .B2(G113), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n374), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n373), .A2(new_n377), .ZN(new_n378));
  OAI211_X1 g192(.A(new_n372), .B(new_n374), .C1(new_n376), .C2(new_n375), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT4), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n367), .A2(new_n381), .A3(G101), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n371), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n291), .A2(G104), .ZN(new_n384));
  OAI21_X1  g198(.A(G101), .B1(new_n366), .B2(new_n384), .ZN(new_n385));
  AND2_X1   g199(.A1(new_n370), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT5), .ZN(new_n387));
  INV_X1    g201(.A(G119), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n387), .A2(new_n388), .A3(G116), .ZN(new_n389));
  OAI211_X1 g203(.A(G113), .B(new_n389), .C1(new_n373), .C2(new_n387), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n386), .A2(new_n379), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n362), .B1(new_n383), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT80), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(KEYINPUT6), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n392), .B(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n383), .A2(new_n362), .A3(new_n391), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(KEYINPUT81), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT81), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n383), .A2(new_n398), .A3(new_n362), .A4(new_n391), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n397), .A2(KEYINPUT6), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n361), .B1(new_n395), .B2(new_n400), .ZN(new_n401));
  AND2_X1   g215(.A1(new_n397), .A2(new_n399), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n362), .B(KEYINPUT8), .ZN(new_n403));
  INV_X1    g217(.A(new_n391), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n386), .B1(new_n379), .B2(new_n390), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n403), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n352), .A2(new_n342), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT7), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n407), .B1(new_n408), .B2(new_n356), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n406), .B(new_n409), .C1(new_n408), .C2(new_n359), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n187), .B1(new_n402), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n330), .B1(new_n401), .B2(new_n411), .ZN(new_n412));
  AND3_X1   g226(.A1(new_n397), .A2(KEYINPUT6), .A3(new_n399), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n383), .A2(new_n391), .ZN(new_n414));
  INV_X1    g228(.A(new_n362), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(new_n394), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n392), .A2(new_n393), .A3(KEYINPUT6), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n360), .B1(new_n413), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n406), .A2(new_n409), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n359), .A2(new_n408), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n397), .A2(new_n399), .ZN(new_n424));
  AOI21_X1  g238(.A(G902), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n420), .A2(new_n425), .A3(new_n329), .ZN(new_n426));
  AND2_X1   g240(.A1(new_n412), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(G214), .B1(G237), .B2(G902), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  AOI22_X1  g244(.A1(new_n345), .A2(G128), .B1(new_n331), .B2(new_n332), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n351), .B1(new_n431), .B2(KEYINPUT78), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n298), .B1(new_n331), .B2(KEYINPUT1), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT78), .ZN(new_n434));
  NOR3_X1   g248(.A1(new_n433), .A2(new_n338), .A3(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n386), .B1(new_n432), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT10), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT64), .ZN(new_n439));
  INV_X1    g253(.A(G137), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n439), .B1(new_n440), .B2(G134), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n303), .A2(KEYINPUT64), .A3(G137), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(KEYINPUT11), .B1(new_n440), .B2(G134), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n440), .A2(KEYINPUT11), .A3(G134), .ZN(new_n446));
  AND4_X1   g260(.A1(new_n216), .A2(new_n443), .A3(new_n445), .A4(new_n446), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n440), .A2(KEYINPUT11), .A3(G134), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n448), .A2(new_n444), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n216), .B1(new_n449), .B2(new_n443), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n337), .A2(new_n339), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n371), .A2(new_n452), .A3(new_n382), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n349), .A2(new_n351), .ZN(new_n454));
  AND3_X1   g268(.A1(new_n370), .A2(KEYINPUT10), .A3(new_n385), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n438), .A2(new_n451), .A3(new_n453), .A4(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(G110), .B(G140), .ZN(new_n458));
  INV_X1    g272(.A(G227), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n459), .A2(G953), .ZN(new_n460));
  XOR2_X1   g274(.A(new_n458), .B(new_n460), .Z(new_n461));
  NAND2_X1  g275(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(KEYINPUT79), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT79), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n457), .A2(new_n464), .A3(new_n461), .ZN(new_n465));
  INV_X1    g279(.A(new_n451), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n453), .A2(new_n456), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n431), .A2(KEYINPUT78), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n434), .B1(new_n433), .B2(new_n338), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n468), .A2(new_n469), .A3(new_n351), .ZN(new_n470));
  AOI21_X1  g284(.A(KEYINPUT10), .B1(new_n470), .B2(new_n386), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n466), .B1(new_n467), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n463), .A2(new_n465), .A3(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n461), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT12), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n370), .A2(new_n385), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n349), .A2(new_n351), .A3(new_n476), .ZN(new_n477));
  AOI211_X1 g291(.A(new_n475), .B(new_n451), .C1(new_n436), .C2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n436), .A2(new_n477), .ZN(new_n479));
  AOI21_X1  g293(.A(KEYINPUT12), .B1(new_n479), .B2(new_n466), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n457), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n474), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n473), .A2(G469), .A3(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(G469), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n481), .A2(new_n462), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n461), .B1(new_n472), .B2(new_n457), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n485), .B(new_n187), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n485), .A2(new_n187), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n484), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(G221), .B1(new_n316), .B2(G902), .ZN(new_n492));
  XOR2_X1   g306(.A(new_n492), .B(KEYINPUT77), .Z(new_n493));
  AND2_X1   g307(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n328), .A2(new_n430), .A3(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n452), .B1(new_n447), .B2(new_n450), .ZN(new_n496));
  OAI21_X1  g310(.A(KEYINPUT65), .B1(new_n303), .B2(G137), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT65), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n498), .A2(new_n440), .A3(G134), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n303), .A2(G137), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n497), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(G131), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT66), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n449), .A2(new_n216), .A3(new_n443), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n501), .A2(KEYINPUT66), .A3(G131), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n351), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT1), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n509), .B1(G143), .B2(new_n221), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(KEYINPUT67), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n345), .A2(new_n346), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n511), .A2(G128), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n508), .B1(new_n513), .B2(new_n333), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n496), .B1(new_n507), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n380), .ZN(new_n516));
  INV_X1    g330(.A(new_n380), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n496), .B(new_n517), .C1(new_n507), .C2(new_n514), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n516), .A2(KEYINPUT28), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n515), .A2(KEYINPUT69), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT69), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n496), .B(new_n521), .C1(new_n507), .C2(new_n514), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n380), .A2(KEYINPUT28), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n520), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n205), .A2(G210), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n525), .B(G101), .ZN(new_n526));
  XNOR2_X1  g340(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n526), .B(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n519), .A2(new_n524), .A3(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT30), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n515), .A2(new_n531), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n496), .B(KEYINPUT30), .C1(new_n507), .C2(new_n514), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n532), .A2(new_n380), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n534), .A2(new_n528), .A3(new_n518), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT31), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n530), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(G472), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n534), .A2(KEYINPUT31), .A3(new_n528), .A4(new_n518), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n537), .A2(new_n538), .A3(new_n187), .A4(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT32), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n529), .B1(new_n519), .B2(new_n524), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n528), .B1(new_n534), .B2(new_n518), .ZN(new_n544));
  NOR3_X1   g358(.A1(new_n543), .A2(new_n544), .A3(KEYINPUT29), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n519), .A2(new_n524), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n546), .A2(KEYINPUT29), .A3(new_n528), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n187), .ZN(new_n548));
  OAI21_X1  g362(.A(G472), .B1(new_n545), .B2(new_n548), .ZN(new_n549));
  AND2_X1   g363(.A1(new_n539), .A2(new_n187), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n550), .A2(KEYINPUT32), .A3(new_n538), .A4(new_n537), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n542), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n317), .B1(G234), .B2(new_n187), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(KEYINPUT22), .B(G137), .ZN(new_n555));
  AND3_X1   g369(.A1(new_n201), .A2(G221), .A3(G234), .ZN(new_n556));
  XOR2_X1   g370(.A(new_n555), .B(new_n556), .Z(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  XOR2_X1   g372(.A(G119), .B(G128), .Z(new_n559));
  XNOR2_X1  g373(.A(KEYINPUT24), .B(G110), .ZN(new_n560));
  OR2_X1    g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(KEYINPUT23), .B1(new_n388), .B2(G128), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT23), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n563), .A2(new_n298), .A3(G119), .ZN(new_n564));
  AOI22_X1  g378(.A1(new_n562), .A2(new_n564), .B1(new_n388), .B2(G128), .ZN(new_n565));
  INV_X1    g379(.A(G110), .ZN(new_n566));
  OR2_X1    g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n236), .A2(new_n238), .A3(new_n561), .A4(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT74), .ZN(new_n569));
  AOI22_X1  g383(.A1(new_n565), .A2(new_n566), .B1(new_n559), .B2(new_n560), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n570), .A2(new_n189), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n259), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n569), .B1(new_n259), .B2(new_n571), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n568), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT75), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n558), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n259), .A2(new_n571), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(KEYINPUT74), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n259), .A2(new_n571), .A3(new_n569), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(KEYINPUT75), .B1(new_n580), .B2(new_n568), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n576), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n574), .A2(new_n575), .A3(new_n557), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n187), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n554), .B1(new_n585), .B2(KEYINPUT25), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n574), .A2(new_n575), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n580), .A2(KEYINPUT75), .A3(new_n568), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n587), .A2(new_n588), .A3(new_n558), .ZN(new_n589));
  AOI211_X1 g403(.A(KEYINPUT25), .B(G902), .C1(new_n589), .C2(new_n583), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n586), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n589), .A2(new_n583), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n553), .A2(G902), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n593), .A2(KEYINPUT76), .A3(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(KEYINPUT76), .B1(new_n593), .B2(new_n594), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n552), .A2(new_n592), .A3(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n495), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(new_n369), .ZN(G3));
  AOI21_X1  g415(.A(new_n318), .B1(new_n309), .B2(new_n314), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT33), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT90), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n321), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n309), .A2(new_n314), .A3(KEYINPUT90), .A4(new_n318), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n604), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(KEYINPUT91), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT91), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n604), .A2(new_n610), .A3(new_n606), .A4(new_n607), .ZN(new_n611));
  INV_X1    g425(.A(new_n321), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n603), .B1(new_n612), .B2(new_n602), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT89), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n322), .A2(KEYINPUT89), .A3(new_n603), .ZN(new_n616));
  AOI22_X1  g430(.A1(new_n609), .A2(new_n611), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n324), .A2(G902), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n323), .A2(new_n324), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n276), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n622), .A2(new_n285), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n550), .A2(new_n537), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(G472), .ZN(new_n626));
  AND2_X1   g440(.A1(new_n626), .A2(new_n540), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n627), .A2(new_n592), .A3(new_n598), .A4(new_n494), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT88), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n412), .A2(new_n426), .A3(new_n629), .ZN(new_n630));
  OAI211_X1 g444(.A(new_n630), .B(new_n428), .C1(new_n629), .C2(new_n426), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n624), .A2(new_n628), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(new_n226), .ZN(new_n633));
  XNOR2_X1  g447(.A(KEYINPUT92), .B(KEYINPUT34), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G6));
  NOR2_X1   g449(.A1(new_n276), .A2(new_n326), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n284), .ZN(new_n637));
  NOR3_X1   g451(.A1(new_n628), .A2(new_n631), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(KEYINPUT35), .B(G107), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G9));
  NOR2_X1   g454(.A1(new_n558), .A2(KEYINPUT36), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n574), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n594), .ZN(new_n643));
  AOI21_X1  g457(.A(G902), .B1(new_n589), .B2(new_n583), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT25), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n553), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n643), .B1(new_n646), .B2(new_n590), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n627), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n495), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(KEYINPUT37), .B(G110), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G12));
  OAI21_X1  g465(.A(new_n428), .B1(new_n426), .B2(new_n629), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n652), .B1(new_n427), .B2(new_n629), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n653), .A2(new_n552), .A3(new_n647), .A4(new_n494), .ZN(new_n654));
  INV_X1    g468(.A(G900), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n278), .B1(new_n280), .B2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n636), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(new_n298), .ZN(G30));
  NAND2_X1  g474(.A1(new_n542), .A2(new_n551), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n516), .A2(new_n518), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n529), .ZN(new_n663));
  OR2_X1    g477(.A1(new_n663), .A2(KEYINPUT94), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(KEYINPUT94), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n664), .A2(new_n535), .A3(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n538), .B1(new_n666), .B2(new_n187), .ZN(new_n667));
  OR2_X1    g481(.A1(new_n661), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g482(.A(new_n668), .B(KEYINPUT95), .Z(new_n669));
  XOR2_X1   g483(.A(KEYINPUT93), .B(KEYINPUT38), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n427), .B(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n276), .A2(new_n327), .ZN(new_n672));
  OR4_X1    g486(.A1(new_n429), .A2(new_n671), .A3(new_n647), .A4(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n656), .B(KEYINPUT39), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n494), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(KEYINPUT40), .ZN(new_n677));
  OR3_X1    g491(.A1(new_n669), .A2(new_n673), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G143), .ZN(G45));
  NAND3_X1  g493(.A1(new_n276), .A2(new_n621), .A3(new_n657), .ZN(new_n680));
  OAI21_X1  g494(.A(KEYINPUT96), .B1(new_n654), .B2(new_n680), .ZN(new_n681));
  AND3_X1   g495(.A1(new_n542), .A2(new_n549), .A3(new_n551), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n682), .A2(new_n631), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n647), .A2(new_n494), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT96), .ZN(new_n685));
  INV_X1    g499(.A(new_n680), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n683), .A2(new_n684), .A3(new_n685), .A4(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n681), .A2(new_n687), .ZN(new_n688));
  XOR2_X1   g502(.A(KEYINPUT97), .B(G146), .Z(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G48));
  AOI21_X1  g504(.A(new_n451), .B1(new_n436), .B2(new_n477), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(KEYINPUT12), .ZN(new_n692));
  AND2_X1   g506(.A1(new_n457), .A2(new_n461), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n472), .A2(new_n457), .ZN(new_n694));
  AOI22_X1  g508(.A1(new_n692), .A2(new_n693), .B1(new_n694), .B2(new_n474), .ZN(new_n695));
  OAI21_X1  g509(.A(G469), .B1(new_n695), .B2(G902), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT98), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n696), .A2(new_n697), .A3(new_n488), .ZN(new_n698));
  OAI211_X1 g512(.A(KEYINPUT98), .B(G469), .C1(new_n695), .C2(G902), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g514(.A(KEYINPUT99), .B1(new_n700), .B2(new_n492), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT99), .ZN(new_n702));
  INV_X1    g516(.A(new_n492), .ZN(new_n703));
  AOI211_X1 g517(.A(new_n702), .B(new_n703), .C1(new_n698), .C2(new_n699), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n701), .A2(new_n704), .A3(new_n631), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n593), .A2(new_n594), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT76), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI211_X1 g522(.A(new_n708), .B(new_n595), .C1(new_n646), .C2(new_n590), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n705), .A2(new_n552), .A3(new_n710), .A4(new_n623), .ZN(new_n711));
  XNOR2_X1  g525(.A(KEYINPUT41), .B(G113), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(G15));
  INV_X1    g527(.A(new_n637), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n705), .A2(new_n552), .A3(new_n710), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G116), .ZN(G18));
  AND2_X1   g530(.A1(new_n328), .A2(new_n647), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n705), .A2(new_n552), .A3(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G119), .ZN(G21));
  INV_X1    g533(.A(KEYINPUT100), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n626), .A2(new_n540), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n720), .B1(new_n709), .B2(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n627), .A2(new_n592), .A3(new_n598), .A4(KEYINPUT100), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n701), .A2(new_n704), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n631), .A2(new_n672), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n724), .A2(new_n284), .A3(new_n725), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G122), .ZN(G24));
  INV_X1    g542(.A(KEYINPUT101), .ZN(new_n729));
  INV_X1    g543(.A(new_n643), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n730), .B1(new_n586), .B2(new_n591), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n729), .B1(new_n731), .B2(new_n721), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n627), .A2(new_n647), .A3(KEYINPUT101), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT102), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n680), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n276), .A2(new_n621), .A3(KEYINPUT102), .A4(new_n657), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n705), .A2(new_n734), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G125), .ZN(G27));
  INV_X1    g554(.A(KEYINPUT105), .ZN(new_n741));
  AND3_X1   g555(.A1(new_n412), .A2(new_n426), .A3(new_n428), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT103), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n742), .A2(new_n743), .A3(new_n492), .A4(new_n491), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n491), .A2(new_n492), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n412), .A2(new_n426), .A3(new_n428), .ZN(new_n746));
  OAI21_X1  g560(.A(KEYINPUT103), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n599), .B1(new_n744), .B2(new_n747), .ZN(new_n748));
  AOI21_X1  g562(.A(KEYINPUT42), .B1(new_n748), .B2(new_n738), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n747), .A2(new_n744), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n738), .A2(KEYINPUT42), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n661), .A2(KEYINPUT104), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT104), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n542), .A2(new_n753), .A3(new_n551), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n752), .A2(new_n549), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n710), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n751), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n741), .B1(new_n749), .B2(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n682), .A2(new_n709), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n738), .A2(new_n759), .A3(new_n750), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT42), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n761), .B1(new_n736), .B2(new_n737), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n763), .A2(new_n710), .A3(new_n750), .A4(new_n755), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n762), .A2(KEYINPUT105), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n758), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G131), .ZN(G33));
  AOI211_X1 g581(.A(new_n658), .B(new_n599), .C1(new_n744), .C2(new_n747), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(new_n303), .ZN(G36));
  AND2_X1   g583(.A1(new_n473), .A2(new_n483), .ZN(new_n770));
  OR2_X1    g584(.A1(new_n770), .A2(KEYINPUT45), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(KEYINPUT45), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n771), .A2(G469), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n490), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT46), .ZN(new_n775));
  OAI21_X1  g589(.A(KEYINPUT106), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT106), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n773), .A2(new_n777), .A3(KEYINPUT46), .A4(new_n490), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n774), .A2(new_n775), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n776), .A2(new_n488), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n492), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n781), .A2(new_n674), .ZN(new_n782));
  OR2_X1    g596(.A1(new_n267), .A2(new_n275), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n783), .A2(new_n248), .A3(new_n621), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(KEYINPUT43), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n786), .A2(new_n721), .A3(new_n647), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT44), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n746), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  OAI211_X1 g603(.A(new_n782), .B(new_n789), .C1(new_n788), .C2(new_n787), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G137), .ZN(G39));
  INV_X1    g605(.A(KEYINPUT47), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n792), .A2(KEYINPUT107), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n781), .A2(new_n793), .ZN(new_n794));
  NOR4_X1   g608(.A1(new_n710), .A2(new_n552), .A3(new_n680), .A4(new_n746), .ZN(new_n795));
  AOI22_X1  g609(.A1(new_n780), .A2(new_n492), .B1(KEYINPUT107), .B2(new_n792), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n794), .B(new_n795), .C1(new_n793), .C2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G140), .ZN(G42));
  AND2_X1   g612(.A1(new_n669), .A2(new_n710), .ZN(new_n799));
  INV_X1    g613(.A(new_n784), .ZN(new_n800));
  AND4_X1   g614(.A1(new_n428), .A2(new_n671), .A3(new_n493), .A4(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n700), .B(KEYINPUT49), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n799), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT54), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT108), .ZN(new_n805));
  INV_X1    g619(.A(new_n768), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n734), .A2(new_n738), .A3(new_n750), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n276), .A2(new_n327), .A3(new_n656), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n684), .A2(new_n552), .A3(new_n742), .A4(new_n808), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n762), .A2(KEYINPUT105), .A3(new_n764), .ZN(new_n811));
  AOI21_X1  g625(.A(KEYINPUT105), .B1(new_n762), .B2(new_n764), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n806), .B(new_n810), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n711), .A2(new_n727), .A3(new_n718), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n495), .B1(new_n599), .B2(new_n648), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n628), .B1(new_n624), .B2(new_n637), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n815), .B1(new_n816), .B2(new_n430), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n814), .A2(new_n715), .A3(new_n817), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n805), .B1(new_n813), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n768), .B1(new_n758), .B2(new_n765), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n711), .A2(new_n715), .A3(new_n727), .A4(new_n718), .ZN(new_n821));
  INV_X1    g635(.A(new_n817), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n820), .A2(KEYINPUT108), .A3(new_n823), .A4(new_n810), .ZN(new_n824));
  INV_X1    g638(.A(new_n659), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n647), .A2(new_n656), .A3(new_n745), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n826), .A2(new_n668), .A3(new_n726), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n688), .A2(new_n739), .A3(new_n825), .A4(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(KEYINPUT52), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n659), .B1(new_n681), .B2(new_n687), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT52), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n830), .A2(new_n831), .A3(new_n739), .A4(new_n827), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n819), .A2(new_n824), .A3(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT53), .ZN(new_n835));
  OR2_X1    g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  OR2_X1    g650(.A1(new_n836), .A2(KEYINPUT110), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT109), .ZN(new_n838));
  AOI22_X1  g652(.A1(new_n829), .A2(new_n832), .B1(new_n838), .B2(new_n828), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n828), .A2(new_n838), .A3(new_n831), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n841), .A2(new_n819), .A3(new_n824), .ZN(new_n842));
  AOI22_X1  g656(.A1(new_n836), .A2(KEYINPUT110), .B1(new_n835), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n804), .B1(new_n837), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n785), .A2(new_n279), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n671), .A2(new_n429), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n845), .A2(new_n725), .A3(new_n724), .A4(new_n846), .ZN(new_n847));
  XOR2_X1   g661(.A(new_n847), .B(KEYINPUT50), .Z(new_n848));
  NOR3_X1   g662(.A1(new_n701), .A2(new_n704), .A3(new_n746), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT113), .ZN(new_n850));
  OR2_X1    g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n279), .B1(new_n849), .B2(new_n850), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n853), .A2(new_n734), .A3(new_n786), .ZN(new_n854));
  INV_X1    g668(.A(new_n276), .ZN(new_n855));
  INV_X1    g669(.A(new_n621), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n853), .A2(new_n799), .A3(new_n855), .A4(new_n856), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n848), .A2(new_n854), .A3(new_n857), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n845), .A2(new_n724), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(new_n742), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n794), .B1(new_n796), .B2(new_n793), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n493), .B1(new_n698), .B2(new_n699), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n860), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT112), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n858), .B(new_n865), .C1(new_n866), .C2(KEYINPUT51), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n853), .A2(new_n786), .ZN(new_n868));
  INV_X1    g682(.A(new_n756), .ZN(new_n869));
  XOR2_X1   g683(.A(KEYINPUT115), .B(KEYINPUT48), .Z(new_n870));
  NAND3_X1  g684(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n853), .A2(new_n799), .A3(new_n276), .A4(new_n621), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n859), .A2(new_n725), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT114), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n874), .B1(new_n277), .B2(G953), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n201), .A2(KEYINPUT114), .A3(G952), .ZN(new_n876));
  AOI22_X1  g690(.A1(new_n873), .A2(new_n653), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n871), .A2(new_n872), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n870), .B1(new_n868), .B2(new_n869), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n848), .A2(new_n866), .A3(new_n854), .A4(new_n857), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT51), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n848), .A2(new_n854), .A3(new_n857), .ZN(new_n883));
  OAI211_X1 g697(.A(new_n881), .B(new_n882), .C1(new_n883), .C2(new_n864), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n867), .A2(new_n880), .A3(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT116), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n867), .A2(KEYINPUT116), .A3(new_n884), .A4(new_n880), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT111), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n762), .A2(new_n764), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n814), .A2(new_n890), .A3(new_n715), .A4(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n891), .ZN(new_n893));
  OAI21_X1  g707(.A(KEYINPUT111), .B1(new_n821), .B2(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n768), .A2(new_n835), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n810), .A2(new_n817), .A3(new_n895), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n892), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  AOI221_X4 g711(.A(KEYINPUT54), .B1(new_n841), .B2(new_n897), .C1(new_n834), .C2(new_n835), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n844), .A2(new_n889), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n277), .A2(new_n201), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT117), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n803), .B1(new_n899), .B2(new_n901), .ZN(G75));
  NAND2_X1  g716(.A1(new_n834), .A2(new_n835), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n841), .A2(new_n897), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n187), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(KEYINPUT56), .B1(new_n905), .B2(G210), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n413), .A2(new_n419), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(new_n360), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT55), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n906), .A2(new_n909), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n201), .A2(G952), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(G51));
  INV_X1    g727(.A(KEYINPUT118), .ZN(new_n914));
  INV_X1    g728(.A(new_n912), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n903), .A2(new_n904), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(KEYINPUT54), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n903), .A2(new_n804), .A3(new_n904), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n489), .B(KEYINPUT57), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n695), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  AOI211_X1 g735(.A(new_n187), .B(new_n773), .C1(new_n903), .C2(new_n904), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n914), .B(new_n915), .C1(new_n921), .C2(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n804), .B1(new_n903), .B2(new_n904), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n920), .B1(new_n898), .B2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n695), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n922), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(KEYINPUT118), .B1(new_n927), .B2(new_n912), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n923), .A2(new_n928), .ZN(G54));
  NAND3_X1  g743(.A1(new_n905), .A2(KEYINPUT58), .A3(G475), .ZN(new_n930));
  INV_X1    g744(.A(new_n265), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n930), .A2(new_n931), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n932), .A2(new_n933), .A3(new_n912), .ZN(G60));
  INV_X1    g748(.A(new_n919), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n617), .B(KEYINPUT119), .Z(new_n936));
  XNOR2_X1  g750(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n324), .A2(new_n187), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n937), .B(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  OR2_X1    g754(.A1(new_n936), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n915), .B1(new_n935), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n939), .B1(new_n844), .B2(new_n898), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n942), .B1(new_n943), .B2(new_n936), .ZN(G63));
  NAND2_X1  g758(.A1(G217), .A2(G902), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT60), .Z(new_n946));
  AOI21_X1  g760(.A(new_n593), .B1(new_n916), .B2(new_n946), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n947), .A2(new_n912), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT121), .ZN(new_n949));
  AOI21_X1  g763(.A(KEYINPUT61), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n916), .A2(new_n642), .A3(new_n946), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n948), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  OAI211_X1 g767(.A(new_n948), .B(new_n951), .C1(new_n949), .C2(KEYINPUT61), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(G66));
  INV_X1    g769(.A(new_n282), .ZN(new_n956));
  OAI21_X1  g770(.A(G953), .B1(new_n956), .B2(new_n355), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n957), .B1(new_n823), .B2(G953), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n907), .B1(G898), .B2(new_n201), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT122), .Z(new_n960));
  XNOR2_X1  g774(.A(new_n958), .B(new_n960), .ZN(G69));
  NAND2_X1  g775(.A1(new_n532), .A2(new_n533), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(new_n254), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n655), .A2(G953), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n790), .A2(new_n797), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n782), .A2(new_n726), .A3(new_n869), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n820), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n830), .A2(new_n739), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(KEYINPUT124), .ZN(new_n969));
  NOR3_X1   g783(.A1(new_n965), .A2(new_n967), .A3(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n964), .B1(new_n970), .B2(G953), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n963), .B1(new_n971), .B2(KEYINPUT125), .ZN(new_n972));
  INV_X1    g786(.A(new_n636), .ZN(new_n973));
  AOI211_X1 g787(.A(new_n746), .B(new_n676), .C1(new_n622), .C2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(new_n759), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n790), .A2(new_n797), .A3(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT124), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n968), .B(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(new_n678), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT62), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n978), .A2(KEYINPUT62), .A3(new_n678), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n976), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g797(.A(KEYINPUT123), .B1(new_n983), .B2(G953), .ZN(new_n984));
  OAI211_X1 g798(.A(new_n972), .B(new_n984), .C1(KEYINPUT125), .C2(new_n971), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n983), .A2(G953), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n963), .B1(new_n986), .B2(KEYINPUT123), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g802(.A(G953), .B1(new_n459), .B2(new_n655), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(new_n989), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n985), .A2(new_n987), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n990), .A2(new_n992), .ZN(G72));
  AND2_X1   g807(.A1(new_n534), .A2(new_n518), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n994), .A2(new_n529), .ZN(new_n995));
  AOI211_X1 g809(.A(new_n818), .B(new_n976), .C1(new_n981), .C2(new_n982), .ZN(new_n996));
  NAND2_X1  g810(.A1(G472), .A2(G902), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n997), .B(KEYINPUT63), .Z(new_n998));
  XOR2_X1   g812(.A(new_n998), .B(KEYINPUT126), .Z(new_n999));
  OAI21_X1  g813(.A(new_n995), .B1(new_n996), .B2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n1000), .B(KEYINPUT127), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n837), .A2(new_n843), .ZN(new_n1002));
  INV_X1    g816(.A(new_n535), .ZN(new_n1003));
  OAI211_X1 g817(.A(new_n1002), .B(new_n998), .C1(new_n1003), .C2(new_n544), .ZN(new_n1004));
  AND2_X1   g818(.A1(new_n970), .A2(new_n823), .ZN(new_n1005));
  OR2_X1    g819(.A1(new_n1005), .A2(new_n999), .ZN(new_n1006));
  AND2_X1   g820(.A1(new_n994), .A2(new_n529), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n912), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  AND3_X1   g822(.A1(new_n1001), .A2(new_n1004), .A3(new_n1008), .ZN(G57));
endmodule


