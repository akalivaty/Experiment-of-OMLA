//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 0 1 0 0 0 1 1 1 0 1 1 1 0 1 0 1 0 1 0 0 1 0 1 1 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:27 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1221, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1271;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT0), .Z(new_n212));
  INV_X1    g0012(.A(G68), .ZN(new_n213));
  INV_X1    g0013(.A(G238), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G87), .ZN(new_n216));
  INV_X1    g0016(.A(G250), .ZN(new_n217));
  INV_X1    g0017(.A(G257), .ZN(new_n218));
  OAI22_X1  g0018(.A1(new_n216), .A2(new_n217), .B1(new_n202), .B2(new_n218), .ZN(new_n219));
  AOI211_X1 g0019(.A(new_n215), .B(new_n219), .C1(G107), .C2(G264), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G116), .A2(G270), .ZN(new_n221));
  AND2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G50), .ZN(new_n223));
  INV_X1    g0023(.A(G226), .ZN(new_n224));
  INV_X1    g0024(.A(G77), .ZN(new_n225));
  INV_X1    g0025(.A(G244), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  AND2_X1   g0027(.A1(G58), .A2(G232), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n209), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT1), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(KEYINPUT64), .ZN(new_n232));
  INV_X1    g0032(.A(KEYINPUT64), .ZN(new_n233));
  NAND3_X1  g0033(.A1(new_n233), .A2(G1), .A3(G13), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n207), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  NOR2_X1   g0035(.A1(G58), .A2(G68), .ZN(new_n236));
  INV_X1    g0036(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g0037(.A1(new_n237), .A2(G50), .ZN(new_n238));
  INV_X1    g0038(.A(new_n238), .ZN(new_n239));
  AOI211_X1 g0039(.A(new_n212), .B(new_n230), .C1(new_n235), .C2(new_n239), .ZN(G361));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G264), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n242), .B(G270), .Z(new_n243));
  XNOR2_X1  g0043(.A(G238), .B(G244), .ZN(new_n244));
  XNOR2_X1  g0044(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G226), .B(G232), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n243), .B(new_n248), .Z(G358));
  XOR2_X1   g0049(.A(G68), .B(G77), .Z(new_n250));
  XNOR2_X1  g0050(.A(G50), .B(G58), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(G97), .B(G107), .Z(new_n253));
  XNOR2_X1  g0053(.A(G87), .B(G116), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n252), .B(new_n255), .ZN(G351));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n232), .A2(new_n234), .A3(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n259), .B1(G1), .B2(new_n207), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(new_n223), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n207), .B1(new_n236), .B2(new_n223), .ZN(new_n262));
  XNOR2_X1  g0062(.A(new_n262), .B(KEYINPUT67), .ZN(new_n263));
  INV_X1    g0063(.A(G150), .ZN(new_n264));
  INV_X1    g0064(.A(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n207), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT8), .ZN(new_n267));
  INV_X1    g0067(.A(G58), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(KEYINPUT66), .A2(G58), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(KEYINPUT66), .A2(G58), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n269), .B1(new_n274), .B2(new_n267), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n207), .A2(G33), .ZN(new_n276));
  OAI221_X1 g0076(.A(new_n263), .B1(new_n264), .B2(new_n266), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n261), .B1(new_n277), .B2(new_n258), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n223), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n278), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT3), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n265), .ZN(new_n285));
  NAND2_X1  g0085(.A1(KEYINPUT3), .A2(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G1698), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G222), .ZN(new_n289));
  INV_X1    g0089(.A(G223), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n287), .B(new_n289), .C1(new_n290), .C2(new_n288), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n232), .A2(new_n234), .B1(G33), .B2(G41), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n291), .B(new_n292), .C1(G77), .C2(new_n287), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n294));
  INV_X1    g0094(.A(G274), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n231), .ZN(new_n298));
  NAND2_X1  g0098(.A1(G33), .A2(G41), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(new_n294), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n293), .B(new_n297), .C1(new_n224), .C2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G169), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n304), .B1(G179), .B2(new_n302), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n283), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT70), .ZN(new_n308));
  OR2_X1    g0108(.A1(new_n308), .A2(KEYINPUT9), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(KEYINPUT9), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n283), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n282), .A2(new_n308), .A3(KEYINPUT9), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT10), .ZN(new_n314));
  INV_X1    g0114(.A(G190), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n302), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n316), .B1(G200), .B2(new_n302), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n313), .A2(new_n314), .A3(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n314), .B1(new_n313), .B2(new_n317), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n307), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n260), .A2(new_n225), .ZN(new_n322));
  XNOR2_X1  g0122(.A(new_n322), .B(KEYINPUT68), .ZN(new_n323));
  NAND2_X1  g0123(.A1(G20), .A2(G77), .ZN(new_n324));
  XNOR2_X1  g0124(.A(KEYINPUT8), .B(G58), .ZN(new_n325));
  XOR2_X1   g0125(.A(KEYINPUT15), .B(G87), .Z(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  OAI221_X1 g0127(.A(new_n324), .B1(new_n266), .B2(new_n325), .C1(new_n327), .C2(new_n276), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n328), .A2(new_n258), .B1(new_n225), .B2(new_n280), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n323), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n288), .A2(G232), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n287), .B(new_n331), .C1(new_n214), .C2(new_n288), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n332), .B(new_n292), .C1(G107), .C2(new_n287), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n333), .B(new_n297), .C1(new_n226), .C2(new_n301), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(new_n303), .ZN(new_n335));
  OR2_X1    g0135(.A1(new_n334), .A2(G179), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n330), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  OR2_X1    g0137(.A1(new_n334), .A2(new_n315), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n334), .A2(G200), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n338), .A2(new_n323), .A3(new_n329), .A4(new_n339), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  OR2_X1    g0141(.A1(new_n341), .A2(KEYINPUT69), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n287), .B1(G232), .B2(new_n288), .ZN(new_n343));
  NOR2_X1   g0143(.A1(G226), .A2(G1698), .ZN(new_n344));
  OAI22_X1  g0144(.A1(new_n343), .A2(new_n344), .B1(new_n265), .B2(new_n202), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(new_n292), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n346), .B(new_n297), .C1(new_n214), .C2(new_n301), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT13), .ZN(new_n348));
  XNOR2_X1  g0148(.A(new_n347), .B(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(KEYINPUT14), .B1(new_n349), .B2(new_n303), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(G179), .ZN(new_n351));
  XNOR2_X1  g0151(.A(new_n347), .B(KEYINPUT13), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT14), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n352), .A2(new_n353), .A3(G169), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n350), .A2(new_n351), .A3(new_n354), .ZN(new_n355));
  OAI22_X1  g0155(.A1(new_n266), .A2(new_n223), .B1(new_n276), .B2(new_n225), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n207), .A2(G68), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n258), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  XNOR2_X1  g0158(.A(new_n358), .B(KEYINPUT11), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(new_n213), .B2(new_n260), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n280), .A2(new_n213), .ZN(new_n361));
  OAI21_X1  g0161(.A(KEYINPUT12), .B1(new_n361), .B2(KEYINPUT71), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(KEYINPUT71), .ZN(new_n363));
  XOR2_X1   g0163(.A(new_n362), .B(new_n363), .Z(new_n364));
  NOR2_X1   g0164(.A1(new_n360), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n355), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n352), .A2(G200), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n349), .A2(G190), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n368), .A2(new_n369), .A3(new_n365), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n341), .A2(KEYINPUT69), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n342), .A2(new_n367), .A3(new_n370), .A4(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n260), .A2(new_n275), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n373), .B1(new_n280), .B2(new_n275), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  AND2_X1   g0175(.A1(KEYINPUT3), .A2(G33), .ZN(new_n376));
  NOR2_X1   g0176(.A1(KEYINPUT3), .A2(G33), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(KEYINPUT7), .B1(new_n378), .B2(new_n207), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n285), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n286), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(G68), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(G159), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n266), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT66), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(new_n268), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n386), .A2(G68), .A3(new_n270), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n237), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n384), .B1(new_n388), .B2(G20), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n382), .A2(KEYINPUT16), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(KEYINPUT72), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT72), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n382), .A2(new_n389), .A3(new_n392), .A4(KEYINPUT16), .ZN(new_n393));
  AND3_X1   g0193(.A1(new_n391), .A2(new_n258), .A3(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n285), .A2(new_n207), .A3(new_n286), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT7), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n213), .B1(new_n397), .B2(new_n380), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT73), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  AOI211_X1 g0201(.A(KEYINPUT73), .B(new_n213), .C1(new_n397), .C2(new_n380), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n401), .A2(new_n389), .A3(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT16), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n375), .B1(new_n394), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n290), .A2(new_n288), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n287), .B(new_n408), .C1(G226), .C2(new_n288), .ZN(new_n409));
  OAI21_X1  g0209(.A(KEYINPUT74), .B1(new_n265), .B2(new_n216), .ZN(new_n410));
  OR3_X1    g0210(.A1(new_n265), .A2(new_n216), .A3(KEYINPUT74), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n296), .B1(new_n412), .B2(new_n292), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT75), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n300), .A2(G232), .A3(new_n294), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n413), .A2(new_n414), .A3(new_n315), .A4(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n412), .A2(new_n292), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n417), .A2(new_n297), .A3(new_n415), .ZN(new_n418));
  INV_X1    g0218(.A(G200), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n413), .A2(new_n315), .A3(new_n415), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n420), .A2(KEYINPUT75), .A3(new_n421), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n407), .A2(KEYINPUT17), .A3(new_n416), .A4(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT17), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n400), .A2(new_n402), .ZN(new_n425));
  AOI21_X1  g0225(.A(KEYINPUT16), .B1(new_n425), .B2(new_n389), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n391), .A2(new_n258), .A3(new_n393), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n416), .B(new_n374), .C1(new_n426), .C2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n422), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n424), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n374), .B1(new_n426), .B2(new_n427), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n418), .A2(G169), .ZN(new_n432));
  INV_X1    g0232(.A(G179), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n432), .B1(new_n433), .B2(new_n418), .ZN(new_n434));
  AND3_X1   g0234(.A1(new_n431), .A2(KEYINPUT18), .A3(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(KEYINPUT18), .B1(new_n431), .B2(new_n434), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n423), .B(new_n430), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  NOR3_X1   g0237(.A1(new_n321), .A2(new_n372), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(G45), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n440), .A2(G1), .ZN(new_n441));
  NOR2_X1   g0241(.A1(KEYINPUT5), .A2(G41), .ZN(new_n442));
  AND2_X1   g0242(.A1(KEYINPUT5), .A2(G41), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n441), .B(G274), .C1(new_n442), .C2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT77), .ZN(new_n445));
  XNOR2_X1  g0245(.A(KEYINPUT5), .B(G41), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT77), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n446), .A2(new_n447), .A3(G274), .A4(new_n441), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n288), .A2(G257), .ZN(new_n450));
  NAND2_X1  g0250(.A1(G264), .A2(G1698), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n450), .B(new_n451), .C1(new_n376), .C2(new_n377), .ZN(new_n452));
  INV_X1    g0252(.A(G303), .ZN(new_n453));
  AND2_X1   g0253(.A1(new_n453), .A2(KEYINPUT79), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n453), .A2(KEYINPUT79), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n292), .B(new_n452), .C1(new_n456), .C2(new_n287), .ZN(new_n457));
  AOI22_X1  g0257(.A1(new_n446), .A2(new_n441), .B1(new_n298), .B2(new_n299), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(G270), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n449), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(G200), .ZN(new_n461));
  INV_X1    g0261(.A(G116), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(G20), .ZN(new_n463));
  NAND2_X1  g0263(.A1(G33), .A2(G283), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n464), .B(new_n207), .C1(G33), .C2(new_n202), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n258), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT20), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n258), .A2(KEYINPUT20), .A3(new_n463), .A4(new_n465), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n232), .A2(new_n234), .A3(new_n279), .A4(new_n257), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n265), .A2(G1), .ZN(new_n471));
  OAI21_X1  g0271(.A(G116), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n279), .A2(new_n462), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n468), .A2(new_n469), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n461), .B(new_n474), .C1(new_n315), .C2(new_n460), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT21), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n460), .A2(G169), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n476), .B1(new_n477), .B2(new_n474), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n468), .A2(new_n469), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n472), .A2(new_n473), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n481), .A2(KEYINPUT21), .A3(G169), .A4(new_n460), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n449), .A2(new_n457), .A3(new_n459), .A4(G179), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n481), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n475), .A2(new_n478), .A3(new_n482), .A4(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT80), .ZN(new_n487));
  XNOR2_X1  g0287(.A(new_n486), .B(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT4), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n489), .A2(G1698), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n490), .B(G244), .C1(new_n377), .C2(new_n376), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n226), .B1(new_n285), .B2(new_n286), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n491), .B(new_n464), .C1(new_n492), .C2(KEYINPUT4), .ZN(new_n493));
  OAI21_X1  g0293(.A(G250), .B1(new_n376), .B2(new_n377), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n288), .B1(new_n494), .B2(KEYINPUT4), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n292), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n458), .A2(G257), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n496), .A2(new_n497), .A3(new_n449), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G200), .ZN(new_n499));
  OAI21_X1  g0299(.A(G107), .B1(new_n379), .B2(new_n381), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n207), .A2(new_n265), .A3(G77), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT6), .ZN(new_n502));
  AND2_X1   g0302(.A1(G97), .A2(G107), .ZN(new_n503));
  NOR2_X1   g0303(.A1(G97), .A2(G107), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n203), .A2(KEYINPUT6), .A3(G97), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n207), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n500), .A2(new_n501), .A3(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n470), .A2(new_n471), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n509), .A2(new_n258), .B1(G97), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n280), .A2(new_n202), .ZN(new_n512));
  XNOR2_X1  g0312(.A(new_n512), .B(KEYINPUT76), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n496), .A2(new_n497), .A3(G190), .A4(new_n449), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n499), .A2(new_n511), .A3(new_n513), .A4(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n498), .A2(new_n303), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n510), .A2(G97), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n203), .B1(new_n397), .B2(new_n380), .ZN(new_n518));
  INV_X1    g0318(.A(new_n501), .ZN(new_n519));
  NOR3_X1   g0319(.A1(new_n518), .A2(new_n519), .A3(new_n507), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n517), .B(new_n513), .C1(new_n520), .C2(new_n259), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n496), .A2(new_n497), .A3(new_n433), .A4(new_n449), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n516), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n441), .A2(new_n295), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n300), .B(new_n524), .C1(G250), .C2(new_n441), .ZN(new_n525));
  NAND2_X1  g0325(.A1(G33), .A2(G116), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n285), .A2(new_n286), .B1(new_n214), .B2(new_n288), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n226), .A2(G1698), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n292), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n525), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(G200), .ZN(new_n533));
  OAI211_X1 g0333(.A(G190), .B(new_n525), .C1(new_n530), .C2(new_n531), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT19), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(new_n276), .B2(new_n202), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n207), .B(G68), .C1(new_n376), .C2(new_n377), .ZN(new_n537));
  OR2_X1    g0337(.A1(KEYINPUT78), .A2(G87), .ZN(new_n538));
  NAND2_X1  g0338(.A1(KEYINPUT78), .A2(G87), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n204), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n541), .A2(new_n207), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n536), .B(new_n537), .C1(new_n540), .C2(new_n542), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n543), .A2(new_n258), .B1(new_n280), .B2(new_n327), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n510), .A2(G87), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n533), .A2(new_n534), .A3(new_n544), .A4(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n515), .A2(new_n523), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n543), .A2(new_n258), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n327), .A2(new_n280), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n510), .A2(new_n326), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  OAI221_X1 g0351(.A(new_n529), .B1(G238), .B2(G1698), .C1(new_n376), .C2(new_n377), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n292), .B1(new_n553), .B2(new_n527), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n554), .A2(new_n433), .A3(new_n525), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n532), .A2(new_n303), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n551), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n547), .A2(new_n558), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n207), .B(G87), .C1(new_n376), .C2(new_n377), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(KEYINPUT22), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT22), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n287), .A2(new_n562), .A3(new_n207), .A4(G87), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(KEYINPUT81), .B1(new_n207), .B2(G107), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT23), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n207), .A2(G33), .A3(G116), .ZN(new_n568));
  OAI211_X1 g0368(.A(KEYINPUT81), .B(KEYINPUT23), .C1(new_n207), .C2(G107), .ZN(new_n569));
  AND3_X1   g0369(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n564), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(KEYINPUT24), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT24), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n564), .A2(new_n573), .A3(new_n570), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n575), .A2(new_n258), .B1(G107), .B2(new_n510), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n217), .A2(new_n288), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n218), .A2(G1698), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n577), .B(new_n578), .C1(new_n376), .C2(new_n377), .ZN(new_n579));
  NAND2_X1  g0379(.A1(G33), .A2(G294), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n292), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n458), .A2(G264), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n449), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n419), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n585), .A2(KEYINPUT83), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(G13), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n588), .A2(G1), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n589), .A2(G20), .A3(new_n203), .ZN(new_n590));
  XOR2_X1   g0390(.A(new_n590), .B(KEYINPUT25), .Z(new_n591));
  AOI22_X1  g0391(.A1(new_n292), .A2(new_n581), .B1(new_n458), .B2(G264), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n592), .A2(new_n315), .A3(new_n449), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n585), .A2(KEYINPUT83), .A3(new_n593), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n576), .A2(new_n587), .A3(new_n591), .A4(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT84), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n584), .A2(G169), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(KEYINPUT82), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n592), .A2(G179), .A3(new_n449), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT82), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n584), .A2(new_n600), .A3(G169), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n598), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  AND3_X1   g0402(.A1(new_n564), .A2(new_n573), .A3(new_n570), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n573), .B1(new_n564), .B2(new_n570), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n258), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n510), .A2(G107), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n605), .A2(new_n606), .A3(new_n591), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n602), .A2(new_n607), .ZN(new_n608));
  AND3_X1   g0408(.A1(new_n595), .A2(new_n596), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n596), .B1(new_n595), .B2(new_n608), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n488), .B(new_n559), .C1(new_n609), .C2(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n439), .A2(new_n611), .ZN(G372));
  NAND2_X1  g0412(.A1(new_n367), .A2(new_n337), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n423), .A2(new_n430), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n613), .A2(new_n614), .A3(new_n370), .ZN(new_n615));
  INV_X1    g0415(.A(new_n436), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n431), .A2(KEYINPUT18), .A3(new_n434), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  OR2_X1    g0419(.A1(new_n319), .A2(new_n320), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n306), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n478), .A2(new_n482), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n608), .A2(new_n622), .A3(new_n485), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n515), .A2(new_n523), .A3(new_n546), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n623), .A2(new_n624), .A3(new_n595), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n516), .A2(new_n521), .A3(new_n522), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n546), .A2(new_n557), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n626), .A2(KEYINPUT26), .A3(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT26), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n546), .A2(new_n557), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n629), .B1(new_n523), .B2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n628), .A2(KEYINPUT85), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(KEYINPUT26), .B1(new_n626), .B2(new_n627), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT85), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n625), .A2(new_n632), .A3(new_n635), .A4(new_n557), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n438), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n621), .A2(new_n637), .ZN(G369));
  NAND3_X1  g0438(.A1(new_n478), .A2(new_n482), .A3(new_n485), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n589), .A2(new_n207), .ZN(new_n640));
  OR2_X1    g0440(.A1(new_n640), .A2(KEYINPUT27), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(KEYINPUT27), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n641), .A2(new_n642), .A3(G213), .ZN(new_n643));
  INV_X1    g0443(.A(G343), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n646), .A2(new_n474), .ZN(new_n647));
  XNOR2_X1  g0447(.A(new_n647), .B(KEYINPUT86), .ZN(new_n648));
  MUX2_X1   g0448(.A(new_n639), .B(new_n488), .S(new_n648), .Z(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(G330), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n608), .A2(new_n646), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n595), .A2(new_n608), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(KEYINPUT84), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n595), .A2(new_n596), .A3(new_n608), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n607), .A2(new_n645), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n651), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n650), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n639), .A2(new_n646), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n655), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n602), .A2(new_n607), .A3(new_n646), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n658), .A2(new_n663), .ZN(G399));
  INV_X1    g0464(.A(new_n210), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n665), .A2(G41), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n540), .A2(new_n462), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n667), .A2(G1), .A3(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n670), .B1(new_n238), .B2(new_n667), .ZN(new_n671));
  XNOR2_X1  g0471(.A(new_n671), .B(KEYINPUT87), .ZN(new_n672));
  XNOR2_X1  g0472(.A(new_n672), .B(KEYINPUT28), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n636), .A2(new_n646), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT90), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n636), .A2(KEYINPUT90), .A3(new_n646), .ZN(new_n677));
  AOI21_X1  g0477(.A(KEYINPUT29), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n639), .B1(new_n607), .B2(new_n602), .ZN(new_n680));
  INV_X1    g0480(.A(new_n594), .ZN(new_n681));
  NOR3_X1   g0481(.A1(new_n607), .A2(new_n681), .A3(new_n586), .ZN(new_n682));
  NOR3_X1   g0482(.A1(new_n680), .A2(new_n682), .A3(new_n547), .ZN(new_n683));
  NOR3_X1   g0483(.A1(new_n523), .A2(new_n630), .A3(new_n629), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n557), .B1(new_n633), .B2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n646), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(KEYINPUT91), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n558), .B1(new_n628), .B2(new_n631), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n645), .B1(new_n625), .B2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT91), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  AND3_X1   g0491(.A1(new_n687), .A2(KEYINPUT29), .A3(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT89), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n460), .A2(new_n433), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n695), .A2(new_n498), .A3(new_n532), .A4(new_n584), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT30), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n592), .A2(new_n554), .A3(new_n525), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n498), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n697), .B1(new_n699), .B2(new_n484), .ZN(new_n700));
  NOR4_X1   g0500(.A1(new_n498), .A2(new_n698), .A3(new_n483), .A4(KEYINPUT30), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n696), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n646), .B1(new_n702), .B2(KEYINPUT88), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT88), .ZN(new_n704));
  OAI211_X1 g0504(.A(new_n704), .B(new_n696), .C1(new_n700), .C2(new_n701), .ZN(new_n705));
  AOI21_X1  g0505(.A(KEYINPUT31), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n582), .A2(new_n583), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(new_n532), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n217), .B1(new_n285), .B2(new_n286), .ZN(new_n709));
  OAI21_X1  g0509(.A(G1698), .B1(new_n709), .B2(new_n489), .ZN(new_n710));
  OAI21_X1  g0510(.A(G244), .B1(new_n376), .B2(new_n377), .ZN(new_n711));
  AOI22_X1  g0511(.A1(new_n711), .A2(new_n489), .B1(G33), .B2(G283), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n710), .A2(new_n712), .A3(new_n491), .ZN(new_n713));
  AOI22_X1  g0513(.A1(new_n713), .A2(new_n292), .B1(new_n448), .B2(new_n445), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n484), .A2(new_n708), .A3(new_n714), .A4(new_n497), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(KEYINPUT30), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n699), .A2(new_n697), .A3(new_n484), .ZN(new_n717));
  AND3_X1   g0517(.A1(new_n695), .A2(new_n532), .A3(new_n498), .ZN(new_n718));
  AOI22_X1  g0518(.A1(new_n716), .A2(new_n717), .B1(new_n718), .B2(new_n584), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT31), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n719), .A2(new_n720), .A3(new_n646), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n694), .B1(new_n706), .B2(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n645), .B1(new_n719), .B2(new_n704), .ZN(new_n723));
  INV_X1    g0523(.A(new_n705), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n720), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n721), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n725), .A2(KEYINPUT89), .A3(new_n726), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n655), .A2(new_n559), .A3(new_n488), .A4(new_n646), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n722), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(G330), .ZN(new_n730));
  AND3_X1   g0530(.A1(new_n679), .A2(new_n693), .A3(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n673), .B1(new_n731), .B2(G1), .ZN(G364));
  NOR2_X1   g0532(.A1(G13), .A2(G33), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(G20), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  OR2_X1    g0536(.A1(new_n649), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n210), .A2(new_n378), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n738), .B1(new_n440), .B2(new_n239), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n739), .B1(new_n252), .B2(new_n440), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n210), .A2(G355), .A3(new_n287), .ZN(new_n741));
  OAI211_X1 g0541(.A(new_n740), .B(new_n741), .C1(G116), .C2(new_n210), .ZN(new_n742));
  AOI22_X1  g0542(.A1(new_n232), .A2(new_n234), .B1(G20), .B2(new_n303), .ZN(new_n743));
  XOR2_X1   g0543(.A(new_n743), .B(KEYINPUT93), .Z(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n735), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n742), .A2(new_n746), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n588), .A2(new_n440), .A3(G20), .ZN(new_n748));
  OR2_X1    g0548(.A1(new_n748), .A2(KEYINPUT92), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(KEYINPUT92), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n749), .A2(G1), .A3(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n666), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n207), .A2(new_n433), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n315), .A2(new_n419), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n287), .B1(new_n756), .B2(G326), .ZN(new_n757));
  INV_X1    g0557(.A(G294), .ZN(new_n758));
  NOR3_X1   g0558(.A1(new_n315), .A2(G179), .A3(G200), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n207), .ZN(new_n760));
  XOR2_X1   g0560(.A(KEYINPUT33), .B(G317), .Z(new_n761));
  NOR2_X1   g0561(.A1(new_n419), .A2(G190), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n753), .A2(new_n762), .ZN(new_n763));
  OAI221_X1 g0563(.A(new_n757), .B1(new_n758), .B2(new_n760), .C1(new_n761), .C2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n207), .A2(G179), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(new_n762), .ZN(new_n766));
  XNOR2_X1  g0566(.A(new_n766), .B(KEYINPUT95), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n764), .B1(G283), .B2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n753), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n769), .A2(new_n315), .A3(G200), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G190), .A2(G200), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n765), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI22_X1  g0573(.A1(new_n770), .A2(G322), .B1(G329), .B2(new_n773), .ZN(new_n774));
  AND2_X1   g0574(.A1(new_n768), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n754), .A2(new_n765), .ZN(new_n776));
  INV_X1    g0576(.A(G311), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n753), .A2(new_n771), .ZN(new_n778));
  OAI221_X1 g0578(.A(new_n775), .B1(new_n453), .B2(new_n776), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n778), .ZN(new_n780));
  AOI22_X1  g0580(.A1(G50), .A2(new_n756), .B1(new_n780), .B2(G77), .ZN(new_n781));
  INV_X1    g0581(.A(new_n770), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n781), .B1(new_n274), .B2(new_n782), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT94), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n772), .A2(new_n383), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT32), .ZN(new_n786));
  INV_X1    g0586(.A(new_n763), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G68), .ZN(new_n788));
  INV_X1    g0588(.A(new_n760), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G97), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n784), .A2(new_n786), .A3(new_n788), .A4(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n378), .B1(new_n767), .B2(G107), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n538), .A2(new_n539), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n792), .B1(new_n793), .B2(new_n776), .ZN(new_n794));
  XOR2_X1   g0594(.A(new_n794), .B(KEYINPUT96), .Z(new_n795));
  OAI21_X1  g0595(.A(new_n779), .B1(new_n791), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(new_n745), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n737), .A2(new_n747), .A3(new_n752), .A4(new_n797), .ZN(new_n798));
  OR2_X1    g0598(.A1(new_n649), .A2(G330), .ZN(new_n799));
  INV_X1    g0599(.A(new_n752), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n799), .A2(new_n650), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n798), .A2(new_n801), .ZN(G396));
  NAND2_X1  g0602(.A1(new_n330), .A2(new_n645), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n337), .A2(new_n340), .A3(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(KEYINPUT99), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n337), .A2(new_n803), .A3(KEYINPUT99), .A4(new_n340), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n337), .A2(new_n646), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(new_n733), .ZN(new_n811));
  XNOR2_X1  g0611(.A(KEYINPUT98), .B(G143), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n770), .A2(new_n812), .B1(new_n780), .B2(G159), .ZN(new_n813));
  INV_X1    g0613(.A(G137), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n813), .B1(new_n814), .B2(new_n755), .C1(new_n264), .C2(new_n763), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(KEYINPUT34), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n767), .A2(G68), .B1(new_n273), .B2(new_n789), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n378), .B1(new_n773), .B2(G132), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n776), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n819), .B1(G50), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n776), .A2(new_n203), .ZN(new_n822));
  INV_X1    g0622(.A(G283), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n782), .A2(new_n758), .B1(new_n763), .B2(new_n823), .ZN(new_n824));
  AOI211_X1 g0624(.A(new_n822), .B(new_n824), .C1(G116), .C2(new_n780), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n767), .A2(G87), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n790), .B1(new_n777), .B2(new_n772), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n287), .B(new_n827), .C1(G303), .C2(new_n756), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n825), .A2(new_n826), .A3(new_n828), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT97), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n745), .B1(new_n821), .B2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n745), .A2(new_n733), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(new_n225), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n811), .A2(new_n752), .A3(new_n831), .A4(new_n833), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n636), .A2(new_n646), .A3(new_n808), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n676), .A2(new_n677), .ZN(new_n836));
  INV_X1    g0636(.A(new_n810), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n835), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n838), .B(new_n730), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n834), .B1(new_n839), .B2(new_n752), .ZN(G384));
  NAND2_X1  g0640(.A1(new_n505), .A2(new_n506), .ZN(new_n841));
  OAI211_X1 g0641(.A(G116), .B(new_n235), .C1(new_n841), .C2(KEYINPUT35), .ZN(new_n842));
  XOR2_X1   g0642(.A(new_n842), .B(KEYINPUT100), .Z(new_n843));
  NAND2_X1  g0643(.A1(new_n841), .A2(KEYINPUT35), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n845), .B(KEYINPUT36), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n239), .A2(G77), .A3(new_n387), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n847), .B1(G50), .B2(new_n213), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n848), .A2(G1), .A3(new_n588), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT40), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT38), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n236), .B1(new_n273), .B2(G68), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n852), .A2(new_n207), .B1(new_n383), .B2(new_n266), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n405), .B1(new_n853), .B2(new_n398), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n391), .A2(new_n258), .A3(new_n393), .A4(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n374), .ZN(new_n856));
  INV_X1    g0656(.A(new_n643), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n858), .B1(new_n614), .B2(new_n618), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n856), .A2(new_n434), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n858), .B(new_n860), .C1(new_n428), .C2(new_n429), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(KEYINPUT37), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n431), .B1(new_n434), .B2(new_n857), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT37), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n863), .B(new_n864), .C1(new_n428), .C2(new_n429), .ZN(new_n865));
  AND2_X1   g0665(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n851), .B1(new_n859), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n858), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n437), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n862), .A2(new_n865), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n869), .A2(KEYINPUT38), .A3(new_n870), .ZN(new_n871));
  AND2_X1   g0671(.A1(new_n867), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n366), .A2(new_n645), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n367), .A2(new_n370), .A3(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n370), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n366), .B(new_n645), .C1(new_n875), .C2(new_n355), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n703), .A2(KEYINPUT31), .A3(new_n705), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n725), .B(new_n878), .C1(new_n611), .C2(new_n645), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n877), .A2(new_n879), .A3(new_n837), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n850), .B1(new_n872), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(KEYINPUT102), .ZN(new_n882));
  AND3_X1   g0682(.A1(new_n877), .A2(new_n879), .A3(new_n837), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n867), .A2(new_n871), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT102), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n885), .A2(new_n886), .A3(new_n850), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n882), .A2(new_n887), .ZN(new_n888));
  AND3_X1   g0688(.A1(new_n869), .A2(KEYINPUT38), .A3(new_n870), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n407), .A2(new_n643), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n437), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n394), .A2(new_n406), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n413), .A2(G179), .A3(new_n415), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n432), .A2(new_n893), .ZN(new_n894));
  AOI22_X1  g0694(.A1(new_n892), .A2(new_n374), .B1(new_n894), .B2(new_n643), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n428), .A2(new_n429), .ZN(new_n896));
  OAI21_X1  g0696(.A(KEYINPUT37), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n865), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT38), .B1(new_n891), .B2(new_n898), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n883), .B(KEYINPUT40), .C1(new_n889), .C2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n888), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n438), .A2(new_n879), .ZN(new_n902));
  XOR2_X1   g0702(.A(new_n901), .B(new_n902), .Z(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(G330), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n438), .B1(new_n678), .B2(new_n692), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n621), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n618), .A2(new_n857), .ZN(new_n909));
  OR2_X1    g0709(.A1(new_n337), .A2(new_n645), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n910), .B(KEYINPUT101), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n835), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n877), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n909), .B1(new_n914), .B2(new_n884), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT39), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n889), .B2(new_n899), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n867), .A2(KEYINPUT39), .A3(new_n871), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n355), .A2(new_n366), .A3(new_n646), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n917), .A2(new_n918), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n915), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n908), .B(new_n922), .ZN(new_n923));
  XOR2_X1   g0723(.A(new_n904), .B(new_n923), .Z(new_n924));
  AOI21_X1  g0724(.A(new_n206), .B1(G13), .B2(new_n207), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n846), .B(new_n849), .C1(new_n924), .C2(new_n925), .ZN(G367));
  OAI22_X1  g0726(.A1(new_n823), .A2(new_n778), .B1(new_n763), .B2(new_n758), .ZN(new_n927));
  AOI211_X1 g0727(.A(new_n287), .B(new_n927), .C1(new_n456), .C2(new_n770), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n756), .A2(G311), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n820), .A2(G116), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT46), .ZN(new_n931));
  INV_X1    g0731(.A(G317), .ZN(new_n932));
  OAI22_X1  g0732(.A1(new_n766), .A2(new_n202), .B1(new_n772), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n933), .B1(G107), .B2(new_n789), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n928), .A2(new_n929), .A3(new_n931), .A4(new_n934), .ZN(new_n935));
  OAI22_X1  g0735(.A1(new_n274), .A2(new_n776), .B1(new_n814), .B2(new_n772), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(KEYINPUT108), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n287), .B1(new_n766), .B2(new_n225), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n938), .A2(KEYINPUT107), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n938), .A2(KEYINPUT107), .ZN(new_n940));
  OAI22_X1  g0740(.A1(new_n760), .A2(new_n213), .B1(new_n778), .B2(new_n223), .ZN(new_n941));
  NOR4_X1   g0741(.A1(new_n937), .A2(new_n939), .A3(new_n940), .A4(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n756), .A2(new_n812), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n942), .B(new_n943), .C1(new_n383), .C2(new_n763), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n782), .A2(new_n264), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n935), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT109), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT47), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n745), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n544), .A2(new_n545), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n645), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n951), .A2(new_n557), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT103), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n627), .A2(KEYINPUT104), .A3(new_n951), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT104), .ZN(new_n955));
  INV_X1    g0755(.A(new_n951), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n955), .B1(new_n630), .B2(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n953), .A2(new_n954), .A3(new_n957), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n958), .A2(new_n736), .ZN(new_n959));
  OAI221_X1 g0759(.A(new_n746), .B1(new_n210), .B2(new_n327), .C1(new_n243), .C2(new_n738), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n949), .A2(new_n752), .A3(new_n959), .A4(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n521), .A2(new_n645), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n515), .A2(new_n523), .A3(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n523), .B2(new_n646), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n663), .A2(new_n965), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n966), .B(KEYINPUT44), .Z(new_n967));
  NOR2_X1   g0767(.A1(new_n663), .A2(new_n965), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT45), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(new_n658), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT105), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n650), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n657), .A2(new_n659), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n973), .A2(new_n661), .A3(new_n974), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n650), .A2(new_n972), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n975), .B(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n731), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n971), .A2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT106), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n979), .B(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n731), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n666), .B(KEYINPUT41), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n751), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n655), .A2(new_n523), .A3(new_n515), .A4(new_n660), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n985), .B(KEYINPUT42), .Z(new_n986));
  OAI21_X1  g0786(.A(new_n523), .B1(new_n963), .B2(new_n608), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n646), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n986), .A2(new_n988), .B1(KEYINPUT43), .B2(new_n958), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n658), .A2(new_n964), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n989), .B(new_n990), .Z(new_n991));
  NOR2_X1   g0791(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n991), .B(new_n992), .Z(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n961), .B1(new_n984), .B2(new_n994), .ZN(G387));
  OR2_X1    g0795(.A1(new_n977), .A2(new_n731), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n996), .A2(new_n666), .A3(new_n978), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n657), .A2(new_n735), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n325), .A2(G50), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT50), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n668), .B1(G68), .B2(G77), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n1000), .A2(new_n1001), .A3(new_n440), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n738), .B1(new_n248), .B2(G45), .ZN(new_n1003));
  NOR3_X1   g0803(.A1(new_n669), .A2(new_n665), .A3(new_n378), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1002), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n665), .A2(new_n203), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n735), .B(new_n745), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n770), .A2(G50), .B1(new_n756), .B2(G159), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1008), .B1(new_n225), .B2(new_n776), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n327), .A2(new_n760), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n287), .B1(new_n778), .B2(new_n213), .ZN(new_n1011));
  NOR3_X1   g0811(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n767), .A2(G97), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n275), .A2(new_n763), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n773), .A2(G150), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .A4(new_n1015), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n456), .A2(new_n780), .B1(new_n787), .B2(G311), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n756), .A2(G322), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1017), .B(new_n1018), .C1(new_n932), .C2(new_n782), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT48), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1020), .B1(new_n823), .B2(new_n760), .C1(new_n758), .C2(new_n776), .ZN(new_n1021));
  XOR2_X1   g0821(.A(KEYINPUT110), .B(KEYINPUT49), .Z(new_n1022));
  XNOR2_X1  g0822(.A(new_n1021), .B(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n287), .B1(new_n773), .B2(G326), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n462), .B2(new_n766), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1016), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n800), .B(new_n1007), .C1(new_n1026), .C2(new_n745), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n977), .A2(new_n751), .B1(new_n998), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n997), .A2(new_n1028), .ZN(G393));
  NAND2_X1  g0829(.A1(new_n971), .A2(new_n978), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n981), .A2(new_n666), .A3(new_n1030), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n778), .A2(new_n758), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n770), .A2(G311), .B1(new_n756), .B2(G317), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(KEYINPUT52), .Z(new_n1034));
  NAND2_X1  g0834(.A1(new_n820), .A2(G283), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n767), .A2(G107), .B1(new_n456), .B2(new_n787), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n287), .B1(new_n773), .B2(G322), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n1032), .B(new_n1038), .C1(G116), .C2(new_n789), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n287), .B1(new_n763), .B2(new_n223), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n760), .A2(new_n225), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n1040), .B(new_n1041), .C1(new_n773), .C2(new_n812), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n767), .A2(G87), .B1(G68), .B2(new_n820), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1042), .B(new_n1043), .C1(new_n325), .C2(new_n778), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n770), .A2(G159), .B1(new_n756), .B2(G150), .ZN(new_n1045));
  XOR2_X1   g0845(.A(KEYINPUT111), .B(KEYINPUT51), .Z(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT112), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1045), .B(new_n1047), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1044), .A2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n745), .B1(new_n1039), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n965), .A2(new_n735), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n746), .B1(new_n202), .B2(new_n210), .C1(new_n255), .C2(new_n738), .ZN(new_n1052));
  AND4_X1   g0852(.A1(new_n752), .A2(new_n1050), .A3(new_n1051), .A4(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n971), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1053), .B1(new_n1054), .B2(new_n751), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1031), .A2(new_n1055), .ZN(G390));
  AOI22_X1  g0856(.A1(new_n917), .A2(new_n918), .B1(new_n913), .B2(new_n919), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n810), .B1(new_n687), .B2(new_n691), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n911), .ZN(new_n1059));
  OAI21_X1  g0859(.A(KEYINPUT113), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n689), .A2(new_n690), .ZN(new_n1061));
  AOI211_X1 g0861(.A(KEYINPUT91), .B(new_n645), .C1(new_n625), .C2(new_n688), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n837), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT113), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1063), .A2(new_n1064), .A3(new_n911), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1060), .A2(new_n877), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n899), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n920), .B1(new_n1067), .B2(new_n871), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1057), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n729), .A2(G330), .A3(new_n837), .A4(new_n877), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT114), .ZN(new_n1071));
  AND4_X1   g0871(.A1(new_n1071), .A2(new_n879), .A3(G330), .A4(new_n837), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1069), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n879), .A2(G330), .A3(new_n837), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1077), .A2(KEYINPUT114), .A3(new_n877), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1075), .B1(new_n1069), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(KEYINPUT116), .ZN(new_n1080));
  INV_X1    g0880(.A(G330), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n905), .B(new_n621), .C1(new_n1081), .C2(new_n902), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n729), .A2(G330), .A3(new_n837), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n877), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1077), .A2(new_n877), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n912), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1060), .A2(new_n1065), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1076), .A2(new_n1084), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1089), .A2(new_n1070), .A3(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1082), .B1(new_n1088), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1057), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1078), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT116), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1098), .A2(new_n1099), .A3(new_n1075), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1080), .A2(new_n1093), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT115), .ZN(new_n1102));
  AND4_X1   g0902(.A1(new_n1102), .A2(new_n1098), .A3(new_n1075), .A4(new_n1092), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n1057), .B(new_n1073), .C1(new_n1066), .C2(new_n1068), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1078), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1102), .B1(new_n1106), .B2(new_n1092), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1101), .B(new_n666), .C1(new_n1103), .C2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1106), .A2(new_n751), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n767), .A2(G68), .B1(G97), .B2(new_n780), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1041), .B1(G294), .B2(new_n773), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1110), .B(new_n1111), .C1(new_n216), .C2(new_n776), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n763), .A2(new_n203), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n755), .A2(new_n823), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n378), .B1(new_n782), .B2(new_n462), .ZN(new_n1115));
  NOR4_X1   g0915(.A1(new_n1112), .A2(new_n1113), .A3(new_n1114), .A4(new_n1115), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n776), .A2(new_n264), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT53), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n787), .A2(G137), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n789), .A2(G159), .ZN(new_n1120));
  XOR2_X1   g0920(.A(KEYINPUT54), .B(G143), .Z(new_n1121));
  INV_X1    g0921(.A(new_n766), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n780), .A2(new_n1121), .B1(new_n1122), .B2(G50), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1118), .A2(new_n1119), .A3(new_n1120), .A4(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(G125), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n772), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(G128), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n755), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(G132), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n287), .B1(new_n782), .B2(new_n1129), .ZN(new_n1130));
  NOR4_X1   g0930(.A1(new_n1124), .A2(new_n1126), .A3(new_n1128), .A4(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n745), .B1(new_n1116), .B2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n800), .B1(new_n832), .B2(new_n275), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n1133), .B(KEYINPUT117), .ZN(new_n1134));
  AND2_X1   g0934(.A1(new_n917), .A2(new_n918), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1132), .B(new_n1134), .C1(new_n1135), .C2(new_n734), .ZN(new_n1136));
  AND3_X1   g0936(.A1(new_n1108), .A2(new_n1109), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(G378));
  INV_X1    g0938(.A(KEYINPUT121), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1082), .A2(new_n1139), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1082), .A2(new_n1139), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1140), .B(new_n1142), .C1(new_n1107), .C2(new_n1103), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n886), .B1(new_n885), .B2(new_n850), .ZN(new_n1144));
  AOI211_X1 g0944(.A(KEYINPUT102), .B(KEYINPUT40), .C1(new_n883), .C2(new_n884), .ZN(new_n1145));
  OAI211_X1 g0945(.A(G330), .B(new_n900), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n922), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n888), .A2(G330), .A3(new_n900), .A4(new_n922), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n282), .A2(new_n857), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1150), .B(new_n1151), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n321), .B(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1153), .B(new_n1154), .ZN(new_n1155));
  AND3_X1   g0955(.A1(new_n1148), .A2(new_n1149), .A3(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1155), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1157));
  OR2_X1    g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1143), .A2(KEYINPUT57), .A3(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(new_n666), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(KEYINPUT122), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1143), .A2(new_n1158), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT57), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT122), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1159), .A2(new_n1165), .A3(new_n666), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1161), .A2(new_n1164), .A3(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1155), .A2(new_n733), .ZN(new_n1168));
  INV_X1    g0968(.A(G124), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n265), .B1(new_n772), .B2(new_n1169), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n760), .A2(new_n264), .B1(new_n755), .B2(new_n1125), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n782), .A2(new_n1127), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1171), .B(new_n1172), .C1(new_n820), .C2(new_n1121), .ZN(new_n1173));
  OAI221_X1 g0973(.A(new_n1173), .B1(new_n1129), .B2(new_n763), .C1(new_n814), .C2(new_n778), .ZN(new_n1174));
  AOI211_X1 g0974(.A(G41), .B(new_n1170), .C1(new_n1174), .C2(KEYINPUT59), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n1175), .B1(KEYINPUT59), .B2(new_n1174), .C1(new_n383), .C2(new_n766), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n223), .B1(new_n376), .B2(G41), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n760), .A2(new_n213), .B1(new_n755), .B2(new_n462), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1178), .B(KEYINPUT118), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n274), .A2(new_n766), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n776), .A2(new_n225), .B1(new_n772), .B2(new_n823), .ZN(new_n1181));
  OR4_X1    g0981(.A1(G41), .A2(new_n1180), .A3(new_n1181), .A4(new_n287), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n1179), .B(new_n1182), .C1(G97), .C2(new_n787), .ZN(new_n1183));
  OAI221_X1 g0983(.A(new_n1183), .B1(new_n203), .B2(new_n782), .C1(new_n327), .C2(new_n778), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1184), .B(KEYINPUT58), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1176), .A2(new_n1177), .A3(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1186), .A2(new_n745), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n832), .A2(new_n223), .ZN(new_n1188));
  AND3_X1   g0988(.A1(new_n1168), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n1158), .A2(new_n751), .B1(new_n752), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1167), .A2(new_n1190), .ZN(G375));
  OAI21_X1  g0991(.A(new_n378), .B1(new_n782), .B2(new_n823), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n1010), .B(new_n1192), .C1(G294), .C2(new_n756), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n778), .A2(new_n203), .B1(new_n772), .B2(new_n453), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(new_n767), .B2(G77), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1193), .B(new_n1195), .C1(new_n202), .C2(new_n776), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(G116), .B2(new_n787), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n755), .A2(new_n1129), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(new_n1198), .B(KEYINPUT123), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1180), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n780), .A2(G150), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n787), .A2(new_n1121), .B1(new_n773), .B2(G128), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .A4(new_n1202), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n760), .A2(new_n223), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n776), .A2(new_n383), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n287), .B1(new_n782), .B2(new_n814), .ZN(new_n1206));
  NOR4_X1   g1006(.A1(new_n1203), .A2(new_n1204), .A3(new_n1205), .A4(new_n1206), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n745), .B1(new_n1197), .B2(new_n1207), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n752), .B(new_n1208), .C1(new_n877), .C2(new_n734), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(new_n213), .B2(new_n832), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1088), .A2(new_n1091), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1210), .B1(new_n1211), .B2(new_n751), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1088), .A2(new_n1082), .A3(new_n1091), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(new_n983), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1212), .B1(new_n1214), .B2(new_n1092), .ZN(G381));
  NOR2_X1   g1015(.A1(G375), .A2(G378), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(G393), .A2(G396), .ZN(new_n1217));
  NOR4_X1   g1017(.A1(G387), .A2(G384), .A3(G390), .A4(G381), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  XOR2_X1   g1019(.A(new_n1219), .B(KEYINPUT124), .Z(G407));
  NAND2_X1  g1020(.A1(new_n1216), .A2(new_n644), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(G407), .A2(G213), .A3(new_n1221), .ZN(G409));
  INV_X1    g1022(.A(KEYINPUT61), .ZN(new_n1223));
  AND2_X1   g1023(.A1(new_n644), .A2(G213), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1167), .A2(G378), .A3(new_n1190), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1143), .A2(new_n983), .A3(new_n1158), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1190), .A2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT125), .ZN(new_n1228));
  AND3_X1   g1028(.A1(new_n1227), .A2(new_n1137), .A3(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1228), .B1(new_n1227), .B2(new_n1137), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1224), .B1(new_n1225), .B2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1213), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n667), .B1(new_n1233), .B2(KEYINPUT60), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1234), .B(new_n1093), .C1(KEYINPUT60), .C2(new_n1233), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(new_n1212), .ZN(new_n1236));
  XNOR2_X1  g1036(.A(new_n1236), .B(G384), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1224), .A2(G2897), .ZN(new_n1238));
  XNOR2_X1  g1038(.A(new_n1237), .B(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1223), .B1(new_n1232), .B2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(KEYINPUT127), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT127), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1242), .B(new_n1223), .C1(new_n1232), .C2(new_n1239), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1232), .A2(new_n1237), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(KEYINPUT62), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT62), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1232), .A2(new_n1246), .A3(new_n1237), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1241), .A2(new_n1243), .A3(new_n1245), .A4(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(G387), .A2(new_n1055), .A3(new_n1031), .ZN(new_n1249));
  OAI211_X1 g1049(.A(G390), .B(new_n961), .C1(new_n984), .C2(new_n994), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(KEYINPUT126), .ZN(new_n1252));
  XOR2_X1   g1052(.A(G393), .B(G396), .Z(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1252), .A2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1251), .A2(new_n1255), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1252), .A2(new_n1249), .A3(new_n1254), .A4(new_n1250), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1248), .A2(new_n1259), .ZN(new_n1260));
  OAI21_X1  g1060(.A(KEYINPUT63), .B1(new_n1232), .B2(new_n1239), .ZN(new_n1261));
  AOI21_X1  g1061(.A(KEYINPUT61), .B1(new_n1261), .B2(new_n1244), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT63), .ZN(new_n1263));
  OAI211_X1 g1063(.A(new_n1262), .B(new_n1258), .C1(new_n1263), .C2(new_n1244), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1260), .A2(new_n1264), .ZN(G405));
  NAND2_X1  g1065(.A1(G375), .A2(new_n1137), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(new_n1225), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1259), .A2(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1258), .A2(new_n1225), .A3(new_n1266), .ZN(new_n1269));
  AND3_X1   g1069(.A1(new_n1268), .A2(new_n1237), .A3(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1237), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1270), .A2(new_n1271), .ZN(G402));
endmodule


