//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 0 0 1 1 1 0 0 1 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 1 0 1 0 1 1 0 1 0 0 0 0 1 1 0 1 1 0 0 1 0 1 0 1 0 0 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:15 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016;
  INV_X1    g000(.A(KEYINPUT84), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(KEYINPUT64), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT64), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G146), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n189), .A2(new_n191), .A3(G143), .ZN(new_n192));
  INV_X1    g006(.A(G143), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G146), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT1), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G128), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT68), .ZN(new_n199));
  XNOR2_X1  g013(.A(KEYINPUT67), .B(G128), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n200), .B1(new_n192), .B2(KEYINPUT1), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n193), .A2(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n189), .A2(new_n191), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n202), .B1(new_n203), .B2(new_n193), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n199), .B1(new_n201), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(new_n202), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT64), .B(G146), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n206), .B1(new_n207), .B2(G143), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n196), .B1(new_n207), .B2(G143), .ZN(new_n209));
  OAI211_X1 g023(.A(KEYINPUT68), .B(new_n208), .C1(new_n209), .C2(new_n200), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n198), .B1(new_n205), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G101), .ZN(new_n212));
  INV_X1    g026(.A(G107), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G104), .ZN(new_n214));
  INV_X1    g028(.A(G104), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G107), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n212), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(new_n217), .B(KEYINPUT81), .ZN(new_n218));
  OAI21_X1  g032(.A(KEYINPUT3), .B1(new_n215), .B2(G107), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(new_n213), .A3(G104), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n219), .A2(new_n221), .A3(new_n212), .A4(new_n216), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n218), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(KEYINPUT10), .B1(new_n211), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n223), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT10), .ZN(new_n226));
  INV_X1    g040(.A(new_n198), .ZN(new_n227));
  INV_X1    g041(.A(new_n195), .ZN(new_n228));
  INV_X1    g042(.A(G128), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n229), .B1(new_n206), .B2(KEYINPUT1), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n227), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n225), .A2(new_n226), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n224), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n219), .A2(new_n221), .A3(new_n216), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT78), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n219), .A2(new_n221), .A3(KEYINPUT78), .A4(new_n216), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n236), .A2(G101), .A3(new_n237), .ZN(new_n238));
  AND2_X1   g052(.A1(new_n222), .A2(KEYINPUT4), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  AND2_X1   g054(.A1(KEYINPUT0), .A2(G128), .ZN(new_n241));
  NOR2_X1   g055(.A1(KEYINPUT0), .A2(G128), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  AOI22_X1  g057(.A1(new_n228), .A2(new_n241), .B1(new_n208), .B2(new_n243), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT79), .B(KEYINPUT4), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n236), .A2(G101), .A3(new_n237), .A4(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n240), .A2(new_n244), .A3(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT80), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n240), .A2(new_n244), .A3(KEYINPUT80), .A4(new_n246), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G137), .ZN(new_n252));
  OAI21_X1  g066(.A(KEYINPUT11), .B1(new_n252), .B2(G134), .ZN(new_n253));
  INV_X1    g067(.A(G134), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n253), .B1(new_n254), .B2(G137), .ZN(new_n255));
  INV_X1    g069(.A(G131), .ZN(new_n256));
  OR2_X1    g070(.A1(new_n256), .A2(KEYINPUT66), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n252), .A2(KEYINPUT65), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT65), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G137), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n258), .A2(new_n260), .A3(KEYINPUT11), .A4(G134), .ZN(new_n261));
  AND3_X1   g075(.A1(new_n255), .A2(new_n257), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n257), .B1(new_n255), .B2(new_n261), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n233), .A2(new_n251), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT82), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT82), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n233), .A2(new_n251), .A3(new_n267), .A4(new_n264), .ZN(new_n268));
  INV_X1    g082(.A(new_n264), .ZN(new_n269));
  AOI22_X1  g083(.A1(new_n224), .A2(new_n232), .B1(new_n249), .B2(new_n250), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  AOI22_X1  g085(.A1(new_n266), .A2(new_n268), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  XNOR2_X1  g086(.A(G110), .B(G140), .ZN(new_n273));
  INV_X1    g087(.A(G227), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n274), .A2(G953), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n273), .B(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n187), .B1(new_n272), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n271), .A2(new_n269), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n267), .B1(new_n270), .B2(new_n264), .ZN(new_n280));
  AND4_X1   g094(.A1(new_n267), .A2(new_n233), .A3(new_n251), .A4(new_n264), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n282), .A2(KEYINPUT84), .A3(new_n276), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n205), .A2(new_n210), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n227), .ZN(new_n285));
  OAI21_X1  g099(.A(KEYINPUT83), .B1(new_n285), .B2(new_n225), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n225), .A2(new_n231), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT83), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n211), .A2(new_n288), .A3(new_n223), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n286), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n269), .ZN(new_n291));
  OR2_X1    g105(.A1(new_n291), .A2(KEYINPUT12), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n266), .A2(new_n268), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n291), .A2(KEYINPUT12), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n292), .A2(new_n293), .A3(new_n277), .A4(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n278), .A2(new_n283), .A3(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G469), .ZN(new_n297));
  INV_X1    g111(.A(G902), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(G469), .A2(G902), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n276), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n272), .A2(new_n277), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n302), .A2(G469), .A3(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n299), .A2(new_n300), .A3(new_n304), .ZN(new_n305));
  XNOR2_X1  g119(.A(KEYINPUT9), .B(G234), .ZN(new_n306));
  OAI21_X1  g120(.A(G221), .B1(new_n306), .B2(G902), .ZN(new_n307));
  AND2_X1   g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT91), .ZN(new_n309));
  NOR2_X1   g123(.A1(G475), .A2(G902), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G125), .ZN(new_n312));
  INV_X1    g126(.A(G140), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(G125), .A2(G140), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(KEYINPUT16), .ZN(new_n317));
  NOR3_X1   g131(.A1(new_n312), .A2(KEYINPUT16), .A3(G140), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n317), .A2(G146), .A3(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT88), .ZN(new_n321));
  AOI21_X1  g135(.A(KEYINPUT19), .B1(new_n316), .B2(new_n321), .ZN(new_n322));
  AND2_X1   g136(.A1(G125), .A2(G140), .ZN(new_n323));
  NOR2_X1   g137(.A1(G125), .A2(G140), .ZN(new_n324));
  OAI211_X1 g138(.A(new_n321), .B(KEYINPUT19), .C1(new_n323), .C2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n322), .A2(new_n326), .ZN(new_n327));
  OAI211_X1 g141(.A(KEYINPUT89), .B(new_n320), .C1(new_n327), .C2(new_n203), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT89), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n321), .B1(new_n323), .B2(new_n324), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT19), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n203), .B1(new_n332), .B2(new_n325), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT16), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n334), .B1(new_n314), .B2(new_n315), .ZN(new_n335));
  NOR3_X1   g149(.A1(new_n335), .A2(new_n188), .A3(new_n318), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n329), .B1(new_n333), .B2(new_n336), .ZN(new_n337));
  NOR2_X1   g151(.A1(G237), .A2(G953), .ZN(new_n338));
  AND3_X1   g152(.A1(new_n338), .A2(G143), .A3(G214), .ZN(new_n339));
  AOI21_X1  g153(.A(G143), .B1(new_n338), .B2(G214), .ZN(new_n340));
  OAI21_X1  g154(.A(G131), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n338), .A2(G214), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n193), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n338), .A2(G143), .A3(G214), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n343), .A2(new_n256), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n328), .A2(new_n337), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n316), .A2(new_n207), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n348), .B1(new_n188), .B2(new_n316), .ZN(new_n349));
  OAI211_X1 g163(.A(KEYINPUT18), .B(G131), .C1(new_n339), .C2(new_n340), .ZN(new_n350));
  NAND2_X1  g164(.A1(KEYINPUT18), .A2(G131), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n343), .A2(new_n344), .A3(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n349), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n347), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(G113), .B(G122), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n355), .B(new_n215), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(KEYINPUT90), .B1(new_n346), .B2(KEYINPUT17), .ZN(new_n359));
  OAI211_X1 g173(.A(KEYINPUT17), .B(G131), .C1(new_n339), .C2(new_n340), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n188), .B1(new_n335), .B2(new_n318), .ZN(new_n361));
  AND3_X1   g175(.A1(new_n320), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT90), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT17), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n341), .A2(new_n345), .A3(new_n363), .A4(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n359), .A2(new_n362), .A3(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n366), .A2(new_n356), .A3(new_n353), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n311), .B1(new_n358), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT20), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n309), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  AND3_X1   g184(.A1(new_n366), .A2(new_n356), .A3(new_n353), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n356), .B1(new_n347), .B2(new_n353), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n310), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n373), .A2(KEYINPUT91), .A3(KEYINPUT20), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n368), .A2(new_n369), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n370), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n356), .B1(new_n366), .B2(new_n353), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n298), .B1(new_n371), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(G475), .ZN(new_n379));
  AND3_X1   g193(.A1(new_n376), .A2(KEYINPUT92), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(KEYINPUT92), .B1(new_n376), .B2(new_n379), .ZN(new_n381));
  OAI21_X1  g195(.A(G214), .B1(G237), .B2(G902), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  XNOR2_X1  g197(.A(KEYINPUT70), .B(G116), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n384), .A2(KEYINPUT14), .A3(G122), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(G122), .ZN(new_n386));
  INV_X1    g200(.A(G116), .ZN(new_n387));
  OR2_X1    g201(.A1(new_n387), .A2(G122), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  OAI211_X1 g203(.A(G107), .B(new_n385), .C1(new_n389), .C2(KEYINPUT14), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n200), .A2(G143), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n229), .A2(G143), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n391), .A2(new_n254), .A3(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n254), .B1(new_n391), .B2(new_n393), .ZN(new_n396));
  OAI221_X1 g210(.A(new_n390), .B1(G107), .B2(new_n389), .C1(new_n395), .C2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n193), .A2(KEYINPUT13), .A3(G128), .ZN(new_n398));
  XOR2_X1   g212(.A(new_n398), .B(KEYINPUT93), .Z(new_n399));
  OAI21_X1  g213(.A(new_n391), .B1(KEYINPUT13), .B2(new_n392), .ZN(new_n400));
  OAI21_X1  g214(.A(G134), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n213), .B1(new_n386), .B2(new_n388), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n389), .A2(G107), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n401), .B(new_n394), .C1(new_n402), .C2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(G217), .ZN(new_n405));
  NOR3_X1   g219(.A1(new_n306), .A2(new_n405), .A3(G953), .ZN(new_n406));
  AND3_X1   g220(.A1(new_n397), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n406), .B1(new_n397), .B2(new_n404), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(G478), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n410), .A2(KEYINPUT15), .ZN(new_n411));
  NOR3_X1   g225(.A1(new_n409), .A2(G902), .A3(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(G953), .ZN(new_n414));
  AND2_X1   g228(.A1(new_n414), .A2(G952), .ZN(new_n415));
  NAND2_X1  g229(.A1(G234), .A2(G237), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n416), .A2(G902), .A3(G953), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(KEYINPUT21), .B(G898), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n418), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n411), .B1(new_n409), .B2(G902), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n413), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NOR4_X1   g239(.A1(new_n380), .A2(new_n381), .A3(new_n383), .A4(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n244), .A2(G125), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n427), .B1(new_n211), .B2(G125), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n414), .A2(G224), .ZN(new_n429));
  AND2_X1   g243(.A1(new_n429), .A2(KEYINPUT7), .ZN(new_n430));
  OR2_X1    g244(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(KEYINPUT2), .A2(G113), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT69), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n432), .B(new_n433), .ZN(new_n434));
  OR2_X1    g248(.A1(KEYINPUT2), .A2(G113), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n387), .A2(KEYINPUT70), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT70), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(G116), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n437), .A2(new_n439), .A3(G119), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n440), .B1(new_n387), .B2(G119), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n436), .A2(new_n441), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n387), .A2(G119), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n443), .B1(new_n384), .B2(G119), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n444), .A2(new_n435), .A3(new_n434), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n240), .A2(new_n446), .A3(new_n246), .ZN(new_n447));
  XNOR2_X1  g261(.A(G110), .B(G122), .ZN(new_n448));
  XOR2_X1   g262(.A(new_n448), .B(KEYINPUT85), .Z(new_n449));
  INV_X1    g263(.A(KEYINPUT5), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n443), .A2(new_n450), .ZN(new_n451));
  OAI211_X1 g265(.A(G113), .B(new_n451), .C1(new_n441), .C2(new_n450), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n452), .A2(new_n218), .A3(new_n445), .A4(new_n222), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n447), .A2(new_n449), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n452), .A2(new_n445), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n223), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n453), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n449), .B(KEYINPUT8), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n428), .A2(new_n430), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n431), .A2(new_n454), .A3(new_n459), .A4(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n298), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n454), .A2(KEYINPUT6), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n449), .B1(new_n447), .B2(new_n453), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AOI211_X1 g280(.A(KEYINPUT6), .B(new_n449), .C1(new_n447), .C2(new_n453), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n428), .B(new_n429), .ZN(new_n469));
  AOI21_X1  g283(.A(KEYINPUT86), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n465), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n471), .A2(KEYINPUT6), .A3(new_n454), .ZN(new_n472));
  INV_X1    g286(.A(new_n467), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n469), .A2(new_n472), .A3(KEYINPUT86), .A4(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n463), .B1(new_n470), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(G210), .B1(G237), .B2(G902), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n476), .A2(KEYINPUT87), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n476), .A2(new_n478), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT87), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n469), .A2(new_n472), .A3(new_n473), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT86), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n462), .B1(new_n484), .B2(new_n474), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n477), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n480), .A2(new_n481), .A3(new_n486), .ZN(new_n487));
  AND3_X1   g301(.A1(new_n426), .A2(new_n479), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n405), .B1(G234), .B2(new_n298), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n229), .A2(KEYINPUT67), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT67), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(G128), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n491), .A2(new_n493), .A3(G119), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n494), .B1(G119), .B2(new_n229), .ZN(new_n495));
  XNOR2_X1  g309(.A(KEYINPUT24), .B(G110), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n200), .A2(KEYINPUT23), .A3(G119), .ZN(new_n498));
  AOI21_X1  g312(.A(KEYINPUT23), .B1(new_n229), .B2(G119), .ZN(new_n499));
  INV_X1    g313(.A(G119), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n499), .B1(new_n500), .B2(G128), .ZN(new_n501));
  INV_X1    g315(.A(G110), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n498), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n497), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT75), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n497), .A2(new_n503), .A3(KEYINPUT75), .ZN(new_n507));
  AND2_X1   g321(.A1(new_n320), .A2(new_n348), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT76), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n506), .A2(KEYINPUT76), .A3(new_n507), .A4(new_n508), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OR2_X1    g327(.A1(new_n495), .A2(new_n496), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n320), .A2(new_n361), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n498), .A2(new_n501), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(G110), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n514), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n513), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g333(.A(KEYINPUT22), .B(G137), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n414), .A2(G221), .A3(G234), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n520), .B(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n513), .A2(new_n518), .A3(new_n522), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(new_n298), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT25), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n522), .B1(new_n513), .B2(new_n518), .ZN(new_n529));
  INV_X1    g343(.A(new_n518), .ZN(new_n530));
  AOI211_X1 g344(.A(new_n530), .B(new_n523), .C1(new_n511), .C2(new_n512), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n532), .A2(KEYINPUT25), .A3(new_n298), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n490), .B1(new_n528), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n489), .A2(G902), .ZN(new_n535));
  XOR2_X1   g349(.A(new_n535), .B(KEYINPUT77), .Z(new_n536));
  AOI21_X1  g350(.A(new_n534), .B1(new_n536), .B2(new_n532), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT28), .ZN(new_n539));
  AOI21_X1  g353(.A(G134), .B1(new_n258), .B2(new_n260), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n254), .A2(G137), .ZN(new_n541));
  OAI21_X1  g355(.A(G131), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n255), .A2(new_n261), .A3(new_n256), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n544), .B1(new_n284), .B2(new_n227), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n228), .A2(new_n241), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n208), .A2(new_n243), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n548), .A2(new_n264), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n446), .B1(new_n545), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n244), .B1(new_n263), .B2(new_n262), .ZN(new_n551));
  INV_X1    g365(.A(new_n446), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n551), .B(new_n552), .C1(new_n211), .C2(new_n544), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n539), .B1(new_n550), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n539), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n338), .A2(G210), .ZN(new_n558));
  XOR2_X1   g372(.A(new_n558), .B(KEYINPUT27), .Z(new_n559));
  XNOR2_X1  g373(.A(KEYINPUT26), .B(G101), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n559), .B(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n557), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT71), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n553), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(KEYINPUT30), .B1(new_n545), .B2(new_n549), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT30), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n551), .B(new_n567), .C1(new_n211), .C2(new_n544), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n565), .B1(new_n569), .B2(new_n446), .ZN(new_n570));
  AOI211_X1 g384(.A(new_n564), .B(new_n552), .C1(new_n566), .C2(new_n568), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n562), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT31), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OAI211_X1 g388(.A(KEYINPUT31), .B(new_n562), .C1(new_n570), .C2(new_n571), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n563), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(G472), .A2(G902), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(KEYINPUT72), .ZN(new_n578));
  OAI21_X1  g392(.A(KEYINPUT32), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n563), .ZN(new_n580));
  INV_X1    g394(.A(new_n575), .ZN(new_n581));
  INV_X1    g395(.A(new_n544), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n285), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n567), .B1(new_n583), .B2(new_n551), .ZN(new_n584));
  INV_X1    g398(.A(new_n568), .ZN(new_n585));
  OAI211_X1 g399(.A(KEYINPUT71), .B(new_n446), .C1(new_n584), .C2(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n552), .B1(new_n566), .B2(new_n568), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n586), .B1(new_n587), .B2(new_n565), .ZN(new_n588));
  AOI21_X1  g402(.A(KEYINPUT31), .B1(new_n588), .B2(new_n562), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n580), .B1(new_n581), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT32), .ZN(new_n591));
  INV_X1    g405(.A(new_n578), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n579), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(G472), .ZN(new_n595));
  OAI21_X1  g409(.A(KEYINPUT74), .B1(new_n554), .B2(new_n556), .ZN(new_n596));
  OR2_X1    g410(.A1(new_n556), .A2(KEYINPUT74), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT29), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n561), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(G902), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n557), .A2(new_n562), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT73), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n557), .A2(KEYINPUT73), .A3(new_n562), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n586), .B(new_n561), .C1(new_n587), .C2(new_n565), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n605), .A2(new_n600), .A3(new_n606), .A4(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n595), .B1(new_n602), .B2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n538), .B1(new_n594), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n308), .A2(new_n488), .A3(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(G101), .ZN(G3));
  OAI21_X1  g427(.A(G472), .B1(new_n576), .B2(G902), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n590), .A2(new_n592), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n616), .A2(new_n538), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n308), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n480), .A2(KEYINPUT94), .A3(new_n486), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT94), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n485), .A2(new_n620), .A3(new_n477), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n619), .A2(new_n382), .A3(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n380), .ZN(new_n623));
  INV_X1    g437(.A(new_n381), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n410), .B(new_n298), .C1(new_n407), .C2(new_n408), .ZN(new_n626));
  NAND2_X1  g440(.A1(G478), .A2(G902), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n409), .B(KEYINPUT33), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n628), .B1(new_n629), .B2(G478), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n625), .A2(new_n630), .ZN(new_n631));
  NOR4_X1   g445(.A1(new_n618), .A2(new_n422), .A3(new_n622), .A4(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(KEYINPUT34), .B(G104), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G6));
  AND3_X1   g448(.A1(new_n619), .A2(new_n382), .A3(new_n621), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n370), .A2(new_n374), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(KEYINPUT95), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT95), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n370), .A2(new_n638), .A3(new_n374), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  AOI22_X1  g454(.A1(new_n640), .A2(new_n375), .B1(G475), .B2(new_n378), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n413), .A2(new_n424), .ZN(new_n642));
  AND3_X1   g456(.A1(new_n641), .A2(new_n423), .A3(new_n642), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n308), .A2(new_n617), .A3(new_n635), .A4(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT35), .B(G107), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G9));
  INV_X1    g460(.A(KEYINPUT96), .ZN(new_n647));
  OR2_X1    g461(.A1(new_n523), .A2(KEYINPUT36), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n519), .B(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n536), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n647), .B1(new_n534), .B2(new_n651), .ZN(new_n652));
  AOI21_X1  g466(.A(KEYINPUT25), .B1(new_n532), .B2(new_n298), .ZN(new_n653));
  NOR4_X1   g467(.A1(new_n529), .A2(new_n531), .A3(new_n527), .A4(G902), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n489), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n651), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n655), .A2(new_n656), .A3(KEYINPUT96), .ZN(new_n657));
  AND4_X1   g471(.A1(new_n615), .A2(new_n614), .A3(new_n652), .A4(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n308), .A2(new_n488), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT37), .B(G110), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G12));
  AOI21_X1  g475(.A(new_n591), .B1(new_n590), .B2(new_n592), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n576), .A2(KEYINPUT32), .A3(new_n578), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n610), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n652), .A2(new_n657), .ZN(new_n665));
  AND3_X1   g479(.A1(new_n664), .A2(new_n635), .A3(new_n665), .ZN(new_n666));
  OR2_X1    g480(.A1(new_n419), .A2(G900), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n417), .ZN(new_n668));
  AND3_X1   g482(.A1(new_n641), .A2(new_n642), .A3(new_n668), .ZN(new_n669));
  AND3_X1   g483(.A1(new_n669), .A2(new_n307), .A3(new_n305), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n666), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G128), .ZN(G30));
  NAND2_X1  g486(.A1(new_n487), .A2(new_n479), .ZN(new_n673));
  XOR2_X1   g487(.A(new_n673), .B(KEYINPUT38), .Z(new_n674));
  INV_X1    g488(.A(new_n588), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n562), .ZN(new_n676));
  AND2_X1   g490(.A1(new_n550), .A2(new_n553), .ZN(new_n677));
  AOI21_X1  g491(.A(G902), .B1(new_n677), .B2(new_n561), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n595), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n679), .B1(new_n579), .B2(new_n593), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n625), .A2(new_n642), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n655), .A2(new_n656), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n682), .A2(new_n383), .A3(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n674), .A2(new_n681), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n668), .B(KEYINPUT39), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n308), .A2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT97), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n685), .B1(new_n689), .B2(KEYINPUT40), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n690), .B1(KEYINPUT40), .B2(new_n689), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G143), .ZN(G45));
  NAND3_X1  g506(.A1(new_n664), .A2(new_n635), .A3(new_n665), .ZN(new_n693));
  OAI211_X1 g507(.A(new_n630), .B(new_n668), .C1(new_n380), .C2(new_n381), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n305), .A2(new_n695), .A3(new_n307), .ZN(new_n696));
  OAI21_X1  g510(.A(KEYINPUT98), .B1(new_n693), .B2(new_n696), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n305), .A2(new_n307), .A3(new_n695), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n622), .B1(new_n594), .B2(new_n610), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT98), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n698), .A2(new_n699), .A3(new_n700), .A4(new_n665), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n697), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(KEYINPUT99), .B(G146), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G48));
  NAND2_X1  g518(.A1(new_n296), .A2(new_n298), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(G469), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n706), .A2(new_n307), .A3(new_n299), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n707), .A2(new_n622), .ZN(new_n708));
  INV_X1    g522(.A(new_n631), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n708), .A2(new_n709), .A3(new_n611), .A4(new_n423), .ZN(new_n710));
  XNOR2_X1  g524(.A(KEYINPUT41), .B(G113), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G15));
  AND4_X1   g526(.A1(new_n537), .A2(new_n706), .A3(new_n307), .A4(new_n299), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n713), .A2(new_n699), .A3(new_n643), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G116), .ZN(G18));
  OR2_X1    g529(.A1(new_n625), .A2(new_n425), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n716), .A2(new_n707), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n717), .A2(new_n665), .A3(new_n699), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G119), .ZN(G21));
  NOR2_X1   g533(.A1(new_n682), .A2(new_n622), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT101), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n562), .B1(new_n598), .B2(KEYINPUT100), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT100), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n596), .A2(new_n597), .A3(new_n723), .ZN(new_n724));
  AOI22_X1  g538(.A1(new_n722), .A2(new_n724), .B1(new_n574), .B2(new_n575), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n721), .B1(new_n725), .B2(new_n578), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n598), .A2(KEYINPUT100), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n727), .A2(new_n561), .A3(new_n724), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n574), .A2(new_n575), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n730), .A2(KEYINPUT101), .A3(new_n592), .ZN(new_n731));
  AND3_X1   g545(.A1(new_n726), .A2(new_n731), .A3(new_n614), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n713), .A2(new_n423), .A3(new_n720), .A4(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G122), .ZN(G24));
  NAND4_X1  g548(.A1(new_n726), .A2(new_n731), .A3(new_n614), .A4(new_n683), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n735), .A2(new_n694), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n708), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G125), .ZN(G27));
  NAND3_X1  g552(.A1(new_n664), .A2(KEYINPUT103), .A3(new_n537), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT103), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n609), .B1(new_n579), .B2(new_n593), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n740), .B1(new_n741), .B2(new_n538), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n303), .A2(KEYINPUT102), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT102), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n272), .A2(new_n745), .A3(new_n277), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n744), .A2(new_n302), .A3(G469), .A4(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n299), .A2(new_n300), .A3(new_n747), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n748), .A2(new_n307), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n383), .B1(new_n487), .B2(new_n479), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT42), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n694), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n749), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  OAI21_X1  g567(.A(KEYINPUT104), .B1(new_n743), .B2(new_n753), .ZN(new_n754));
  AND3_X1   g568(.A1(new_n750), .A2(new_n748), .A3(new_n307), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n755), .A2(new_n611), .A3(new_n695), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n751), .ZN(new_n757));
  AND4_X1   g571(.A1(new_n307), .A2(new_n752), .A3(new_n750), .A4(new_n748), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT104), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n758), .A2(new_n759), .A3(new_n742), .A4(new_n739), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n754), .A2(new_n757), .A3(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G131), .ZN(G33));
  NAND3_X1  g576(.A1(new_n755), .A2(new_n611), .A3(new_n669), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G134), .ZN(G36));
  INV_X1    g578(.A(new_n307), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n744), .A2(new_n302), .A3(KEYINPUT45), .A4(new_n746), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n302), .A2(new_n303), .ZN(new_n767));
  OAI211_X1 g581(.A(new_n766), .B(G469), .C1(new_n767), .C2(KEYINPUT45), .ZN(new_n768));
  AOI21_X1  g582(.A(KEYINPUT46), .B1(new_n768), .B2(new_n300), .ZN(new_n769));
  INV_X1    g583(.A(new_n299), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n768), .A2(KEYINPUT46), .A3(new_n300), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n765), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n773), .A2(new_n686), .ZN(new_n774));
  INV_X1    g588(.A(new_n750), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n624), .A2(new_n630), .A3(new_n623), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT105), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(KEYINPUT43), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n616), .A2(new_n683), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT44), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n775), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  OAI211_X1 g597(.A(new_n774), .B(new_n783), .C1(new_n782), .C2(new_n781), .ZN(new_n784));
  XNOR2_X1  g598(.A(KEYINPUT106), .B(G137), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n784), .B(new_n785), .ZN(G39));
  NOR4_X1   g600(.A1(new_n775), .A2(new_n664), .A3(new_n537), .A4(new_n694), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n773), .A2(KEYINPUT47), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n773), .A2(KEYINPUT47), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G140), .ZN(G42));
  NOR2_X1   g605(.A1(G952), .A2(G953), .ZN(new_n792));
  AOI22_X1  g606(.A1(new_n666), .A2(new_n670), .B1(new_n736), .B2(new_n708), .ZN(new_n793));
  INV_X1    g607(.A(new_n668), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n683), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n749), .A2(KEYINPUT108), .A3(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n748), .A2(new_n307), .A3(new_n795), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT108), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n680), .A2(new_n682), .A3(new_n622), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n796), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n702), .A2(new_n793), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(KEYINPUT110), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT109), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n803), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n702), .A2(new_n793), .A3(KEYINPUT52), .A4(new_n801), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(new_n804), .ZN(new_n809));
  INV_X1    g623(.A(new_n806), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n802), .A2(KEYINPUT110), .A3(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n807), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  AND4_X1   g626(.A1(new_n710), .A2(new_n718), .A3(new_n733), .A4(new_n714), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT113), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n761), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n308), .B(new_n488), .C1(new_n611), .C2(new_n658), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n673), .A2(new_n383), .A3(new_n422), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n413), .A2(KEYINPUT107), .A3(new_n424), .ZN(new_n818));
  AOI21_X1  g632(.A(KEYINPUT107), .B1(new_n413), .B2(new_n424), .ZN(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n624), .A2(new_n623), .A3(new_n818), .A4(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n631), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n308), .A2(new_n817), .A3(new_n617), .A4(new_n822), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n816), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n794), .B1(new_n820), .B2(new_n818), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n641), .A2(new_n652), .A3(new_n825), .A4(new_n657), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n775), .A2(new_n741), .A3(new_n826), .ZN(new_n827));
  AOI22_X1  g641(.A1(new_n827), .A2(new_n308), .B1(new_n736), .B2(new_n755), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n824), .A2(KEYINPUT112), .A3(new_n763), .A4(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT112), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n736), .A2(new_n755), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n741), .A2(new_n826), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n832), .A2(new_n308), .A3(new_n750), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n763), .A2(new_n831), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n816), .A2(new_n823), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n830), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n829), .A2(new_n836), .A3(KEYINPUT53), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n814), .B1(new_n761), .B2(new_n813), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n812), .A2(new_n815), .A3(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT54), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n834), .A2(new_n835), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n761), .A2(new_n842), .A3(new_n813), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n802), .A2(new_n805), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(new_n808), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT53), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n840), .A2(new_n841), .A3(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(KEYINPUT111), .B1(new_n847), .B2(new_n848), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT111), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n844), .A2(new_n846), .A3(new_n852), .A4(KEYINPUT53), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n802), .A2(KEYINPUT110), .A3(new_n810), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n810), .B1(new_n802), .B2(KEYINPUT110), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n843), .B1(new_n856), .B2(new_n809), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n851), .B(new_n853), .C1(new_n857), .C2(KEYINPUT53), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n850), .B1(KEYINPUT54), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n788), .A2(new_n789), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n706), .A2(new_n299), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n860), .B1(new_n307), .B2(new_n861), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n732), .A2(new_n537), .ZN(new_n863));
  AND4_X1   g677(.A1(new_n418), .A2(new_n779), .A3(new_n750), .A4(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT114), .ZN(new_n866));
  OR3_X1    g680(.A1(new_n674), .A2(new_n382), .A3(new_n707), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n779), .A2(new_n418), .A3(new_n863), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT50), .ZN(new_n870));
  OR2_X1    g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n775), .A2(new_n707), .A3(new_n417), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n681), .A2(new_n538), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n625), .A2(new_n630), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n779), .A2(new_n872), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n875), .B1(new_n876), .B2(new_n735), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n877), .B1(new_n869), .B2(new_n870), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n865), .A2(KEYINPUT51), .A3(new_n871), .A4(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n872), .A2(new_n709), .A3(new_n873), .ZN(new_n880));
  INV_X1    g694(.A(new_n708), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n880), .B(new_n415), .C1(new_n868), .C2(new_n881), .ZN(new_n882));
  OR2_X1    g696(.A1(new_n876), .A2(new_n743), .ZN(new_n883));
  OR2_X1    g697(.A1(new_n883), .A2(KEYINPUT48), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(KEYINPUT48), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n882), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n879), .A2(new_n886), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n871), .A2(new_n878), .ZN(new_n888));
  AOI21_X1  g702(.A(KEYINPUT51), .B1(new_n888), .B2(new_n865), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n792), .B1(new_n859), .B2(new_n890), .ZN(new_n891));
  NOR4_X1   g705(.A1(new_n674), .A2(new_n765), .A3(new_n383), .A4(new_n776), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n861), .A2(KEYINPUT49), .ZN(new_n893));
  OR2_X1    g707(.A1(new_n861), .A2(KEYINPUT49), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n892), .A2(new_n873), .A3(new_n893), .A4(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(KEYINPUT115), .B1(new_n891), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n851), .A2(new_n853), .ZN(new_n898));
  AOI21_X1  g712(.A(KEYINPUT53), .B1(new_n812), .B2(new_n844), .ZN(new_n899));
  OAI21_X1  g713(.A(KEYINPUT54), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(new_n850), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n900), .A2(new_n890), .A3(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n792), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT115), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n904), .A2(new_n905), .A3(new_n895), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n897), .A2(new_n906), .ZN(G75));
  XOR2_X1   g721(.A(new_n469), .B(KEYINPUT117), .Z(new_n908));
  NAND2_X1  g722(.A1(new_n840), .A2(new_n849), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n909), .A2(G210), .A3(G902), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT56), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n468), .B(KEYINPUT116), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(KEYINPUT55), .Z(new_n913));
  AND3_X1   g727(.A1(new_n910), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n913), .B1(new_n910), .B2(new_n911), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n908), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n910), .A2(new_n911), .ZN(new_n917));
  INV_X1    g731(.A(new_n913), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(new_n908), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n910), .A2(new_n911), .A3(new_n913), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n414), .A2(G952), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  AND3_X1   g738(.A1(new_n916), .A2(new_n922), .A3(new_n924), .ZN(G51));
  INV_X1    g739(.A(new_n815), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n926), .A2(new_n837), .A3(new_n838), .ZN(new_n927));
  AOI22_X1  g741(.A1(new_n927), .A2(new_n812), .B1(new_n848), .B2(new_n847), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(new_n841), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n300), .B(KEYINPUT118), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT57), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(new_n296), .ZN(new_n933));
  OR3_X1    g747(.A1(new_n928), .A2(new_n298), .A3(new_n768), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n923), .B1(new_n933), .B2(new_n934), .ZN(G54));
  NAND4_X1  g749(.A1(new_n909), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n371), .A2(new_n372), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n936), .A2(new_n937), .ZN(new_n939));
  NOR3_X1   g753(.A1(new_n938), .A2(new_n939), .A3(new_n923), .ZN(G60));
  XOR2_X1   g754(.A(new_n627), .B(KEYINPUT59), .Z(new_n941));
  NOR2_X1   g755(.A1(new_n629), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n929), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(new_n924), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n629), .B1(new_n859), .B2(new_n941), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT119), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  OAI211_X1 g761(.A(KEYINPUT119), .B(new_n629), .C1(new_n859), .C2(new_n941), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n944), .B1(new_n947), .B2(new_n948), .ZN(G63));
  INV_X1    g763(.A(KEYINPUT61), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT120), .ZN(new_n951));
  NAND2_X1  g765(.A1(G217), .A2(G902), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT60), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n951), .B1(new_n928), .B2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n953), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n909), .A2(KEYINPUT120), .A3(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(new_n532), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n954), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n924), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n649), .B1(new_n954), .B2(new_n956), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n950), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n960), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n962), .A2(new_n958), .A3(KEYINPUT61), .A4(new_n924), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n961), .A2(new_n963), .ZN(G66));
  INV_X1    g778(.A(new_n421), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n414), .B1(new_n965), .B2(G224), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n813), .A2(new_n824), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT121), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n967), .B(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n966), .B1(new_n969), .B2(new_n414), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n912), .B1(G898), .B2(new_n414), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n971), .B(KEYINPUT122), .Z(new_n972));
  XNOR2_X1  g786(.A(new_n970), .B(new_n972), .ZN(G69));
  XNOR2_X1  g787(.A(new_n569), .B(new_n327), .ZN(new_n974));
  INV_X1    g788(.A(new_n974), .ZN(new_n975));
  OAI211_X1 g789(.A(G900), .B(G953), .C1(new_n975), .C2(G227), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n976), .B1(G227), .B2(new_n975), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT123), .ZN(new_n978));
  AND3_X1   g792(.A1(new_n702), .A2(new_n978), .A3(new_n793), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n978), .B1(new_n702), .B2(new_n793), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n691), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT62), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n982), .A2(KEYINPUT62), .A3(new_n691), .ZN(new_n986));
  AND2_X1   g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n611), .A2(new_n750), .A3(new_n822), .ZN(new_n988));
  OAI211_X1 g802(.A(new_n784), .B(new_n790), .C1(new_n689), .C2(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n974), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(new_n763), .ZN(new_n991));
  NOR3_X1   g805(.A1(new_n743), .A2(new_n622), .A3(new_n682), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n991), .B1(new_n774), .B2(new_n992), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n784), .A2(new_n790), .A3(new_n993), .A4(new_n761), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n994), .A2(new_n981), .ZN(new_n995));
  AOI21_X1  g809(.A(G953), .B1(new_n995), .B2(new_n975), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n977), .B1(new_n990), .B2(new_n996), .ZN(G72));
  NOR2_X1   g811(.A1(new_n675), .A2(new_n562), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n998), .B(KEYINPUT124), .Z(new_n999));
  NOR3_X1   g813(.A1(new_n969), .A2(new_n994), .A3(new_n981), .ZN(new_n1000));
  NAND2_X1  g814(.A1(G472), .A2(G902), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n1001), .B(KEYINPUT63), .Z(new_n1002));
  INV_X1    g816(.A(new_n1002), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n999), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT125), .ZN(new_n1005));
  AND3_X1   g819(.A1(new_n1004), .A2(new_n1005), .A3(new_n924), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n1005), .B1(new_n1004), .B2(new_n924), .ZN(new_n1007));
  AOI211_X1 g821(.A(new_n969), .B(new_n989), .C1(new_n985), .C2(new_n986), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n1008), .A2(new_n1003), .ZN(new_n1009));
  OAI22_X1  g823(.A1(new_n1006), .A2(new_n1007), .B1(new_n1009), .B2(new_n676), .ZN(new_n1010));
  INV_X1    g824(.A(new_n998), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n1011), .A2(new_n676), .A3(new_n1002), .ZN(new_n1012));
  XOR2_X1   g826(.A(new_n1012), .B(KEYINPUT126), .Z(new_n1013));
  NAND2_X1  g827(.A1(new_n858), .A2(new_n1013), .ZN(new_n1014));
  OR2_X1    g828(.A1(new_n1014), .A2(KEYINPUT127), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1014), .A2(KEYINPUT127), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1010), .B1(new_n1015), .B2(new_n1016), .ZN(G57));
endmodule


