//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 1 0 1 1 0 0 1 1 1 0 0 1 0 1 0 0 0 0 0 0 1 1 0 1 1 1 0 0 1 0 0 1 1 0 1 1 0 0 1 1 1 1 1 0 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:42 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1265, new_n1266, new_n1267,
    new_n1268, new_n1269, new_n1270, new_n1271, new_n1272, new_n1273,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  XNOR2_X1  g0001(.A(new_n201), .B(KEYINPUT64), .ZN(new_n202));
  INV_X1    g0002(.A(G77), .ZN(new_n203));
  AND2_X1   g0003(.A1(new_n202), .A2(new_n203), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  OR3_X1    g0014(.A1(KEYINPUT65), .A2(G58), .A3(G68), .ZN(new_n215));
  OAI21_X1  g0015(.A(KEYINPUT65), .B1(G58), .B2(G68), .ZN(new_n216));
  NAND3_X1  g0016(.A1(new_n215), .A2(G50), .A3(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n219), .A2(new_n209), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  XOR2_X1   g0021(.A(KEYINPUT66), .B(G238), .Z(new_n222));
  INV_X1    g0022(.A(G68), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G107), .A2(G264), .ZN(new_n228));
  NAND4_X1  g0028(.A1(new_n225), .A2(new_n226), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n211), .B1(new_n224), .B2(new_n229), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n214), .B(new_n221), .C1(KEYINPUT1), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  INV_X1    g0043(.A(G50), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(G68), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n223), .A2(G50), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n243), .B(new_n249), .ZN(G351));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n219), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n202), .A2(new_n209), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT8), .B(G58), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n209), .A2(G33), .ZN(new_n255));
  INV_X1    g0055(.A(G150), .ZN(new_n256));
  NOR2_X1   g0056(.A1(G20), .A2(G33), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  OAI22_X1  g0058(.A1(new_n254), .A2(new_n255), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n252), .B1(new_n253), .B2(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(new_n219), .A3(new_n251), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n244), .B1(new_n208), .B2(G20), .ZN(new_n264));
  INV_X1    g0064(.A(new_n261), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n263), .A2(new_n264), .B1(new_n244), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n260), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g0067(.A(new_n267), .B(KEYINPUT9), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT10), .ZN(new_n269));
  INV_X1    g0069(.A(G41), .ZN(new_n270));
  INV_X1    g0070(.A(G45), .ZN(new_n271));
  AOI21_X1  g0071(.A(G1), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G33), .A2(G41), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n273), .A2(G1), .A3(G13), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n272), .A2(new_n274), .A3(G274), .ZN(new_n275));
  INV_X1    g0075(.A(G226), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n275), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT3), .B(G33), .ZN(new_n280));
  NOR2_X1   g0080(.A1(G222), .A2(G1698), .ZN(new_n281));
  INV_X1    g0081(.A(G1698), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(G223), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n280), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(KEYINPUT3), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT3), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n274), .B1(new_n289), .B2(new_n203), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n279), .B1(new_n284), .B2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G200), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n293), .B1(G190), .B2(new_n291), .ZN(new_n294));
  AND3_X1   g0094(.A1(new_n268), .A2(new_n269), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n269), .B1(new_n268), .B2(new_n294), .ZN(new_n296));
  OR2_X1    g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G179), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n291), .A2(new_n298), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n299), .B(new_n267), .C1(G169), .C2(new_n291), .ZN(new_n300));
  INV_X1    g0100(.A(G244), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n222), .A2(G1698), .ZN(new_n302));
  INV_X1    g0102(.A(G232), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(new_n282), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n289), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n219), .B1(G33), .B2(G41), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n306), .B1(new_n280), .B2(G107), .ZN(new_n307));
  OAI221_X1 g0107(.A(new_n275), .B1(new_n301), .B2(new_n278), .C1(new_n305), .C2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(G200), .ZN(new_n309));
  OAI22_X1  g0109(.A1(new_n254), .A2(new_n258), .B1(new_n209), .B2(new_n203), .ZN(new_n310));
  XNOR2_X1  g0110(.A(KEYINPUT15), .B(G87), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n311), .A2(new_n255), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n252), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n208), .A2(G20), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G77), .ZN(new_n315));
  OAI221_X1 g0115(.A(new_n313), .B1(G77), .B2(new_n261), .C1(new_n262), .C2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G190), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n309), .B(new_n317), .C1(new_n318), .C2(new_n308), .ZN(new_n319));
  INV_X1    g0119(.A(G169), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n317), .B1(new_n308), .B2(new_n320), .ZN(new_n321));
  OR2_X1    g0121(.A1(new_n308), .A2(G179), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n297), .A2(new_n300), .A3(new_n319), .A4(new_n323), .ZN(new_n324));
  OR2_X1    g0124(.A1(new_n324), .A2(KEYINPUT67), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n276), .A2(new_n282), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n303), .A2(G1698), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n280), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(G33), .A2(G97), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n274), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT13), .ZN(new_n332));
  INV_X1    g0132(.A(G238), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n275), .B1(new_n333), .B2(new_n278), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n331), .A2(new_n332), .A3(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(KEYINPUT13), .B1(new_n330), .B2(new_n334), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(KEYINPUT68), .B1(new_n339), .B2(new_n292), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT68), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n338), .A2(new_n341), .A3(G200), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n336), .A2(G190), .A3(new_n337), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n314), .A2(G68), .ZN(new_n345));
  OR3_X1    g0145(.A1(new_n262), .A2(KEYINPUT69), .A3(new_n345), .ZN(new_n346));
  OAI21_X1  g0146(.A(KEYINPUT69), .B1(new_n262), .B2(new_n345), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n257), .A2(G50), .B1(G20), .B2(new_n223), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n349), .B1(new_n203), .B2(new_n255), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n252), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT11), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n265), .A2(new_n223), .ZN(new_n354));
  XNOR2_X1  g0154(.A(new_n354), .B(KEYINPUT12), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n350), .A2(KEYINPUT11), .A3(new_n252), .ZN(new_n356));
  AND4_X1   g0156(.A1(new_n348), .A2(new_n353), .A3(new_n355), .A4(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n344), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(KEYINPUT70), .B1(new_n343), .B2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT70), .ZN(new_n361));
  AOI211_X1 g0161(.A(new_n361), .B(new_n358), .C1(new_n340), .C2(new_n342), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n363), .B1(new_n324), .B2(KEYINPUT67), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT77), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n254), .B1(new_n208), .B2(G20), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n366), .A2(new_n263), .B1(new_n265), .B2(new_n254), .ZN(new_n367));
  OR2_X1    g0167(.A1(G223), .A2(G1698), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n276), .A2(G1698), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n286), .A2(new_n368), .A3(new_n288), .A4(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(G33), .A2(G87), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n274), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n274), .A2(G232), .A3(new_n277), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n275), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(new_n318), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n292), .B1(new_n372), .B2(new_n374), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(KEYINPUT75), .B1(new_n285), .B2(KEYINPUT3), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT74), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(new_n287), .B2(G33), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT75), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n382), .A2(new_n287), .A3(G33), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n285), .A2(KEYINPUT74), .A3(KEYINPUT3), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n379), .A2(new_n381), .A3(new_n383), .A4(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT7), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n386), .A2(G20), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n287), .A2(G33), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n285), .A2(KEYINPUT3), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n209), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n386), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n388), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(G68), .ZN(new_n394));
  XNOR2_X1  g0194(.A(G58), .B(G68), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(G20), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n257), .A2(G159), .ZN(new_n397));
  AND2_X1   g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(KEYINPUT16), .B1(new_n394), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT73), .ZN(new_n400));
  AND3_X1   g0200(.A1(new_n286), .A2(new_n288), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n400), .B1(new_n286), .B2(new_n288), .ZN(new_n402));
  NOR2_X1   g0202(.A1(KEYINPUT7), .A2(G20), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  NOR3_X1   g0204(.A1(new_n401), .A2(new_n402), .A3(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(G20), .B1(new_n286), .B2(new_n288), .ZN(new_n406));
  OAI21_X1  g0206(.A(G68), .B1(new_n406), .B2(new_n386), .ZN(new_n407));
  OAI211_X1 g0207(.A(KEYINPUT16), .B(new_n398), .C1(new_n405), .C2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n252), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n367), .B(new_n378), .C1(new_n399), .C2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT17), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n367), .ZN(new_n413));
  INV_X1    g0213(.A(new_n252), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n396), .A2(new_n397), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n223), .B1(new_n391), .B2(KEYINPUT7), .ZN(new_n416));
  OAI21_X1  g0216(.A(KEYINPUT73), .B1(new_n389), .B2(new_n390), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n286), .A2(new_n288), .A3(new_n400), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n417), .A2(new_n418), .A3(new_n403), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n415), .B1(new_n416), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n414), .B1(new_n420), .B2(KEYINPUT16), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT16), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n223), .B1(new_n388), .B2(new_n392), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n422), .B1(new_n423), .B2(new_n415), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n413), .B1(new_n421), .B2(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(KEYINPUT17), .B1(new_n425), .B2(new_n378), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n365), .B1(new_n412), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT18), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n367), .B1(new_n399), .B2(new_n409), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n375), .A2(new_n298), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n320), .B1(new_n372), .B2(new_n374), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n430), .A2(KEYINPUT76), .A3(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n432), .B1(KEYINPUT76), .B2(new_n430), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n428), .B1(new_n429), .B2(new_n433), .ZN(new_n434));
  NOR4_X1   g0234(.A1(new_n372), .A2(new_n374), .A3(KEYINPUT76), .A4(G179), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT76), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n436), .B1(new_n375), .B2(new_n298), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n435), .B1(new_n437), .B2(new_n431), .ZN(new_n438));
  NOR3_X1   g0238(.A1(new_n425), .A2(new_n438), .A3(KEYINPUT18), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n434), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n410), .A2(new_n411), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n425), .A2(KEYINPUT17), .A3(new_n378), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n441), .A2(KEYINPUT77), .A3(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n427), .A2(new_n440), .A3(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n320), .B1(new_n336), .B2(new_n337), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT14), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n339), .A2(G179), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n338), .A2(G169), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n447), .B1(new_n450), .B2(KEYINPUT71), .ZN(new_n451));
  AOI211_X1 g0251(.A(KEYINPUT71), .B(new_n320), .C1(new_n336), .C2(new_n337), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n451), .A2(KEYINPUT72), .A3(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT72), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT71), .ZN(new_n456));
  OAI21_X1  g0256(.A(KEYINPUT14), .B1(new_n446), .B2(new_n456), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n455), .B1(new_n457), .B2(new_n452), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n449), .B1(new_n454), .B2(new_n458), .ZN(new_n459));
  OR2_X1    g0259(.A1(new_n459), .A2(new_n357), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n325), .A2(new_n364), .A3(new_n445), .A4(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n262), .B1(new_n208), .B2(G33), .ZN(new_n462));
  INV_X1    g0262(.A(new_n311), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT80), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n280), .A2(new_n209), .A3(G68), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT19), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n209), .B1(new_n329), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n468), .B1(G87), .B2(new_n206), .ZN(new_n469));
  INV_X1    g0269(.A(G97), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n467), .B1(new_n255), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n466), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n252), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n463), .A2(new_n261), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n465), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  AOI211_X1 g0276(.A(KEYINPUT80), .B(new_n474), .C1(new_n472), .C2(new_n252), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n464), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT81), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OAI211_X1 g0280(.A(KEYINPUT81), .B(new_n464), .C1(new_n476), .C2(new_n477), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT82), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n480), .A2(KEYINPUT82), .A3(new_n481), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n271), .A2(G1), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n274), .A2(G274), .A3(new_n486), .ZN(new_n487));
  OAI21_X1  g0287(.A(G250), .B1(new_n271), .B2(G1), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n487), .B1(new_n306), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(G33), .A2(G116), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n301), .A2(G1698), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n491), .B1(G238), .B2(G1698), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n490), .B1(new_n492), .B2(new_n289), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n489), .B1(new_n493), .B2(new_n306), .ZN(new_n494));
  OR2_X1    g0294(.A1(new_n494), .A2(new_n320), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(G179), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n484), .A2(new_n485), .A3(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(G87), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n414), .B(new_n261), .C1(G1), .C2(new_n285), .ZN(new_n500));
  OAI22_X1  g0300(.A1(new_n476), .A2(new_n477), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n494), .A2(G190), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n502), .B1(new_n292), .B2(new_n494), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n498), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n280), .A2(new_n209), .A3(G87), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(KEYINPUT22), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT22), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n280), .A2(new_n509), .A3(new_n209), .A4(G87), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT24), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT23), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n513), .B1(new_n209), .B2(G107), .ZN(new_n514));
  INV_X1    g0314(.A(G107), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n515), .A2(KEYINPUT23), .A3(G20), .ZN(new_n516));
  INV_X1    g0316(.A(new_n490), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n514), .A2(new_n516), .B1(new_n517), .B2(new_n209), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n511), .A2(new_n512), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n512), .B1(new_n511), .B2(new_n518), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n252), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(KEYINPUT25), .B1(new_n265), .B2(new_n515), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n265), .A2(KEYINPUT25), .A3(new_n515), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n462), .A2(G107), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n521), .A2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(G274), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n306), .A2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT79), .ZN(new_n529));
  XNOR2_X1  g0329(.A(KEYINPUT5), .B(G41), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n528), .A2(new_n529), .A3(new_n486), .A4(new_n530), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n530), .A2(G274), .A3(new_n274), .A4(new_n486), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(KEYINPUT79), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n306), .B1(new_n486), .B2(new_n530), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G264), .ZN(new_n537));
  MUX2_X1   g0337(.A(G250), .B(G257), .S(G1698), .Z(new_n538));
  AOI22_X1  g0338(.A1(new_n538), .A2(new_n280), .B1(G33), .B2(G294), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n537), .B1(new_n274), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g0340(.A(G169), .B1(new_n535), .B2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(G264), .ZN(new_n542));
  AOI211_X1 g0342(.A(new_n542), .B(new_n306), .C1(new_n486), .C2(new_n530), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n538), .A2(new_n280), .ZN(new_n544));
  NAND2_X1  g0344(.A1(G33), .A2(G294), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n274), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g0346(.A(KEYINPUT84), .B1(new_n543), .B2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT84), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n537), .B(new_n548), .C1(new_n539), .C2(new_n274), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n547), .A2(new_n549), .A3(new_n534), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n541), .B1(new_n550), .B2(new_n298), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n526), .A2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(G303), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n274), .B1(new_n289), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(G257), .A2(G1698), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n282), .A2(G264), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n280), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n536), .A2(G270), .B1(new_n554), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n320), .B1(new_n534), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(G33), .A2(G283), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n560), .B(new_n209), .C1(G33), .C2(new_n470), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n561), .B(new_n252), .C1(new_n209), .C2(G116), .ZN(new_n562));
  XNOR2_X1  g0362(.A(new_n562), .B(KEYINPUT20), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n261), .A2(G116), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(G116), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n565), .B1(new_n500), .B2(new_n566), .ZN(new_n567));
  NOR3_X1   g0367(.A1(new_n563), .A2(KEYINPUT83), .A3(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT83), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT20), .ZN(new_n570));
  XNOR2_X1  g0370(.A(new_n562), .B(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n564), .B1(new_n462), .B2(G116), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n569), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n559), .B1(new_n568), .B2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT21), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  OAI21_X1  g0376(.A(KEYINPUT83), .B1(new_n563), .B2(new_n567), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n571), .A2(new_n569), .A3(new_n572), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n534), .A2(new_n558), .A3(G179), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n579), .A2(KEYINPUT21), .A3(new_n559), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n552), .A2(new_n576), .A3(new_n582), .A4(new_n583), .ZN(new_n584));
  AND2_X1   g0384(.A1(new_n550), .A2(new_n292), .ZN(new_n585));
  NOR3_X1   g0385(.A1(new_n535), .A2(new_n540), .A3(G190), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n521), .B(new_n525), .C1(new_n585), .C2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n515), .A2(KEYINPUT6), .A3(G97), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n470), .A2(new_n515), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n589), .A2(new_n205), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n588), .B1(new_n590), .B2(KEYINPUT6), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n591), .A2(G20), .B1(G77), .B2(new_n257), .ZN(new_n592));
  INV_X1    g0392(.A(new_n393), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n592), .B1(new_n593), .B2(new_n515), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n252), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n261), .A2(new_n470), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(new_n462), .B2(new_n470), .ZN(new_n597));
  XNOR2_X1  g0397(.A(new_n597), .B(KEYINPUT78), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n531), .A2(new_n533), .B1(G257), .B2(new_n536), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT4), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n282), .A2(G244), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n601), .B1(new_n289), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n280), .A2(G250), .A3(G1698), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n603), .A2(new_n560), .A3(new_n604), .ZN(new_n605));
  NOR3_X1   g0405(.A1(new_n289), .A2(new_n601), .A3(new_n602), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n306), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  AND2_X1   g0407(.A1(new_n600), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n298), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n600), .A2(new_n607), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n320), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n599), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n608), .A2(G190), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n610), .A2(G200), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n613), .A2(new_n595), .A3(new_n598), .A4(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n534), .A2(new_n558), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(G200), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n534), .A2(new_n558), .A3(G190), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n617), .A2(new_n577), .A3(new_n578), .A4(new_n618), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n587), .A2(new_n612), .A3(new_n615), .A4(new_n619), .ZN(new_n620));
  NOR4_X1   g0420(.A1(new_n461), .A2(new_n506), .A3(new_n584), .A4(new_n620), .ZN(G372));
  INV_X1    g0421(.A(new_n612), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n498), .A2(KEYINPUT26), .A3(new_n505), .A4(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n504), .B1(new_n482), .B2(new_n497), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n622), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT26), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n482), .A2(new_n497), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n583), .A2(new_n582), .ZN(new_n631));
  AOI21_X1  g0431(.A(KEYINPUT21), .B1(new_n579), .B2(new_n559), .ZN(new_n632));
  OAI21_X1  g0432(.A(KEYINPUT85), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT85), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n576), .A2(new_n634), .A3(new_n582), .A4(new_n583), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n552), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n612), .A2(new_n615), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n624), .A2(new_n638), .A3(new_n587), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n630), .B1(new_n637), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n461), .B1(new_n628), .B2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n440), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n343), .A2(new_n359), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n460), .B1(new_n323), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n427), .A2(new_n443), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n643), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n297), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n300), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n642), .A2(new_n651), .ZN(G369));
  NAND4_X1  g0452(.A1(new_n576), .A2(new_n582), .A3(new_n583), .A4(new_n619), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n653), .A2(KEYINPUT86), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n655), .A2(KEYINPUT27), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(KEYINPUT27), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n656), .A2(G213), .A3(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(G343), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n579), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n653), .A2(KEYINPUT86), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n654), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT87), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n636), .A2(new_n579), .A3(new_n660), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n663), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n664), .B1(new_n663), .B2(new_n665), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n552), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n526), .A2(new_n660), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n669), .B1(new_n587), .B2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n660), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n671), .B1(new_n669), .B2(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n668), .A2(G330), .A3(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT88), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n668), .A2(KEYINPUT88), .A3(G330), .A4(new_n673), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n576), .A2(new_n582), .A3(new_n583), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n673), .A2(new_n680), .A3(new_n672), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n669), .A2(new_n672), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  OR2_X1    g0483(.A1(new_n679), .A2(new_n683), .ZN(G399));
  INV_X1    g0484(.A(new_n212), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(G41), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR3_X1   g0487(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(G1), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n217), .B2(new_n687), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT28), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n625), .A2(KEYINPUT26), .ZN(new_n692));
  INV_X1    g0492(.A(new_n584), .ZN(new_n693));
  OAI211_X1 g0493(.A(new_n692), .B(new_n629), .C1(new_n639), .C2(new_n693), .ZN(new_n694));
  NOR3_X1   g0494(.A1(new_n506), .A2(KEYINPUT26), .A3(new_n612), .ZN(new_n695));
  OAI211_X1 g0495(.A(KEYINPUT29), .B(new_n672), .C1(new_n694), .C2(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n660), .B1(new_n641), .B2(new_n628), .ZN(new_n697));
  OAI211_X1 g0497(.A(new_n696), .B(KEYINPUT89), .C1(new_n697), .C2(KEYINPUT29), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n620), .A2(new_n584), .ZN(new_n699));
  AOI22_X1  g0499(.A1(new_n482), .A2(new_n483), .B1(new_n495), .B2(new_n496), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n504), .B1(new_n700), .B2(new_n485), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n699), .A2(new_n701), .A3(new_n672), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n494), .A2(G179), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n550), .A2(new_n703), .A3(new_n616), .A4(new_n610), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n547), .A2(new_n549), .A3(new_n494), .ZN(new_n705));
  NOR3_X1   g0505(.A1(new_n705), .A2(new_n610), .A3(new_n580), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n704), .B1(new_n706), .B2(KEYINPUT30), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n547), .A2(new_n549), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n708), .A2(new_n608), .A3(new_n494), .A4(new_n581), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT30), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  OAI211_X1 g0511(.A(KEYINPUT31), .B(new_n660), .C1(new_n707), .C2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n709), .A2(new_n710), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n706), .A2(KEYINPUT30), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n714), .A2(new_n715), .A3(new_n704), .ZN(new_n716));
  AOI21_X1  g0516(.A(KEYINPUT31), .B1(new_n716), .B2(new_n660), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n713), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n702), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(G330), .ZN(new_n720));
  OR2_X1    g0520(.A1(new_n694), .A2(new_n695), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT89), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n721), .A2(new_n722), .A3(KEYINPUT29), .A4(new_n672), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n698), .A2(new_n720), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(KEYINPUT90), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT90), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n698), .A2(new_n723), .A3(new_n726), .A4(new_n720), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n691), .B1(new_n728), .B2(G1), .ZN(G364));
  INV_X1    g0529(.A(G13), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(G20), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n208), .B1(new_n731), .B2(G45), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n686), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n219), .B1(G20), .B2(new_n320), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n209), .A2(new_n298), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G200), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(new_n318), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(G326), .ZN(new_n742));
  INV_X1    g0542(.A(G294), .ZN(new_n743));
  NOR3_X1   g0543(.A1(new_n318), .A2(G179), .A3(G200), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(new_n209), .ZN(new_n745));
  OAI22_X1  g0545(.A1(new_n741), .A2(new_n742), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  XNOR2_X1  g0546(.A(new_n746), .B(KEYINPUT92), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n738), .A2(G190), .A3(new_n292), .ZN(new_n748));
  INV_X1    g0548(.A(G322), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(G190), .A2(G200), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n738), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(G311), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n289), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n209), .A2(G179), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(new_n751), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AOI211_X1 g0557(.A(new_n750), .B(new_n754), .C1(G329), .C2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n739), .A2(G190), .ZN(new_n759));
  INV_X1    g0559(.A(G317), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(KEYINPUT33), .ZN(new_n761));
  OR2_X1    g0561(.A1(new_n760), .A2(KEYINPUT33), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n759), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n755), .A2(G190), .A3(G200), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n755), .A2(new_n318), .A3(G200), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI22_X1  g0567(.A1(new_n765), .A2(G303), .B1(new_n767), .B2(G283), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n747), .A2(new_n758), .A3(new_n763), .A4(new_n768), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n741), .A2(new_n244), .B1(new_n766), .B2(new_n515), .ZN(new_n770));
  INV_X1    g0570(.A(new_n759), .ZN(new_n771));
  OAI22_X1  g0571(.A1(new_n771), .A2(new_n223), .B1(new_n764), .B2(new_n499), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n745), .B(KEYINPUT91), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G97), .ZN(new_n775));
  INV_X1    g0575(.A(G159), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n756), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n777), .B(KEYINPUT32), .ZN(new_n778));
  INV_X1    g0578(.A(G58), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n280), .B1(new_n748), .B2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n752), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n780), .B1(G77), .B2(new_n781), .ZN(new_n782));
  NAND4_X1  g0582(.A1(new_n773), .A2(new_n775), .A3(new_n778), .A4(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n737), .B1(new_n769), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G13), .A2(G33), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(G20), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(new_n736), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n212), .A2(G355), .A3(new_n280), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n401), .A2(new_n402), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n685), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n792), .B1(G45), .B2(new_n217), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n249), .A2(new_n271), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n789), .B1(G116), .B2(new_n212), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n735), .B(new_n784), .C1(new_n788), .C2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n663), .A2(new_n665), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n787), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n796), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n668), .A2(G330), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(new_n735), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n668), .A2(G330), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n800), .B1(new_n802), .B2(new_n803), .ZN(G396));
  NOR2_X1   g0604(.A1(new_n323), .A2(new_n660), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n319), .B1(new_n317), .B2(new_n672), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n805), .B1(new_n323), .B2(new_n806), .ZN(new_n807));
  OR2_X1    g0607(.A1(new_n697), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n628), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n669), .B1(new_n633), .B2(new_n635), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n629), .B1(new_n810), .B2(new_n639), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n672), .B(new_n807), .C1(new_n809), .C2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n808), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n734), .B1(new_n813), .B2(new_n720), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n814), .B1(new_n720), .B2(new_n813), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n736), .A2(new_n785), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n735), .B1(new_n203), .B2(new_n816), .ZN(new_n817));
  AND2_X1   g0617(.A1(new_n771), .A2(KEYINPUT93), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n771), .A2(KEYINPUT93), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n821), .A2(G283), .B1(G116), .B2(new_n781), .ZN(new_n822));
  AND2_X1   g0622(.A1(new_n822), .A2(KEYINPUT94), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n822), .A2(KEYINPUT94), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n289), .B1(new_n756), .B2(new_n753), .C1(new_n741), .C2(new_n553), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n499), .A2(new_n766), .B1(new_n764), .B2(new_n515), .ZN(new_n826));
  NOR4_X1   g0626(.A1(new_n823), .A2(new_n824), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n775), .B1(new_n743), .B2(new_n748), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT95), .ZN(new_n829));
  INV_X1    g0629(.A(new_n748), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n830), .A2(G143), .B1(new_n781), .B2(G159), .ZN(new_n831));
  INV_X1    g0631(.A(G137), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n831), .B1(new_n771), .B2(new_n256), .C1(new_n832), .C2(new_n741), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT34), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n745), .A2(new_n779), .B1(new_n766), .B2(new_n223), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(G50), .B2(new_n765), .ZN(new_n837));
  INV_X1    g0637(.A(G132), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n837), .B(new_n791), .C1(new_n838), .C2(new_n756), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n835), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n833), .A2(new_n834), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n827), .A2(new_n829), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n817), .B1(new_n786), .B2(new_n807), .C1(new_n842), .C2(new_n737), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n815), .A2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(G384));
  INV_X1    g0645(.A(KEYINPUT97), .ZN(new_n846));
  INV_X1    g0646(.A(new_n408), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n252), .B1(new_n420), .B2(KEYINPUT16), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n847), .B1(new_n848), .B2(KEYINPUT96), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT96), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n850), .B(new_n252), .C1(new_n420), .C2(KEYINPUT16), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n413), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n846), .B1(new_n852), .B2(new_n658), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n398), .B1(new_n405), .B2(new_n407), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n414), .B1(new_n854), .B2(new_n422), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n408), .B1(new_n855), .B2(new_n850), .ZN(new_n856));
  INV_X1    g0656(.A(new_n851), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n367), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n658), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n858), .A2(KEYINPUT97), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n853), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n444), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT98), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n444), .A2(KEYINPUT98), .A3(new_n861), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n410), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n867), .B1(new_n858), .B2(new_n433), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n868), .A2(new_n853), .A3(new_n860), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(KEYINPUT37), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n410), .B1(new_n425), .B2(new_n438), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n425), .A2(new_n658), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT99), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT37), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n429), .A2(new_n433), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n429), .A2(new_n859), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n877), .A2(new_n878), .A3(new_n875), .A4(new_n410), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(KEYINPUT99), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n876), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n870), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(KEYINPUT38), .B1(new_n866), .B2(new_n882), .ZN(new_n883));
  AND3_X1   g0683(.A1(new_n444), .A2(KEYINPUT98), .A3(new_n861), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT98), .B1(new_n444), .B2(new_n861), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n882), .B(KEYINPUT38), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(KEYINPUT39), .B1(new_n883), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n441), .A2(new_n442), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n872), .B1(new_n643), .B2(new_n889), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n879), .B(new_n874), .ZN(new_n891));
  OAI21_X1  g0691(.A(KEYINPUT37), .B1(new_n871), .B2(new_n872), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT101), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OAI211_X1 g0694(.A(KEYINPUT101), .B(KEYINPUT37), .C1(new_n871), .C2(new_n872), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n890), .B1(new_n891), .B2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT38), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT39), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n886), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n888), .A2(KEYINPUT100), .A3(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n460), .A2(new_n660), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n882), .B1(new_n884), .B2(new_n885), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n898), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n900), .B1(new_n905), .B2(new_n886), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT100), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n902), .A2(new_n903), .A3(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT102), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n459), .B1(new_n360), .B2(new_n362), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n357), .A2(new_n672), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n912), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n644), .B(new_n914), .C1(new_n459), .C2(new_n357), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n805), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n917), .B1(new_n812), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n905), .A2(new_n886), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n919), .A2(new_n920), .B1(new_n643), .B2(new_n658), .ZN(new_n921));
  AND3_X1   g0721(.A1(new_n909), .A2(new_n910), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n910), .B1(new_n909), .B2(new_n921), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n698), .A2(new_n723), .ZN(new_n925));
  INV_X1    g0725(.A(new_n461), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n651), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  XOR2_X1   g0727(.A(new_n924), .B(new_n927), .Z(new_n928));
  INV_X1    g0728(.A(G330), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n886), .A2(new_n899), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n916), .A2(new_n719), .A3(new_n807), .ZN(new_n931));
  OAI21_X1  g0731(.A(KEYINPUT40), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT40), .ZN(new_n933));
  INV_X1    g0733(.A(new_n931), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n920), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n932), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n461), .B1(new_n702), .B2(new_n718), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n929), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n937), .B2(new_n936), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n928), .A2(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT104), .ZN(new_n941));
  OAI22_X1  g0741(.A1(new_n928), .A2(new_n939), .B1(new_n208), .B2(new_n731), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT103), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n942), .A2(new_n943), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n941), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n591), .A2(KEYINPUT35), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n591), .A2(KEYINPUT35), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n947), .A2(G116), .A3(new_n220), .A4(new_n948), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT36), .ZN(new_n950));
  OAI21_X1  g0750(.A(G77), .B1(new_n779), .B2(new_n223), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n245), .B1(new_n217), .B2(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n952), .A2(G1), .A3(new_n730), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n946), .A2(new_n950), .A3(new_n953), .ZN(G367));
  INV_X1    g0754(.A(new_n792), .ZN(new_n955));
  OAI221_X1 g0755(.A(new_n788), .B1(new_n212), .B2(new_n311), .C1(new_n955), .C2(new_n239), .ZN(new_n956));
  OAI21_X1  g0756(.A(KEYINPUT107), .B1(new_n764), .B2(new_n566), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n821), .A2(G294), .B1(KEYINPUT46), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(KEYINPUT46), .B2(new_n957), .ZN(new_n959));
  AOI22_X1  g0759(.A1(new_n830), .A2(G303), .B1(new_n781), .B2(G283), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n760), .B2(new_n756), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n790), .B1(new_n741), .B2(new_n753), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n745), .A2(new_n515), .B1(new_n766), .B2(new_n470), .ZN(new_n963));
  NOR4_X1   g0763(.A1(new_n959), .A2(new_n961), .A3(new_n962), .A4(new_n963), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT108), .Z(new_n965));
  NAND2_X1  g0765(.A1(new_n821), .A2(G159), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n752), .A2(new_n244), .B1(new_n756), .B2(new_n832), .ZN(new_n967));
  AOI211_X1 g0767(.A(new_n289), .B(new_n967), .C1(G150), .C2(new_n830), .ZN(new_n968));
  INV_X1    g0768(.A(G143), .ZN(new_n969));
  OAI22_X1  g0769(.A1(new_n741), .A2(new_n969), .B1(new_n766), .B2(new_n203), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(G58), .B2(new_n765), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n774), .A2(G68), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n966), .A2(new_n968), .A3(new_n971), .A4(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n965), .A2(new_n973), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n974), .B(KEYINPUT47), .Z(new_n975));
  OAI211_X1 g0775(.A(new_n734), .B(new_n956), .C1(new_n975), .C2(new_n737), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n501), .A2(new_n660), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n629), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n978), .B1(new_n624), .B2(new_n977), .ZN(new_n979));
  AND2_X1   g0779(.A1(new_n979), .A2(new_n787), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n976), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n674), .A2(new_n675), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n599), .A2(new_n660), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n638), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n622), .A2(new_n660), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n680), .A2(new_n672), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n987), .B(new_n682), .C1(new_n671), .C2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT45), .ZN(new_n990));
  OR2_X1    g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n989), .A2(new_n990), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n987), .ZN(new_n994));
  AOI21_X1  g0794(.A(KEYINPUT44), .B1(new_n683), .B2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT44), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n996), .B(new_n987), .C1(new_n681), .C2(new_n682), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n993), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  AND3_X1   g0798(.A1(new_n983), .A2(new_n998), .A3(new_n677), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n998), .B1(new_n983), .B2(new_n677), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n673), .B(new_n988), .Z(new_n1002));
  XNOR2_X1  g0802(.A(new_n801), .B(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(new_n725), .B2(new_n727), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1001), .B1(new_n1004), .B2(KEYINPUT106), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1003), .ZN(new_n1006));
  AND3_X1   g0806(.A1(new_n728), .A2(KEYINPUT106), .A3(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n728), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n686), .B(KEYINPUT41), .Z(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n733), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n681), .A2(new_n994), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n1012), .A2(KEYINPUT42), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(KEYINPUT42), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n612), .B1(new_n985), .B2(new_n552), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n1013), .A2(new_n1014), .B1(new_n672), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT43), .ZN(new_n1017));
  AND2_X1   g0817(.A1(new_n979), .A2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n979), .A2(new_n1017), .ZN(new_n1019));
  NOR3_X1   g0819(.A1(new_n1016), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT105), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1016), .A2(KEYINPUT105), .A3(new_n1018), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1020), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n679), .A2(new_n987), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1025), .B(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n982), .B1(new_n1011), .B2(new_n1028), .ZN(G387));
  INV_X1    g0829(.A(new_n728), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n1003), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n728), .A2(new_n1006), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1031), .A2(new_n686), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n765), .A2(G77), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n741), .B2(new_n776), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n254), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1035), .B1(new_n1036), .B2(new_n759), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n774), .A2(new_n463), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n748), .A2(new_n244), .B1(new_n752), .B2(new_n223), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(G150), .B2(new_n757), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n790), .B1(G97), .B2(new_n767), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n1037), .A2(new_n1038), .A3(new_n1040), .A4(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(G283), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n745), .A2(new_n1043), .B1(new_n764), .B2(new_n743), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n830), .A2(G317), .B1(new_n781), .B2(G303), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1045), .B1(new_n749), .B2(new_n741), .C1(new_n820), .C2(new_n753), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT48), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1044), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(new_n1047), .B2(new_n1046), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT49), .ZN(new_n1050));
  AND2_X1   g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n790), .B1(new_n566), .B2(new_n766), .C1(new_n742), .C2(new_n756), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT110), .Z(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1042), .B1(new_n1051), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT111), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n737), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n1056), .B2(new_n1055), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n271), .B1(new_n223), .B2(new_n203), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n688), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT109), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1059), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  AND3_X1   g0862(.A1(new_n1036), .A2(KEYINPUT50), .A3(new_n244), .ZN(new_n1063));
  AOI21_X1  g0863(.A(KEYINPUT50), .B1(new_n1036), .B2(new_n244), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n1062), .B1(new_n1061), .B2(new_n1060), .C1(new_n1063), .C2(new_n1064), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1065), .B(new_n792), .C1(new_n236), .C2(new_n271), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1060), .A2(new_n212), .A3(new_n280), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1066), .B(new_n1067), .C1(G107), .C2(new_n212), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n735), .B1(new_n1068), .B2(new_n788), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1058), .B(new_n1069), .C1(new_n673), .C2(new_n799), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1033), .B(new_n1070), .C1(new_n732), .C2(new_n1003), .ZN(G393));
  NOR2_X1   g0871(.A1(new_n987), .A2(new_n799), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT112), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n788), .B1(new_n470), .B2(new_n212), .C1(new_n955), .C2(new_n243), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n734), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n745), .A2(new_n566), .B1(new_n752), .B2(new_n743), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n821), .B2(G303), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT114), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(G317), .A2(new_n740), .B1(new_n830), .B2(G311), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1079), .B(new_n1080), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n289), .B1(new_n756), .B2(new_n749), .C1(new_n515), .C2(new_n766), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(G283), .B2(new_n765), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1078), .A2(new_n1081), .A3(new_n1083), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(G150), .A2(new_n740), .B1(new_n830), .B2(G159), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT51), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n223), .A2(new_n764), .B1(new_n766), .B2(new_n499), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n752), .A2(new_n254), .B1(new_n756), .B2(new_n969), .ZN(new_n1088));
  NOR3_X1   g0888(.A1(new_n1087), .A2(new_n790), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n774), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n1089), .B1(new_n203), .B2(new_n1090), .C1(new_n820), .C2(new_n244), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1084), .B1(new_n1086), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1075), .B1(new_n1092), .B2(new_n736), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n1001), .A2(new_n733), .B1(new_n1073), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT106), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1032), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1004), .A2(KEYINPUT106), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1096), .A2(new_n1097), .A3(new_n1001), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n686), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1094), .B1(new_n1099), .B2(new_n1100), .ZN(G390));
  OAI21_X1  g0901(.A(new_n927), .B1(new_n461), .B2(new_n720), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n805), .B1(new_n697), .B2(new_n807), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n719), .A2(G330), .A3(new_n807), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1105), .A2(new_n917), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1105), .A2(new_n917), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1104), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n916), .B(KEYINPUT116), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1105), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1107), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n806), .A2(new_n323), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n672), .B(new_n1114), .C1(new_n694), .C2(new_n695), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n918), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT115), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1115), .A2(KEYINPUT115), .A3(new_n918), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1109), .B1(new_n1113), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1103), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(KEYINPUT118), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n903), .ZN(new_n1125));
  OAI211_X1 g0925(.A(KEYINPUT117), .B(new_n1125), .C1(new_n1104), .C2(new_n917), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT117), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1127), .B1(new_n919), .B2(new_n903), .ZN(new_n1128));
  AND3_X1   g0928(.A1(new_n886), .A2(new_n899), .A3(new_n900), .ZN(new_n1129));
  NOR3_X1   g0929(.A1(new_n906), .A2(new_n1129), .A3(new_n907), .ZN(new_n1130));
  AOI211_X1 g0930(.A(KEYINPUT100), .B(new_n900), .C1(new_n905), .C2(new_n886), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n1126), .B(new_n1128), .C1(new_n1130), .C2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1118), .A2(new_n1119), .A3(new_n1110), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n886), .A2(new_n899), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1133), .A2(new_n1134), .A3(new_n1125), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1132), .A2(new_n1135), .A3(new_n1107), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1107), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1124), .A2(new_n1139), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1123), .B(KEYINPUT118), .C1(new_n1137), .C2(new_n1138), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1140), .A2(new_n686), .A3(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n816), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n223), .A2(new_n766), .B1(new_n764), .B2(new_n499), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(G97), .A2(new_n781), .B1(new_n757), .B2(G294), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1145), .B(new_n289), .C1(new_n566), .C2(new_n748), .ZN(new_n1146));
  AOI211_X1 g0946(.A(new_n1144), .B(new_n1146), .C1(G283), .C2(new_n740), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n821), .A2(G107), .B1(G77), .B2(new_n774), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n821), .A2(G137), .B1(G159), .B2(new_n774), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(KEYINPUT54), .B(G143), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n289), .B1(new_n781), .B2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n764), .A2(new_n256), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT53), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n830), .A2(G132), .B1(new_n757), .B2(G125), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n740), .A2(G128), .B1(new_n767), .B2(G50), .ZN(new_n1156));
  AND4_X1   g0956(.A1(new_n1152), .A2(new_n1154), .A3(new_n1155), .A4(new_n1156), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n1147), .A2(new_n1148), .B1(new_n1149), .B2(new_n1157), .ZN(new_n1158));
  OAI221_X1 g0958(.A(new_n734), .B1(new_n1036), .B2(new_n1143), .C1(new_n1158), .C2(new_n737), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n902), .A2(new_n908), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1159), .B1(new_n1160), .B2(new_n785), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(new_n1139), .B2(new_n733), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1142), .A2(new_n1162), .ZN(G378));
  OAI21_X1  g0963(.A(new_n300), .B1(new_n295), .B2(new_n296), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1164), .A2(new_n267), .A3(new_n859), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n267), .A2(new_n859), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n300), .B(new_n1166), .C1(new_n295), .C2(new_n296), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1165), .A2(new_n1167), .A3(new_n1169), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT120), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1171), .A2(KEYINPUT120), .A3(new_n1172), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n933), .B1(new_n934), .B2(new_n1134), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n916), .A2(new_n719), .A3(new_n933), .A4(new_n807), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(new_n905), .B2(new_n886), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1177), .B(G330), .C1(new_n1178), .C2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1173), .B1(new_n936), .B2(G330), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n922), .A2(new_n923), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n909), .A2(new_n921), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(KEYINPUT102), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1183), .A2(new_n1182), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n909), .A2(new_n910), .A3(new_n921), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  AND2_X1   g0989(.A1(new_n1184), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1132), .A2(new_n1135), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1191), .A2(new_n1106), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1192), .A2(new_n1136), .A3(new_n1122), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(new_n1103), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1190), .A2(new_n1194), .A3(KEYINPUT57), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(new_n686), .ZN(new_n1196));
  AOI21_X1  g0996(.A(KEYINPUT57), .B1(new_n1190), .B2(new_n1194), .ZN(new_n1197));
  OR2_X1    g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1175), .A2(new_n785), .A3(new_n1176), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n734), .B1(G50), .B2(new_n1143), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n766), .A2(new_n779), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1201), .B(KEYINPUT119), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n972), .A2(new_n1202), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n1034), .B1(new_n771), .B2(new_n470), .C1(new_n566), .C2(new_n741), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n790), .A2(new_n270), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n830), .A2(G107), .B1(new_n757), .B2(G283), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1206), .B1(new_n311), .B2(new_n752), .ZN(new_n1207));
  NOR4_X1   g1007(.A1(new_n1203), .A2(new_n1204), .A3(new_n1205), .A4(new_n1207), .ZN(new_n1208));
  OR2_X1    g1008(.A1(new_n1208), .A2(KEYINPUT58), .ZN(new_n1209));
  INV_X1    g1009(.A(G128), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n748), .A2(new_n1210), .B1(new_n752), .B2(new_n832), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(G132), .B2(new_n759), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n740), .A2(G125), .B1(new_n765), .B2(new_n1151), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1212), .B(new_n1213), .C1(new_n1090), .C2(new_n256), .ZN(new_n1214));
  OR2_X1    g1014(.A1(new_n1214), .A2(KEYINPUT59), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(KEYINPUT59), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n767), .A2(G159), .ZN(new_n1217));
  AOI211_X1 g1017(.A(G33), .B(G41), .C1(new_n757), .C2(G124), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .A4(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1208), .A2(KEYINPUT58), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1205), .B(new_n244), .C1(G33), .C2(G41), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1209), .A2(new_n1219), .A3(new_n1220), .A4(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1200), .B1(new_n1222), .B2(new_n736), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1199), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1184), .A2(new_n1189), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1224), .B1(new_n1225), .B2(new_n732), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  AND2_X1   g1027(.A1(new_n1198), .A2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(G375));
  OAI21_X1  g1029(.A(new_n734), .B1(G68), .B2(new_n1143), .ZN(new_n1230));
  OAI221_X1 g1030(.A(new_n791), .B1(new_n776), .B2(new_n764), .C1(new_n838), .C2(new_n741), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n830), .A2(G137), .B1(new_n781), .B2(G150), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1232), .B(new_n1233), .C1(new_n1210), .C2(new_n756), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n1202), .B1(new_n244), .B2(new_n1090), .C1(new_n820), .C2(new_n1150), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n203), .A2(new_n766), .B1(new_n764), .B2(new_n470), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(G294), .B2(new_n740), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n280), .B1(new_n757), .B2(G303), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n830), .A2(G283), .B1(new_n781), .B2(G107), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1237), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1038), .B1(new_n820), .B2(new_n566), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n1234), .A2(new_n1235), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT121), .ZN(new_n1243));
  OR2_X1    g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n737), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1230), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1246), .B1(new_n1110), .B2(new_n786), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1247), .B1(new_n1121), .B2(new_n732), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT122), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(new_n1248), .B(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1102), .A2(new_n1121), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1123), .A2(new_n1010), .A3(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1250), .A2(new_n1252), .ZN(G381));
  NOR2_X1   g1053(.A1(G381), .A2(G384), .ZN(new_n1254));
  INV_X1    g1054(.A(G390), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(G393), .A2(G396), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1254), .A2(new_n1255), .A3(new_n1256), .ZN(new_n1257));
  NOR3_X1   g1057(.A1(new_n1257), .A2(G387), .A3(G378), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1228), .A2(new_n1258), .ZN(G407));
  INV_X1    g1059(.A(G213), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1260), .A2(G343), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(G378), .A2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1228), .A2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(KEYINPUT123), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT123), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1228), .A2(new_n1266), .A3(new_n1263), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1265), .A2(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1260), .B1(new_n1228), .B2(new_n1258), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(KEYINPUT124), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT124), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1268), .A2(new_n1269), .A3(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1271), .A2(new_n1273), .ZN(G409));
  INV_X1    g1074(.A(KEYINPUT125), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n998), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1276), .B1(new_n676), .B2(new_n678), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n983), .A2(new_n998), .A3(new_n677), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1279), .B1(new_n1032), .B2(new_n1095), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1030), .B1(new_n1280), .B2(new_n1097), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n732), .B1(new_n1281), .B2(new_n1009), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n981), .B1(new_n1282), .B2(new_n1027), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1275), .B1(new_n1283), .B2(G390), .ZN(new_n1284));
  XNOR2_X1  g1084(.A(G393), .B(G396), .ZN(new_n1285));
  OAI211_X1 g1085(.A(G390), .B(new_n982), .C1(new_n1011), .C2(new_n1028), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(G387), .A2(new_n1255), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(new_n1284), .A2(new_n1285), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1287), .A2(KEYINPUT125), .A3(new_n1286), .A4(new_n1285), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1288), .A2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT63), .ZN(new_n1292));
  OAI211_X1 g1092(.A(G378), .B(new_n1227), .C1(new_n1196), .C2(new_n1197), .ZN(new_n1293));
  AND3_X1   g1093(.A1(new_n1190), .A2(new_n1194), .A3(new_n1010), .ZN(new_n1294));
  OAI211_X1 g1094(.A(new_n1142), .B(new_n1162), .C1(new_n1294), .C2(new_n1226), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1293), .A2(new_n1295), .ZN(new_n1296));
  OAI21_X1  g1096(.A(KEYINPUT60), .B1(new_n1102), .B2(new_n1121), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n1251), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1102), .A2(new_n1121), .A3(KEYINPUT60), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1298), .A2(new_n686), .A3(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1250), .A2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n844), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1250), .A2(new_n1300), .A3(G384), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1296), .A2(new_n1262), .A3(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1291), .B1(new_n1292), .B2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1296), .A2(new_n1262), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1261), .A2(G2897), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1304), .A2(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1302), .A2(new_n1303), .A3(new_n1309), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1313), .ZN(new_n1314));
  AOI21_X1  g1114(.A(KEYINPUT61), .B1(new_n1308), .B2(new_n1314), .ZN(new_n1315));
  OAI211_X1 g1115(.A(new_n1307), .B(new_n1315), .C1(new_n1292), .C2(new_n1306), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT61), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1261), .B1(new_n1293), .B2(new_n1295), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1317), .B1(new_n1318), .B2(new_n1313), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT62), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1306), .A2(new_n1320), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1318), .A2(KEYINPUT62), .A3(new_n1305), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1319), .B1(new_n1321), .B2(new_n1322), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1291), .B1(new_n1323), .B2(KEYINPUT126), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1322), .ZN(new_n1325));
  AOI21_X1  g1125(.A(KEYINPUT62), .B1(new_n1318), .B2(new_n1305), .ZN(new_n1326));
  OAI211_X1 g1126(.A(KEYINPUT126), .B(new_n1315), .C1(new_n1325), .C2(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1327), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1316), .B1(new_n1324), .B2(new_n1328), .ZN(G405));
  AOI21_X1  g1129(.A(KEYINPUT125), .B1(G387), .B2(new_n1255), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1285), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1286), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1009), .B1(new_n1098), .B2(new_n728), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1027), .B1(new_n1333), .B2(new_n733), .ZN(new_n1334));
  AOI21_X1  g1134(.A(G390), .B1(new_n1334), .B2(new_n982), .ZN(new_n1335));
  OAI22_X1  g1135(.A1(new_n1330), .A2(new_n1331), .B1(new_n1332), .B2(new_n1335), .ZN(new_n1336));
  AND3_X1   g1136(.A1(new_n1336), .A2(new_n1305), .A3(new_n1289), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1305), .B1(new_n1336), .B2(new_n1289), .ZN(new_n1338));
  OAI21_X1  g1138(.A(KEYINPUT127), .B1(new_n1337), .B2(new_n1338), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1304), .B1(new_n1288), .B2(new_n1290), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT127), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1336), .A2(new_n1305), .A3(new_n1289), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1340), .A2(new_n1341), .A3(new_n1342), .ZN(new_n1343));
  NOR2_X1   g1143(.A1(new_n1228), .A2(G378), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1293), .ZN(new_n1345));
  NOR2_X1   g1145(.A1(new_n1344), .A2(new_n1345), .ZN(new_n1346));
  AND3_X1   g1146(.A1(new_n1339), .A2(new_n1343), .A3(new_n1346), .ZN(new_n1347));
  AOI21_X1  g1147(.A(new_n1346), .B1(new_n1339), .B2(new_n1343), .ZN(new_n1348));
  NOR2_X1   g1148(.A1(new_n1347), .A2(new_n1348), .ZN(G402));
endmodule


