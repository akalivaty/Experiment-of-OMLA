

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735;

  NOR2_X1 U367 ( .A1(n521), .A2(n645), .ZN(n532) );
  XNOR2_X2 U368 ( .A(n561), .B(n382), .ZN(n543) );
  XNOR2_X2 U369 ( .A(n414), .B(n413), .ZN(n478) );
  XNOR2_X2 U370 ( .A(KEYINPUT3), .B(G119), .ZN(n414) );
  NOR2_X1 U371 ( .A1(n588), .A2(n676), .ZN(n573) );
  NOR2_X1 U372 ( .A1(n504), .A2(n503), .ZN(n391) );
  XNOR2_X1 U373 ( .A(n480), .B(n479), .ZN(n711) );
  XNOR2_X1 U374 ( .A(n484), .B(G134), .ZN(n451) );
  XNOR2_X2 U375 ( .A(n353), .B(KEYINPUT45), .ZN(n703) );
  INV_X1 U376 ( .A(n601), .ZN(n360) );
  INV_X1 U377 ( .A(G237), .ZN(n422) );
  XNOR2_X1 U378 ( .A(n355), .B(n354), .ZN(n448) );
  INV_X1 U379 ( .A(KEYINPUT8), .ZN(n354) );
  NAND2_X1 U380 ( .A1(n723), .A2(G234), .ZN(n355) );
  XOR2_X1 U381 ( .A(KEYINPUT71), .B(G131), .Z(n465) );
  OR2_X1 U382 ( .A1(n393), .A2(KEYINPUT2), .ZN(n372) );
  NOR2_X1 U383 ( .A1(G953), .A2(G237), .ZN(n460) );
  XNOR2_X1 U384 ( .A(n352), .B(n373), .ZN(n601) );
  INV_X1 U385 ( .A(KEYINPUT48), .ZN(n373) );
  XNOR2_X1 U386 ( .A(n580), .B(n569), .ZN(n661) );
  XNOR2_X1 U387 ( .A(n496), .B(n495), .ZN(n504) );
  XNOR2_X1 U388 ( .A(G119), .B(G128), .ZN(n395) );
  XNOR2_X1 U389 ( .A(KEYINPUT88), .B(KEYINPUT4), .ZN(n482) );
  AND2_X2 U390 ( .A1(n380), .A2(n379), .ZN(n693) );
  NAND2_X1 U391 ( .A1(n603), .A2(KEYINPUT2), .ZN(n379) );
  XNOR2_X1 U392 ( .A(n386), .B(KEYINPUT67), .ZN(n380) );
  XNOR2_X1 U393 ( .A(n381), .B(n522), .ZN(n677) );
  XNOR2_X1 U394 ( .A(n362), .B(n361), .ZN(n599) );
  INV_X1 U395 ( .A(KEYINPUT39), .ZN(n361) );
  NAND2_X1 U396 ( .A1(n365), .A2(n575), .ZN(n362) );
  AND2_X1 U397 ( .A1(n661), .A2(n574), .ZN(n365) );
  NAND2_X1 U398 ( .A1(n375), .A2(n374), .ZN(n581) );
  AND2_X1 U399 ( .A1(n543), .A2(n376), .ZN(n375) );
  NOR2_X1 U400 ( .A1(n563), .A2(n500), .ZN(n376) );
  BUF_X1 U401 ( .A(n504), .Z(n580) );
  INV_X1 U402 ( .A(KEYINPUT0), .ZN(n368) );
  XNOR2_X1 U403 ( .A(n449), .B(n377), .ZN(n700) );
  XNOR2_X1 U404 ( .A(n451), .B(n378), .ZN(n377) );
  XNOR2_X1 U405 ( .A(n479), .B(n450), .ZN(n378) );
  BUF_X1 U406 ( .A(n693), .Z(n699) );
  XNOR2_X1 U407 ( .A(n577), .B(KEYINPUT85), .ZN(n578) );
  NOR2_X1 U408 ( .A1(n731), .A2(n732), .ZN(n579) );
  XOR2_X1 U409 ( .A(KEYINPUT100), .B(KEYINPUT104), .Z(n462) );
  XOR2_X1 U410 ( .A(KEYINPUT11), .B(KEYINPUT103), .Z(n459) );
  XOR2_X1 U411 ( .A(G122), .B(G104), .Z(n469) );
  XNOR2_X1 U412 ( .A(G113), .B(G143), .ZN(n468) );
  XNOR2_X1 U413 ( .A(n451), .B(n347), .ZN(n719) );
  XOR2_X1 U414 ( .A(G146), .B(G125), .Z(n486) );
  INV_X1 U415 ( .A(G113), .ZN(n413) );
  AND2_X1 U416 ( .A1(n359), .A2(n350), .ZN(n383) );
  NAND2_X1 U417 ( .A1(G234), .A2(G237), .ZN(n432) );
  XNOR2_X1 U418 ( .A(n391), .B(n390), .ZN(n589) );
  INV_X1 U419 ( .A(KEYINPUT19), .ZN(n390) );
  XOR2_X1 U420 ( .A(G116), .B(KEYINPUT98), .Z(n411) );
  AND2_X1 U421 ( .A1(n601), .A2(n393), .ZN(n718) );
  XNOR2_X1 U422 ( .A(G122), .B(G116), .ZN(n452) );
  XNOR2_X1 U423 ( .A(n719), .B(G146), .ZN(n430) );
  XNOR2_X1 U424 ( .A(n478), .B(KEYINPUT16), .ZN(n480) );
  AND2_X1 U425 ( .A1(n567), .A2(n566), .ZN(n568) );
  NOR2_X1 U426 ( .A1(n665), .A2(n664), .ZN(n571) );
  NAND2_X1 U427 ( .A1(n700), .A2(n453), .ZN(n455) );
  AND2_X1 U428 ( .A1(n363), .A2(n648), .ZN(n575) );
  XNOR2_X1 U429 ( .A(n423), .B(n364), .ZN(n363) );
  INV_X1 U430 ( .A(KEYINPUT30), .ZN(n364) );
  INV_X1 U431 ( .A(KEYINPUT64), .ZN(n394) );
  XNOR2_X1 U432 ( .A(n400), .B(n356), .ZN(n611) );
  XNOR2_X1 U433 ( .A(n399), .B(n472), .ZN(n356) );
  NAND2_X1 U434 ( .A1(n693), .A2(G475), .ZN(n619) );
  OR2_X1 U435 ( .A1(n723), .A2(G952), .ZN(n620) );
  NOR2_X1 U436 ( .A1(n581), .A2(n580), .ZN(n582) );
  NAND2_X1 U437 ( .A1(n527), .A2(n526), .ZN(n528) );
  NOR2_X1 U438 ( .A1(n646), .A2(n545), .ZN(n546) );
  INV_X1 U439 ( .A(KEYINPUT31), .ZN(n533) );
  INV_X1 U440 ( .A(G110), .ZN(n520) );
  XNOR2_X1 U441 ( .A(n537), .B(KEYINPUT99), .ZN(n371) );
  XNOR2_X1 U442 ( .A(n369), .B(KEYINPUT108), .ZN(n735) );
  NAND2_X1 U443 ( .A1(n517), .A2(n370), .ZN(n369) );
  AND2_X1 U444 ( .A1(n539), .A2(n646), .ZN(n370) );
  XNOR2_X1 U445 ( .A(n358), .B(n357), .ZN(n701) );
  INV_X1 U446 ( .A(n700), .ZN(n357) );
  NAND2_X1 U447 ( .A1(n699), .A2(G478), .ZN(n358) );
  XNOR2_X1 U448 ( .A(n406), .B(n405), .ZN(n560) );
  AND2_X1 U449 ( .A1(n570), .A2(n649), .ZN(n345) );
  AND2_X1 U450 ( .A1(n540), .A2(n735), .ZN(n346) );
  XOR2_X1 U451 ( .A(n465), .B(n408), .Z(n347) );
  AND2_X1 U452 ( .A1(n646), .A2(n536), .ZN(n348) );
  AND2_X1 U453 ( .A1(n536), .A2(n535), .ZN(n349) );
  AND2_X1 U454 ( .A1(n372), .A2(n387), .ZN(n350) );
  INV_X1 U455 ( .A(n624), .ZN(n374) );
  XNOR2_X1 U456 ( .A(n430), .B(n418), .ZN(n604) );
  XOR2_X1 U457 ( .A(n520), .B(KEYINPUT114), .Z(n351) );
  NAND2_X1 U458 ( .A1(n597), .A2(n596), .ZN(n352) );
  NAND2_X1 U459 ( .A1(n360), .A2(n681), .ZN(n359) );
  NAND2_X1 U460 ( .A1(n559), .A2(n558), .ZN(n353) );
  NOR2_X1 U461 ( .A1(n677), .A2(n366), .ZN(n524) );
  NOR2_X2 U462 ( .A1(n614), .A2(n702), .ZN(n615) );
  NOR2_X2 U463 ( .A1(n691), .A2(n702), .ZN(n692) );
  INV_X1 U464 ( .A(n555), .ZN(n553) );
  NAND2_X1 U465 ( .A1(n550), .A2(n551), .ZN(n555) );
  INV_X1 U466 ( .A(n514), .ZN(n366) );
  AND2_X1 U467 ( .A1(n514), .A2(n367), .ZN(n534) );
  INV_X1 U468 ( .A(n655), .ZN(n367) );
  NAND2_X1 U469 ( .A1(n514), .A2(n349), .ZN(n537) );
  XNOR2_X2 U470 ( .A(n512), .B(n368), .ZN(n514) );
  NOR2_X1 U471 ( .A1(n371), .A2(n639), .ZN(n538) );
  NAND2_X1 U472 ( .A1(n371), .A2(n638), .ZN(n626) );
  NAND2_X1 U473 ( .A1(n371), .A2(n374), .ZN(n625) );
  INV_X1 U474 ( .A(n703), .ZN(n385) );
  AND2_X1 U475 ( .A1(n703), .A2(n718), .ZN(n603) );
  AND2_X2 U476 ( .A1(n517), .A2(n348), .ZN(n518) );
  XNOR2_X1 U477 ( .A(n551), .B(n351), .ZN(G12) );
  NAND2_X1 U478 ( .A1(n519), .A2(n560), .ZN(n551) );
  NAND2_X1 U479 ( .A1(n385), .A2(n681), .ZN(n384) );
  NAND2_X1 U480 ( .A1(n384), .A2(n383), .ZN(n386) );
  NAND2_X1 U481 ( .A1(n532), .A2(n543), .ZN(n381) );
  INV_X1 U482 ( .A(KEYINPUT6), .ZN(n382) );
  XNOR2_X2 U483 ( .A(n421), .B(n420), .ZN(n561) );
  XNOR2_X2 U484 ( .A(n409), .B(G128), .ZN(n484) );
  INV_X1 U485 ( .A(n602), .ZN(n387) );
  XNOR2_X1 U486 ( .A(n388), .B(n541), .ZN(n559) );
  NAND2_X1 U487 ( .A1(n346), .A2(n389), .ZN(n388) );
  NAND2_X1 U488 ( .A1(n730), .A2(KEYINPUT44), .ZN(n389) );
  XNOR2_X2 U489 ( .A(n528), .B(KEYINPUT35), .ZN(n730) );
  NAND2_X1 U490 ( .A1(n589), .A2(n511), .ZN(n512) );
  XOR2_X1 U491 ( .A(n425), .B(n424), .Z(n392) );
  NOR2_X1 U492 ( .A1(n643), .A2(n600), .ZN(n393) );
  INV_X1 U493 ( .A(G137), .ZN(n407) );
  XNOR2_X1 U494 ( .A(n407), .B(KEYINPUT4), .ZN(n408) );
  INV_X1 U495 ( .A(KEYINPUT82), .ZN(n542) );
  INV_X1 U496 ( .A(KEYINPUT33), .ZN(n522) );
  XNOR2_X1 U497 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U498 ( .A(n392), .B(n481), .ZN(n429) );
  XNOR2_X1 U499 ( .A(n430), .B(n429), .ZN(n694) );
  XNOR2_X1 U500 ( .A(n694), .B(n695), .ZN(n696) );
  XNOR2_X1 U501 ( .A(n534), .B(n533), .ZN(n639) );
  XNOR2_X1 U502 ( .A(n697), .B(n696), .ZN(n698) );
  XNOR2_X2 U503 ( .A(n394), .B(G953), .ZN(n723) );
  NAND2_X1 U504 ( .A1(G221), .A2(n448), .ZN(n400) );
  XOR2_X1 U505 ( .A(G110), .B(G137), .Z(n396) );
  XNOR2_X1 U506 ( .A(n396), .B(n395), .ZN(n398) );
  XOR2_X1 U507 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n397) );
  XOR2_X1 U508 ( .A(G140), .B(KEYINPUT10), .Z(n401) );
  XNOR2_X1 U509 ( .A(n486), .B(n401), .ZN(n721) );
  INV_X1 U510 ( .A(n721), .ZN(n472) );
  INV_X1 U511 ( .A(G902), .ZN(n453) );
  NAND2_X1 U512 ( .A1(n611), .A2(n453), .ZN(n406) );
  XNOR2_X1 U513 ( .A(G902), .B(KEYINPUT15), .ZN(n602) );
  NAND2_X1 U514 ( .A1(G234), .A2(n602), .ZN(n402) );
  XNOR2_X1 U515 ( .A(KEYINPUT20), .B(n402), .ZN(n442) );
  NAND2_X1 U516 ( .A1(n442), .A2(G217), .ZN(n404) );
  XNOR2_X1 U517 ( .A(KEYINPUT25), .B(KEYINPUT78), .ZN(n403) );
  XNOR2_X1 U518 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X2 U519 ( .A(G143), .B(KEYINPUT66), .ZN(n409) );
  NAND2_X1 U520 ( .A1(n460), .A2(G210), .ZN(n410) );
  XNOR2_X1 U521 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U522 ( .A(n412), .B(KEYINPUT5), .Z(n417) );
  XOR2_X1 U523 ( .A(G101), .B(KEYINPUT70), .Z(n426) );
  INV_X1 U524 ( .A(n478), .ZN(n415) );
  XNOR2_X1 U525 ( .A(n426), .B(n415), .ZN(n416) );
  XNOR2_X1 U526 ( .A(n417), .B(n416), .ZN(n418) );
  NAND2_X1 U527 ( .A1(n604), .A2(n453), .ZN(n421) );
  INV_X1 U528 ( .A(KEYINPUT75), .ZN(n419) );
  XNOR2_X1 U529 ( .A(n419), .B(G472), .ZN(n420) );
  NAND2_X1 U530 ( .A1(n453), .A2(n422), .ZN(n493) );
  NAND2_X1 U531 ( .A1(n493), .A2(G214), .ZN(n660) );
  NAND2_X1 U532 ( .A1(n561), .A2(n660), .ZN(n423) );
  XOR2_X1 U533 ( .A(G107), .B(G140), .Z(n425) );
  NAND2_X1 U534 ( .A1(G227), .A2(n723), .ZN(n424) );
  XNOR2_X1 U535 ( .A(n426), .B(KEYINPUT73), .ZN(n428) );
  XOR2_X1 U536 ( .A(G104), .B(KEYINPUT77), .Z(n427) );
  XNOR2_X1 U537 ( .A(n427), .B(n520), .ZN(n710) );
  XNOR2_X1 U538 ( .A(n428), .B(n710), .ZN(n481) );
  NOR2_X1 U539 ( .A1(n694), .A2(G902), .ZN(n431) );
  XNOR2_X2 U540 ( .A(n431), .B(G469), .ZN(n565) );
  XOR2_X1 U541 ( .A(KEYINPUT14), .B(KEYINPUT91), .Z(n433) );
  XNOR2_X1 U542 ( .A(n433), .B(n432), .ZN(n437) );
  NAND2_X1 U543 ( .A1(n437), .A2(G952), .ZN(n434) );
  XNOR2_X1 U544 ( .A(n434), .B(KEYINPUT92), .ZN(n675) );
  NOR2_X1 U545 ( .A1(G953), .A2(n675), .ZN(n436) );
  INV_X1 U546 ( .A(KEYINPUT93), .ZN(n435) );
  XNOR2_X1 U547 ( .A(n436), .B(n435), .ZN(n505) );
  NAND2_X1 U548 ( .A1(n437), .A2(G902), .ZN(n438) );
  XOR2_X1 U549 ( .A(n438), .B(KEYINPUT95), .Z(n506) );
  OR2_X1 U550 ( .A1(n723), .A2(n506), .ZN(n439) );
  NOR2_X1 U551 ( .A1(G900), .A2(n439), .ZN(n440) );
  NOR2_X1 U552 ( .A1(n505), .A2(n440), .ZN(n441) );
  XNOR2_X1 U553 ( .A(KEYINPUT83), .B(n441), .ZN(n447) );
  XOR2_X1 U554 ( .A(KEYINPUT97), .B(KEYINPUT21), .Z(n444) );
  NAND2_X1 U555 ( .A1(G221), .A2(n442), .ZN(n443) );
  XNOR2_X1 U556 ( .A(n444), .B(n443), .ZN(n446) );
  INV_X1 U557 ( .A(KEYINPUT96), .ZN(n445) );
  XNOR2_X1 U558 ( .A(n446), .B(n445), .ZN(n649) );
  NAND2_X1 U559 ( .A1(n447), .A2(n649), .ZN(n499) );
  NOR2_X1 U560 ( .A1(n565), .A2(n499), .ZN(n574) );
  NAND2_X1 U561 ( .A1(n575), .A2(n574), .ZN(n477) );
  XOR2_X1 U562 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n450) );
  NAND2_X1 U563 ( .A1(G217), .A2(n448), .ZN(n449) );
  XNOR2_X1 U564 ( .A(n452), .B(G107), .ZN(n479) );
  INV_X1 U565 ( .A(G478), .ZN(n454) );
  XNOR2_X1 U566 ( .A(n455), .B(n454), .ZN(n530) );
  INV_X1 U567 ( .A(n530), .ZN(n476) );
  XOR2_X1 U568 ( .A(KEYINPUT106), .B(KEYINPUT13), .Z(n457) );
  XNOR2_X1 U569 ( .A(KEYINPUT105), .B(G475), .ZN(n456) );
  XNOR2_X1 U570 ( .A(n457), .B(n456), .ZN(n475) );
  XNOR2_X1 U571 ( .A(KEYINPUT101), .B(KEYINPUT102), .ZN(n458) );
  XNOR2_X1 U572 ( .A(n459), .B(n458), .ZN(n464) );
  NAND2_X1 U573 ( .A1(G214), .A2(n460), .ZN(n461) );
  XNOR2_X1 U574 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U575 ( .A(n464), .B(n463), .ZN(n467) );
  XNOR2_X1 U576 ( .A(n465), .B(KEYINPUT12), .ZN(n466) );
  XNOR2_X1 U577 ( .A(n467), .B(n466), .ZN(n471) );
  XOR2_X1 U578 ( .A(n469), .B(n468), .Z(n470) );
  XNOR2_X1 U579 ( .A(n471), .B(n470), .ZN(n473) );
  XNOR2_X1 U580 ( .A(n473), .B(n472), .ZN(n617) );
  NOR2_X1 U581 ( .A1(G902), .A2(n617), .ZN(n474) );
  XNOR2_X1 U582 ( .A(n475), .B(n474), .ZN(n529) );
  NAND2_X1 U583 ( .A1(n476), .A2(n529), .ZN(n525) );
  NOR2_X1 U584 ( .A1(n477), .A2(n525), .ZN(n498) );
  XNOR2_X1 U585 ( .A(n711), .B(n481), .ZN(n492) );
  NAND2_X1 U586 ( .A1(n723), .A2(G224), .ZN(n483) );
  XNOR2_X1 U587 ( .A(n483), .B(n482), .ZN(n485) );
  XNOR2_X1 U588 ( .A(n485), .B(n484), .ZN(n490) );
  XNOR2_X1 U589 ( .A(KEYINPUT18), .B(n486), .ZN(n488) );
  XOR2_X1 U590 ( .A(KEYINPUT79), .B(KEYINPUT17), .Z(n487) );
  XNOR2_X1 U591 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U592 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U593 ( .A(n492), .B(n491), .ZN(n686) );
  NAND2_X1 U594 ( .A1(n686), .A2(n602), .ZN(n496) );
  NAND2_X1 U595 ( .A1(n493), .A2(G210), .ZN(n494) );
  XNOR2_X1 U596 ( .A(n494), .B(KEYINPUT90), .ZN(n495) );
  INV_X1 U597 ( .A(n580), .ZN(n497) );
  NAND2_X1 U598 ( .A1(n498), .A2(n497), .ZN(n585) );
  XNOR2_X1 U599 ( .A(n585), .B(G143), .ZN(G45) );
  XNOR2_X1 U600 ( .A(n565), .B(KEYINPUT1), .ZN(n521) );
  INV_X1 U601 ( .A(n521), .ZN(n516) );
  NAND2_X1 U602 ( .A1(n660), .A2(n560), .ZN(n500) );
  NAND2_X1 U603 ( .A1(n530), .A2(n529), .ZN(n624) );
  XNOR2_X1 U604 ( .A(n499), .B(KEYINPUT72), .ZN(n563) );
  OR2_X1 U605 ( .A1(n516), .A2(n581), .ZN(n501) );
  XNOR2_X1 U606 ( .A(KEYINPUT43), .B(n501), .ZN(n502) );
  AND2_X1 U607 ( .A1(n580), .A2(n502), .ZN(n600) );
  XOR2_X1 U608 ( .A(n600), .B(G140), .Z(G42) );
  INV_X1 U609 ( .A(n660), .ZN(n503) );
  INV_X1 U610 ( .A(n505), .ZN(n510) );
  INV_X1 U611 ( .A(n506), .ZN(n508) );
  XOR2_X1 U612 ( .A(G898), .B(KEYINPUT94), .Z(n707) );
  NAND2_X1 U613 ( .A1(G953), .A2(n707), .ZN(n713) );
  INV_X1 U614 ( .A(n713), .ZN(n507) );
  NAND2_X1 U615 ( .A1(n508), .A2(n507), .ZN(n509) );
  NAND2_X1 U616 ( .A1(n510), .A2(n509), .ZN(n511) );
  INV_X1 U617 ( .A(n529), .ZN(n513) );
  AND2_X1 U618 ( .A1(n513), .A2(n530), .ZN(n570) );
  NAND2_X1 U619 ( .A1(n514), .A2(n345), .ZN(n515) );
  XNOR2_X1 U620 ( .A(n515), .B(KEYINPUT22), .ZN(n547) );
  INV_X1 U621 ( .A(n547), .ZN(n517) );
  INV_X1 U622 ( .A(n516), .ZN(n646) );
  INV_X1 U623 ( .A(n561), .ZN(n536) );
  INV_X1 U624 ( .A(n536), .ZN(n652) );
  XNOR2_X1 U625 ( .A(n518), .B(KEYINPUT68), .ZN(n519) );
  INV_X1 U626 ( .A(n560), .ZN(n648) );
  NAND2_X1 U627 ( .A1(n648), .A2(n649), .ZN(n645) );
  XNOR2_X1 U628 ( .A(KEYINPUT74), .B(KEYINPUT34), .ZN(n523) );
  XNOR2_X1 U629 ( .A(n524), .B(n523), .ZN(n527) );
  XOR2_X1 U630 ( .A(n525), .B(KEYINPUT80), .Z(n526) );
  NOR2_X1 U631 ( .A1(n530), .A2(n529), .ZN(n638) );
  INV_X1 U632 ( .A(n638), .ZN(n598) );
  NAND2_X1 U633 ( .A1(n598), .A2(n624), .ZN(n531) );
  XNOR2_X1 U634 ( .A(n531), .B(KEYINPUT107), .ZN(n666) );
  NAND2_X1 U635 ( .A1(n652), .A2(n532), .ZN(n655) );
  NOR2_X1 U636 ( .A1(n565), .A2(n645), .ZN(n535) );
  OR2_X1 U637 ( .A1(n666), .A2(n538), .ZN(n540) );
  NOR2_X1 U638 ( .A1(n543), .A2(n560), .ZN(n539) );
  INV_X1 U639 ( .A(KEYINPUT86), .ZN(n541) );
  XNOR2_X1 U640 ( .A(n543), .B(n542), .ZN(n544) );
  NAND2_X1 U641 ( .A1(n544), .A2(n560), .ZN(n545) );
  XNOR2_X1 U642 ( .A(n546), .B(KEYINPUT81), .ZN(n548) );
  NOR2_X1 U643 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U644 ( .A(n549), .B(KEYINPUT32), .ZN(n733) );
  INV_X1 U645 ( .A(n733), .ZN(n550) );
  OR2_X1 U646 ( .A1(n730), .A2(KEYINPUT44), .ZN(n552) );
  NAND2_X1 U647 ( .A1(n553), .A2(n552), .ZN(n557) );
  INV_X1 U648 ( .A(KEYINPUT44), .ZN(n554) );
  NAND2_X1 U649 ( .A1(n555), .A2(n554), .ZN(n556) );
  NAND2_X1 U650 ( .A1(n557), .A2(n556), .ZN(n558) );
  NAND2_X1 U651 ( .A1(n561), .A2(n560), .ZN(n562) );
  NOR2_X1 U652 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U653 ( .A(n564), .B(KEYINPUT28), .ZN(n567) );
  INV_X1 U654 ( .A(n565), .ZN(n566) );
  XNOR2_X1 U655 ( .A(n568), .B(KEYINPUT109), .ZN(n588) );
  XNOR2_X1 U656 ( .A(KEYINPUT76), .B(KEYINPUT38), .ZN(n569) );
  NAND2_X1 U657 ( .A1(n661), .A2(n660), .ZN(n665) );
  INV_X1 U658 ( .A(n570), .ZN(n664) );
  XNOR2_X1 U659 ( .A(n571), .B(KEYINPUT41), .ZN(n676) );
  XNOR2_X1 U660 ( .A(KEYINPUT110), .B(KEYINPUT42), .ZN(n572) );
  XNOR2_X1 U661 ( .A(n573), .B(n572), .ZN(n731) );
  NOR2_X1 U662 ( .A1(n624), .A2(n599), .ZN(n576) );
  XNOR2_X1 U663 ( .A(KEYINPUT40), .B(n576), .ZN(n732) );
  XNOR2_X1 U664 ( .A(KEYINPUT46), .B(KEYINPUT65), .ZN(n577) );
  XNOR2_X1 U665 ( .A(n579), .B(n578), .ZN(n597) );
  XOR2_X1 U666 ( .A(KEYINPUT36), .B(n582), .Z(n583) );
  NOR2_X1 U667 ( .A1(n646), .A2(n583), .ZN(n641) );
  NAND2_X1 U668 ( .A1(KEYINPUT47), .A2(n666), .ZN(n584) );
  NAND2_X1 U669 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U670 ( .A(KEYINPUT84), .B(n586), .ZN(n587) );
  NOR2_X1 U671 ( .A1(n641), .A2(n587), .ZN(n595) );
  INV_X1 U672 ( .A(n588), .ZN(n590) );
  NAND2_X1 U673 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U674 ( .A(n591), .B(KEYINPUT47), .ZN(n593) );
  INV_X1 U675 ( .A(n591), .ZN(n634) );
  NAND2_X1 U676 ( .A1(n634), .A2(n666), .ZN(n592) );
  NAND2_X1 U677 ( .A1(n593), .A2(n592), .ZN(n594) );
  AND2_X1 U678 ( .A1(n595), .A2(n594), .ZN(n596) );
  NOR2_X1 U679 ( .A1(n599), .A2(n598), .ZN(n643) );
  INV_X1 U680 ( .A(KEYINPUT2), .ZN(n681) );
  NAND2_X1 U681 ( .A1(n693), .A2(G472), .ZN(n608) );
  XNOR2_X1 U682 ( .A(KEYINPUT111), .B(KEYINPUT112), .ZN(n605) );
  XOR2_X1 U683 ( .A(n605), .B(KEYINPUT62), .Z(n606) );
  XNOR2_X1 U684 ( .A(n604), .B(n606), .ZN(n607) );
  XNOR2_X1 U685 ( .A(n608), .B(n607), .ZN(n609) );
  NAND2_X1 U686 ( .A1(n609), .A2(n620), .ZN(n610) );
  XNOR2_X1 U687 ( .A(n610), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U688 ( .A1(n693), .A2(G217), .ZN(n613) );
  XNOR2_X1 U689 ( .A(n611), .B(KEYINPUT123), .ZN(n612) );
  XNOR2_X1 U690 ( .A(n613), .B(n612), .ZN(n614) );
  INV_X1 U691 ( .A(n620), .ZN(n702) );
  XNOR2_X1 U692 ( .A(n615), .B(KEYINPUT124), .ZN(G66) );
  XOR2_X1 U693 ( .A(KEYINPUT89), .B(KEYINPUT59), .Z(n616) );
  XNOR2_X1 U694 ( .A(n617), .B(n616), .ZN(n618) );
  XNOR2_X1 U695 ( .A(n619), .B(n618), .ZN(n621) );
  NAND2_X1 U696 ( .A1(n621), .A2(n620), .ZN(n623) );
  XNOR2_X1 U697 ( .A(KEYINPUT69), .B(KEYINPUT60), .ZN(n622) );
  XNOR2_X1 U698 ( .A(n623), .B(n622), .ZN(G60) );
  XNOR2_X1 U699 ( .A(n625), .B(G104), .ZN(G6) );
  XOR2_X1 U700 ( .A(G107), .B(KEYINPUT26), .Z(n627) );
  XNOR2_X1 U701 ( .A(n627), .B(n626), .ZN(n629) );
  XOR2_X1 U702 ( .A(KEYINPUT27), .B(KEYINPUT113), .Z(n628) );
  XNOR2_X1 U703 ( .A(n629), .B(n628), .ZN(G9) );
  XOR2_X1 U704 ( .A(KEYINPUT29), .B(KEYINPUT116), .Z(n631) );
  NAND2_X1 U705 ( .A1(n634), .A2(n638), .ZN(n630) );
  XNOR2_X1 U706 ( .A(n631), .B(n630), .ZN(n633) );
  XOR2_X1 U707 ( .A(G128), .B(KEYINPUT115), .Z(n632) );
  XNOR2_X1 U708 ( .A(n633), .B(n632), .ZN(G30) );
  NAND2_X1 U709 ( .A1(n634), .A2(n374), .ZN(n635) );
  XNOR2_X1 U710 ( .A(n635), .B(G146), .ZN(G48) );
  XOR2_X1 U711 ( .A(G113), .B(KEYINPUT117), .Z(n637) );
  NAND2_X1 U712 ( .A1(n639), .A2(n374), .ZN(n636) );
  XNOR2_X1 U713 ( .A(n637), .B(n636), .ZN(G15) );
  NAND2_X1 U714 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U715 ( .A(n640), .B(G116), .ZN(G18) );
  XNOR2_X1 U716 ( .A(G125), .B(n641), .ZN(n642) );
  XNOR2_X1 U717 ( .A(n642), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U718 ( .A(G134), .B(n643), .Z(G36) );
  XNOR2_X1 U719 ( .A(KEYINPUT51), .B(KEYINPUT118), .ZN(n644) );
  XNOR2_X1 U720 ( .A(n644), .B(KEYINPUT119), .ZN(n658) );
  NAND2_X1 U721 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U722 ( .A(n647), .B(KEYINPUT50), .ZN(n654) );
  NOR2_X1 U723 ( .A1(n649), .A2(n648), .ZN(n650) );
  XOR2_X1 U724 ( .A(KEYINPUT49), .B(n650), .Z(n651) );
  NOR2_X1 U725 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U726 ( .A1(n654), .A2(n653), .ZN(n656) );
  NAND2_X1 U727 ( .A1(n656), .A2(n655), .ZN(n657) );
  XOR2_X1 U728 ( .A(n658), .B(n657), .Z(n659) );
  NOR2_X1 U729 ( .A1(n676), .A2(n659), .ZN(n672) );
  NOR2_X1 U730 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U731 ( .A(n662), .B(KEYINPUT120), .ZN(n663) );
  NOR2_X1 U732 ( .A1(n664), .A2(n663), .ZN(n668) );
  NOR2_X1 U733 ( .A1(n666), .A2(n665), .ZN(n667) );
  NOR2_X1 U734 ( .A1(n668), .A2(n667), .ZN(n669) );
  NOR2_X1 U735 ( .A1(n677), .A2(n669), .ZN(n670) );
  XOR2_X1 U736 ( .A(KEYINPUT121), .B(n670), .Z(n671) );
  NOR2_X1 U737 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U738 ( .A(n673), .B(KEYINPUT52), .ZN(n674) );
  NOR2_X1 U739 ( .A1(n675), .A2(n674), .ZN(n679) );
  NOR2_X1 U740 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U741 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U742 ( .A(KEYINPUT122), .B(n680), .ZN(n684) );
  XNOR2_X1 U743 ( .A(n603), .B(n681), .ZN(n682) );
  NOR2_X1 U744 ( .A1(n682), .A2(G953), .ZN(n683) );
  NAND2_X1 U745 ( .A1(n684), .A2(n683), .ZN(n685) );
  XOR2_X1 U746 ( .A(KEYINPUT53), .B(n685), .Z(G75) );
  NAND2_X1 U747 ( .A1(n693), .A2(G210), .ZN(n690) );
  XOR2_X1 U748 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n687) );
  XNOR2_X1 U749 ( .A(n687), .B(KEYINPUT87), .ZN(n688) );
  XNOR2_X1 U750 ( .A(n686), .B(n688), .ZN(n689) );
  XNOR2_X1 U751 ( .A(n690), .B(n689), .ZN(n691) );
  XNOR2_X1 U752 ( .A(n692), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U753 ( .A1(n699), .A2(G469), .ZN(n697) );
  XOR2_X1 U754 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n695) );
  NOR2_X1 U755 ( .A1(n702), .A2(n698), .ZN(G54) );
  NOR2_X1 U756 ( .A1(n702), .A2(n701), .ZN(G63) );
  INV_X1 U757 ( .A(n703), .ZN(n704) );
  NOR2_X1 U758 ( .A1(n704), .A2(G953), .ZN(n709) );
  NAND2_X1 U759 ( .A1(G953), .A2(G224), .ZN(n705) );
  XOR2_X1 U760 ( .A(KEYINPUT61), .B(n705), .Z(n706) );
  NOR2_X1 U761 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X1 U762 ( .A1(n709), .A2(n708), .ZN(n716) );
  XOR2_X1 U763 ( .A(n710), .B(G101), .Z(n712) );
  XNOR2_X1 U764 ( .A(n711), .B(n712), .ZN(n714) );
  NAND2_X1 U765 ( .A1(n714), .A2(n713), .ZN(n715) );
  XOR2_X1 U766 ( .A(n716), .B(n715), .Z(n717) );
  XNOR2_X1 U767 ( .A(KEYINPUT125), .B(n717), .ZN(G69) );
  INV_X1 U768 ( .A(n718), .ZN(n722) );
  XOR2_X1 U769 ( .A(n719), .B(KEYINPUT126), .Z(n720) );
  XNOR2_X1 U770 ( .A(n721), .B(n720), .ZN(n725) );
  XNOR2_X1 U771 ( .A(n722), .B(n725), .ZN(n724) );
  NAND2_X1 U772 ( .A1(n724), .A2(n723), .ZN(n729) );
  XNOR2_X1 U773 ( .A(G227), .B(n725), .ZN(n726) );
  NAND2_X1 U774 ( .A1(n726), .A2(G900), .ZN(n727) );
  NAND2_X1 U775 ( .A1(n727), .A2(G953), .ZN(n728) );
  NAND2_X1 U776 ( .A1(n729), .A2(n728), .ZN(G72) );
  XOR2_X1 U777 ( .A(n730), .B(G122), .Z(G24) );
  XOR2_X1 U778 ( .A(n731), .B(G137), .Z(G39) );
  XOR2_X1 U779 ( .A(G131), .B(n732), .Z(G33) );
  XNOR2_X1 U780 ( .A(G119), .B(KEYINPUT127), .ZN(n734) );
  XNOR2_X1 U781 ( .A(n734), .B(n733), .ZN(G21) );
  XNOR2_X1 U782 ( .A(G101), .B(n735), .ZN(G3) );
endmodule

