//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 0 1 0 1 1 0 0 1 0 1 0 0 1 1 1 1 0 1 1 1 1 1 1 1 0 1 0 1 1 1 1 0 1 1 0 1 1 0 1 1 1 1 1 1 1 1 0 1 0 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:31 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012;
  INV_X1    g000(.A(KEYINPUT66), .ZN(new_n187));
  INV_X1    g001(.A(G116), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G119), .ZN(new_n189));
  INV_X1    g003(.A(G119), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(KEYINPUT66), .A3(G116), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n188), .A2(G119), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT2), .B(G113), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n190), .A2(G116), .ZN(new_n196));
  OAI21_X1  g010(.A(G113), .B1(new_n196), .B2(KEYINPUT5), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n193), .A2(KEYINPUT67), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT67), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n189), .A2(new_n191), .A3(new_n199), .A4(new_n192), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n197), .B1(new_n201), .B2(KEYINPUT5), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n195), .B1(new_n202), .B2(KEYINPUT88), .ZN(new_n203));
  INV_X1    g017(.A(G104), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT3), .B1(new_n204), .B2(G107), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT3), .ZN(new_n206));
  INV_X1    g020(.A(G107), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(new_n207), .A3(G104), .ZN(new_n208));
  INV_X1    g022(.A(G101), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n204), .A2(G107), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n205), .A2(new_n208), .A3(new_n209), .A4(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n207), .A2(G104), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(new_n210), .ZN(new_n213));
  AOI21_X1  g027(.A(KEYINPUT81), .B1(new_n213), .B2(G101), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT81), .ZN(new_n215));
  AOI211_X1 g029(.A(new_n215), .B(new_n209), .C1(new_n212), .C2(new_n210), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n211), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT83), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI211_X1 g033(.A(KEYINPUT83), .B(new_n211), .C1(new_n214), .C2(new_n216), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT88), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT5), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n223), .B1(new_n198), .B2(new_n200), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n222), .B1(new_n224), .B2(new_n197), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n203), .A2(new_n221), .A3(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n205), .A2(new_n208), .A3(new_n210), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G101), .ZN(new_n228));
  OAI21_X1  g042(.A(KEYINPUT80), .B1(new_n228), .B2(KEYINPUT4), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT80), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT4), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n227), .A2(new_n230), .A3(new_n231), .A4(G101), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n228), .A2(KEYINPUT79), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT79), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n227), .A2(new_n235), .A3(G101), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n234), .A2(KEYINPUT4), .A3(new_n211), .A4(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT87), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n198), .A2(new_n194), .A3(new_n200), .ZN(new_n239));
  INV_X1    g053(.A(new_n195), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n233), .A2(new_n237), .A3(new_n238), .A4(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n233), .A2(new_n237), .A3(new_n241), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(KEYINPUT87), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n226), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  XNOR2_X1  g059(.A(G110), .B(G122), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n226), .A2(new_n244), .A3(new_n246), .A4(new_n242), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n248), .A2(KEYINPUT6), .A3(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT6), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n245), .A2(new_n251), .A3(new_n247), .ZN(new_n252));
  INV_X1    g066(.A(G128), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n253), .A2(KEYINPUT1), .ZN(new_n254));
  INV_X1    g068(.A(G146), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G143), .ZN(new_n256));
  INV_X1    g070(.A(G143), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G146), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n254), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n257), .A2(G146), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT64), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n261), .B1(new_n255), .B2(G143), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n257), .A2(KEYINPUT64), .A3(G146), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n260), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n253), .B1(new_n256), .B2(KEYINPUT1), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n259), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(G125), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AND2_X1   g083(.A1(KEYINPUT0), .A2(G128), .ZN(new_n270));
  AND3_X1   g084(.A1(new_n256), .A2(new_n258), .A3(new_n270), .ZN(new_n271));
  AND3_X1   g085(.A1(new_n257), .A2(KEYINPUT64), .A3(G146), .ZN(new_n272));
  AOI21_X1  g086(.A(KEYINPUT64), .B1(new_n257), .B2(G146), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n256), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NOR2_X1   g088(.A1(KEYINPUT0), .A2(G128), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n270), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n271), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n269), .B1(new_n268), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(G224), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n279), .A2(G953), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n278), .B(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n250), .A2(new_n252), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT7), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n278), .B(new_n284), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n249), .A2(new_n285), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n246), .B(KEYINPUT8), .ZN(new_n287));
  INV_X1    g101(.A(new_n220), .ZN(new_n288));
  XNOR2_X1  g102(.A(G104), .B(G107), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n215), .B1(new_n289), .B2(new_n209), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n213), .A2(KEYINPUT81), .A3(G101), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(KEYINPUT83), .B1(new_n292), .B2(new_n211), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n288), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n193), .A2(new_n223), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n295), .A2(new_n197), .ZN(new_n296));
  NOR3_X1   g110(.A1(new_n294), .A2(new_n195), .A3(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n217), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n298), .B1(new_n203), .B2(new_n225), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n287), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(G902), .B1(new_n286), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n282), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(G210), .B1(G237), .B2(G902), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n282), .A2(new_n303), .A3(new_n301), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n305), .A2(KEYINPUT89), .A3(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(G214), .B1(G237), .B2(G902), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n303), .B1(new_n282), .B2(new_n301), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT89), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n307), .A2(new_n308), .A3(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT90), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n312), .B(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G217), .ZN(new_n315));
  XOR2_X1   g129(.A(KEYINPUT74), .B(G902), .Z(new_n316));
  AOI21_X1  g130(.A(new_n315), .B1(new_n316), .B2(G234), .ZN(new_n317));
  NOR3_X1   g131(.A1(new_n268), .A2(KEYINPUT16), .A3(G140), .ZN(new_n318));
  XNOR2_X1  g132(.A(G125), .B(G140), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n318), .B1(new_n319), .B2(KEYINPUT16), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n320), .B(G146), .ZN(new_n321));
  XNOR2_X1  g135(.A(G119), .B(G128), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n322), .B(KEYINPUT75), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT24), .B(G110), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(G110), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n190), .A2(G128), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n328), .A2(KEYINPUT76), .ZN(new_n329));
  OAI21_X1  g143(.A(KEYINPUT23), .B1(new_n253), .B2(G119), .ZN(new_n330));
  OR2_X1    g144(.A1(KEYINPUT76), .A2(KEYINPUT23), .ZN(new_n331));
  AOI22_X1  g145(.A1(new_n329), .A2(new_n330), .B1(new_n328), .B2(new_n331), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n321), .B(new_n326), .C1(new_n327), .C2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n327), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n334), .B1(new_n323), .B2(new_n325), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n320), .A2(G146), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT77), .ZN(new_n337));
  INV_X1    g151(.A(G140), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G125), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n268), .A2(G140), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n337), .B1(new_n341), .B2(G146), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n319), .A2(KEYINPUT77), .A3(new_n255), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n335), .A2(new_n336), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n333), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g160(.A(KEYINPUT22), .B(G137), .ZN(new_n347));
  INV_X1    g161(.A(G953), .ZN(new_n348));
  AND3_X1   g162(.A1(new_n348), .A2(G221), .A3(G234), .ZN(new_n349));
  XOR2_X1   g163(.A(new_n347), .B(new_n349), .Z(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n346), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n333), .A2(new_n345), .A3(new_n350), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n352), .A2(new_n316), .A3(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT25), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n317), .B1(new_n356), .B2(KEYINPUT78), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  AND2_X1   g172(.A1(new_n352), .A2(new_n353), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n359), .A2(KEYINPUT25), .A3(new_n316), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n360), .A2(KEYINPUT78), .A3(new_n356), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n317), .A2(G902), .ZN(new_n362));
  AOI22_X1  g176(.A1(new_n358), .A2(new_n361), .B1(new_n362), .B2(new_n359), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT71), .ZN(new_n365));
  NOR2_X1   g179(.A1(G237), .A2(G953), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(G210), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n367), .B(KEYINPUT27), .ZN(new_n368));
  XNOR2_X1  g182(.A(KEYINPUT26), .B(G101), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n368), .B(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT11), .ZN(new_n371));
  INV_X1    g185(.A(G134), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n371), .B1(new_n372), .B2(G137), .ZN(new_n373));
  INV_X1    g187(.A(G137), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n374), .A2(KEYINPUT11), .A3(G134), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n372), .A2(G137), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n373), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(G131), .ZN(new_n378));
  INV_X1    g192(.A(G131), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n373), .A2(new_n375), .A3(new_n379), .A4(new_n376), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n374), .A2(KEYINPUT65), .A3(G134), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT65), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n383), .B1(new_n372), .B2(G137), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n374), .A2(G134), .ZN(new_n385));
  OAI211_X1 g199(.A(G131), .B(new_n382), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  AND2_X1   g200(.A1(new_n386), .A2(new_n380), .ZN(new_n387));
  AOI22_X1  g201(.A1(new_n381), .A2(new_n277), .B1(new_n387), .B2(new_n266), .ZN(new_n388));
  AND2_X1   g202(.A1(new_n239), .A2(new_n240), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NOR3_X1   g204(.A1(new_n388), .A2(new_n389), .A3(KEYINPUT69), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT69), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n277), .A2(new_n381), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n266), .A2(new_n380), .A3(new_n386), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n392), .B1(new_n395), .B2(new_n241), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n390), .B1(new_n391), .B2(new_n396), .ZN(new_n397));
  XOR2_X1   g211(.A(KEYINPUT68), .B(KEYINPUT28), .Z(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n395), .A2(new_n241), .ZN(new_n400));
  NOR3_X1   g214(.A1(new_n400), .A2(KEYINPUT70), .A3(KEYINPUT28), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT70), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT28), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n402), .B1(new_n390), .B2(new_n403), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n370), .B1(new_n399), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT30), .ZN(new_n407));
  AND3_X1   g221(.A1(new_n393), .A2(new_n394), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n407), .B1(new_n393), .B2(new_n394), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n241), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n410), .A2(new_n390), .A3(new_n370), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(KEYINPUT31), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT31), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n410), .A2(new_n413), .A3(new_n390), .A4(new_n370), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n365), .B1(new_n406), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n370), .ZN(new_n417));
  INV_X1    g231(.A(new_n398), .ZN(new_n418));
  OAI21_X1  g232(.A(KEYINPUT69), .B1(new_n388), .B2(new_n389), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n395), .A2(new_n392), .A3(new_n241), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n418), .B1(new_n421), .B2(new_n390), .ZN(new_n422));
  OAI21_X1  g236(.A(KEYINPUT70), .B1(new_n400), .B2(KEYINPUT28), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n390), .A2(new_n402), .A3(new_n403), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n417), .B1(new_n422), .B2(new_n425), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n426), .A2(KEYINPUT71), .A3(new_n412), .A4(new_n414), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n416), .A2(new_n427), .ZN(new_n428));
  NOR2_X1   g242(.A1(G472), .A2(G902), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  XNOR2_X1  g244(.A(KEYINPUT72), .B(KEYINPUT32), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n430), .A2(KEYINPUT73), .A3(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT73), .ZN(new_n434));
  INV_X1    g248(.A(new_n429), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n435), .B1(new_n416), .B2(new_n427), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n434), .B1(new_n436), .B2(new_n431), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n433), .A2(new_n437), .ZN(new_n438));
  AND2_X1   g252(.A1(new_n410), .A2(new_n390), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n417), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n395), .A2(new_n241), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n390), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n425), .B1(KEYINPUT28), .B2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT29), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n370), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NOR3_X1   g259(.A1(new_n422), .A2(new_n425), .A3(KEYINPUT29), .ZN(new_n446));
  OAI221_X1 g260(.A(new_n316), .B1(KEYINPUT29), .B2(new_n440), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  AOI22_X1  g261(.A1(new_n447), .A2(G472), .B1(new_n436), .B2(KEYINPUT32), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n364), .B1(new_n438), .B2(new_n448), .ZN(new_n449));
  XNOR2_X1  g263(.A(KEYINPUT9), .B(G234), .ZN(new_n450));
  OAI21_X1  g264(.A(G221), .B1(new_n450), .B2(G902), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(G902), .ZN(new_n453));
  XNOR2_X1  g267(.A(G143), .B(G146), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n259), .B1(new_n265), .B2(new_n454), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n455), .B(new_n211), .C1(new_n214), .C2(new_n216), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT10), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT82), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n456), .A2(KEYINPUT82), .A3(new_n457), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n274), .A2(new_n276), .ZN(new_n462));
  INV_X1    g276(.A(new_n271), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n235), .B1(new_n227), .B2(G101), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n211), .A2(KEYINPUT4), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n464), .B1(new_n467), .B2(new_n236), .ZN(new_n468));
  AOI22_X1  g282(.A1(new_n460), .A2(new_n461), .B1(new_n233), .B2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n381), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT84), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n266), .A2(KEYINPUT10), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n471), .B1(new_n221), .B2(new_n473), .ZN(new_n474));
  AOI211_X1 g288(.A(KEYINPUT84), .B(new_n472), .C1(new_n219), .C2(new_n220), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n469), .B(new_n470), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  NOR3_X1   g290(.A1(new_n288), .A2(new_n293), .A3(new_n266), .ZN(new_n477));
  INV_X1    g291(.A(new_n456), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n381), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(KEYINPUT12), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT12), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n481), .B(new_n381), .C1(new_n477), .C2(new_n478), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n476), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  XNOR2_X1  g297(.A(G110), .B(G140), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n348), .A2(G227), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n484), .B(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT85), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n474), .A2(new_n475), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n460), .A2(new_n461), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n468), .A2(new_n233), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n381), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n486), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n493), .A2(new_n476), .A3(new_n494), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n487), .A2(new_n488), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n488), .B1(new_n487), .B2(new_n495), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n453), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G469), .ZN(new_n499));
  INV_X1    g313(.A(G469), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n494), .B1(new_n493), .B2(new_n476), .ZN(new_n501));
  AND4_X1   g315(.A1(new_n476), .A2(new_n480), .A3(new_n482), .A4(new_n494), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n500), .B(new_n316), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(KEYINPUT86), .ZN(new_n504));
  INV_X1    g318(.A(new_n476), .ZN(new_n505));
  OAI21_X1  g319(.A(KEYINPUT84), .B1(new_n294), .B2(new_n472), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n221), .A2(new_n473), .A3(new_n471), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n470), .B1(new_n508), .B2(new_n469), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n486), .B1(new_n505), .B2(new_n509), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n476), .A2(new_n480), .A3(new_n482), .A4(new_n494), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT86), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n512), .A2(new_n513), .A3(new_n500), .A4(new_n316), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n504), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n452), .B1(new_n499), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT97), .ZN(new_n517));
  INV_X1    g331(.A(G478), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n518), .A2(KEYINPUT15), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(KEYINPUT13), .B1(new_n257), .B2(G128), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n521), .B1(new_n253), .B2(G143), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n257), .A2(KEYINPUT13), .A3(G128), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n372), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n257), .A2(G128), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n253), .A2(G143), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n525), .A2(new_n526), .A3(new_n372), .ZN(new_n527));
  INV_X1    g341(.A(G122), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(G116), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n188), .A2(G122), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n529), .A2(new_n530), .A3(new_n207), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n207), .B1(new_n529), .B2(new_n530), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n527), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OR2_X1    g348(.A1(new_n524), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n527), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n372), .B1(new_n525), .B2(new_n526), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n531), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(KEYINPUT14), .B1(new_n528), .B2(G116), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n528), .A2(G116), .ZN(new_n541));
  OAI21_X1  g355(.A(KEYINPUT95), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT95), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n188), .A2(G122), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n543), .B(new_n530), .C1(new_n544), .C2(KEYINPUT14), .ZN(new_n545));
  OR2_X1    g359(.A1(new_n530), .A2(KEYINPUT14), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n542), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(G107), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n539), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT96), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n535), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n538), .B1(G107), .B2(new_n547), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n524), .A2(new_n534), .ZN(new_n553));
  OAI21_X1  g367(.A(KEYINPUT96), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  NOR3_X1   g369(.A1(new_n450), .A2(new_n315), .A3(G953), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n551), .A2(new_n554), .A3(new_n556), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n520), .B1(new_n560), .B2(new_n316), .ZN(new_n561));
  INV_X1    g375(.A(new_n316), .ZN(new_n562));
  AOI211_X1 g376(.A(new_n562), .B(new_n519), .C1(new_n558), .C2(new_n559), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n517), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n559), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n556), .B1(new_n551), .B2(new_n554), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n316), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n519), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n560), .A2(new_n316), .A3(new_n520), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n568), .A2(new_n569), .A3(KEYINPUT97), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n564), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g385(.A1(G475), .A2(G902), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n572), .B(KEYINPUT94), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n320), .B(new_n255), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n366), .A2(G214), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n575), .A2(KEYINPUT91), .A3(new_n257), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n257), .A2(KEYINPUT91), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n577), .A2(G214), .A3(new_n366), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n579), .A2(KEYINPUT17), .A3(G131), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n575), .B(new_n577), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n379), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n579), .A2(G131), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n574), .B(new_n580), .C1(new_n584), .C2(KEYINPUT17), .ZN(new_n585));
  XNOR2_X1  g399(.A(G113), .B(G122), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(new_n204), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n341), .A2(G146), .ZN(new_n588));
  NAND2_X1  g402(.A1(KEYINPUT18), .A2(G131), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  AOI22_X1  g404(.A1(new_n344), .A2(new_n588), .B1(new_n590), .B2(new_n579), .ZN(new_n591));
  NOR3_X1   g405(.A1(new_n579), .A2(KEYINPUT92), .A3(new_n590), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT92), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n593), .B1(new_n581), .B2(new_n589), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n591), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  AND3_X1   g409(.A1(new_n585), .A2(new_n587), .A3(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT93), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT19), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n341), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n319), .A2(KEYINPUT19), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n597), .B1(new_n601), .B2(new_n255), .ZN(new_n602));
  AOI211_X1 g416(.A(KEYINPUT93), .B(G146), .C1(new_n599), .C2(new_n600), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n584), .B(new_n336), .C1(new_n602), .C2(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n587), .B1(new_n604), .B2(new_n595), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n573), .B1(new_n596), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(KEYINPUT20), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT20), .ZN(new_n608));
  OAI211_X1 g422(.A(new_n608), .B(new_n573), .C1(new_n596), .C2(new_n605), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n587), .B1(new_n585), .B2(new_n595), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n453), .B1(new_n596), .B2(new_n610), .ZN(new_n611));
  AOI22_X1  g425(.A1(new_n607), .A2(new_n609), .B1(G475), .B2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  AND2_X1   g427(.A1(new_n348), .A2(G952), .ZN(new_n614));
  INV_X1    g428(.A(G234), .ZN(new_n615));
  INV_X1    g429(.A(G237), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  AOI211_X1 g432(.A(new_n348), .B(new_n316), .C1(G234), .C2(G237), .ZN(new_n619));
  XNOR2_X1  g433(.A(KEYINPUT21), .B(G898), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NOR3_X1   g435(.A1(new_n571), .A2(new_n613), .A3(new_n621), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n516), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n314), .A2(new_n449), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(KEYINPUT98), .B(G101), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G3));
  NAND2_X1  g440(.A1(new_n428), .A2(new_n316), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(G472), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n430), .ZN(new_n629));
  AOI22_X1  g443(.A1(new_n498), .A2(G469), .B1(new_n504), .B2(new_n514), .ZN(new_n630));
  NOR4_X1   g444(.A1(new_n629), .A2(new_n630), .A3(new_n364), .A4(new_n452), .ZN(new_n631));
  AND3_X1   g445(.A1(new_n282), .A2(new_n303), .A3(new_n301), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n308), .B1(new_n632), .B2(new_n309), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT33), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n560), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n558), .A2(KEYINPUT33), .A3(new_n559), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n635), .A2(G478), .A3(new_n316), .A4(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n567), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n637), .B1(G478), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n613), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n633), .A2(new_n621), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n631), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(new_n204), .ZN(new_n643));
  XNOR2_X1  g457(.A(KEYINPUT99), .B(KEYINPUT34), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G6));
  NAND2_X1  g459(.A1(new_n305), .A2(new_n306), .ZN(new_n646));
  INV_X1    g460(.A(new_n621), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n613), .B1(new_n564), .B2(new_n570), .ZN(new_n648));
  AND4_X1   g462(.A1(new_n308), .A2(new_n646), .A3(new_n647), .A4(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n631), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT35), .B(G107), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G9));
  NOR2_X1   g466(.A1(new_n351), .A2(KEYINPUT36), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n346), .B(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n362), .ZN(new_n655));
  INV_X1    g469(.A(new_n361), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n655), .B1(new_n656), .B2(new_n357), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n629), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n314), .A2(new_n623), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT37), .B(G110), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G12));
  INV_X1    g476(.A(G900), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n618), .B1(new_n619), .B2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n648), .A2(new_n657), .A3(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n666), .B1(new_n438), .B2(new_n448), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n630), .A2(new_n452), .A3(new_n633), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G128), .ZN(G30));
  XOR2_X1   g484(.A(new_n664), .B(KEYINPUT39), .Z(new_n671));
  NAND2_X1  g485(.A1(new_n516), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(KEYINPUT100), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(KEYINPUT40), .ZN(new_n674));
  OR2_X1    g488(.A1(new_n672), .A2(KEYINPUT100), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT40), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n672), .A2(KEYINPUT100), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n307), .A2(new_n311), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(KEYINPUT38), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n439), .A2(new_n417), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n442), .ZN(new_n683));
  AOI21_X1  g497(.A(G902), .B1(new_n683), .B2(new_n417), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  AOI22_X1  g499(.A1(new_n436), .A2(KEYINPUT32), .B1(G472), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n438), .A2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n612), .B1(new_n564), .B2(new_n570), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n658), .A2(new_n308), .A3(new_n689), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n680), .A2(new_n688), .A3(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n674), .A2(new_n678), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G143), .ZN(G45));
  AOI21_X1  g507(.A(new_n658), .B1(new_n438), .B2(new_n448), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n639), .A2(new_n613), .A3(new_n665), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n694), .A2(new_n668), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G146), .ZN(G48));
  INV_X1    g512(.A(new_n512), .ZN(new_n699));
  OAI21_X1  g513(.A(G469), .B1(new_n699), .B2(new_n562), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n515), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n701), .A2(new_n452), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n449), .A2(new_n641), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(KEYINPUT41), .B(G113), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G15));
  NAND3_X1  g519(.A1(new_n449), .A2(new_n649), .A3(new_n702), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G116), .ZN(G18));
  NOR3_X1   g521(.A1(new_n701), .A2(new_n452), .A3(new_n633), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n694), .A2(new_n708), .A3(new_n622), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G119), .ZN(G21));
  OAI211_X1 g524(.A(new_n689), .B(new_n308), .C1(new_n632), .C2(new_n309), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT101), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n646), .A2(KEYINPUT101), .A3(new_n308), .A4(new_n689), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n443), .A2(new_n370), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n429), .B1(new_n716), .B2(new_n415), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n628), .A2(new_n363), .A3(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n715), .A2(new_n702), .A3(new_n719), .A4(new_n647), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G122), .ZN(G24));
  NAND3_X1  g535(.A1(new_n628), .A2(new_n657), .A3(new_n717), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n722), .A2(new_n695), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n708), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G125), .ZN(G27));
  INV_X1    g539(.A(KEYINPUT102), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n483), .A2(new_n726), .A3(new_n486), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n495), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n726), .B1(new_n483), .B2(new_n486), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n453), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(G469), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n452), .B1(new_n515), .B2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n308), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n733), .B1(new_n307), .B2(new_n311), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n436), .A2(KEYINPUT32), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n364), .B1(new_n448), .B2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT42), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n695), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n736), .A2(KEYINPUT103), .A3(new_n739), .A4(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT103), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n739), .A2(new_n741), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n743), .B1(new_n744), .B2(new_n735), .ZN(new_n745));
  AND2_X1   g559(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n736), .A2(new_n449), .A3(new_n696), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(new_n740), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G131), .ZN(G33));
  NAND4_X1  g564(.A1(new_n736), .A2(new_n449), .A3(new_n648), .A4(new_n665), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G134), .ZN(G36));
  NAND2_X1  g566(.A1(new_n639), .A2(new_n612), .ZN(new_n753));
  NAND2_X1  g567(.A1(KEYINPUT104), .A2(KEYINPUT43), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n639), .A2(new_n612), .A3(new_n756), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n658), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n629), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT44), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n758), .A2(KEYINPUT44), .A3(new_n629), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n761), .A2(new_n734), .A3(new_n762), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n500), .A2(new_n453), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n728), .A2(new_n729), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(KEYINPUT45), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(G469), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n496), .A2(new_n497), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n769), .A2(KEYINPUT45), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n765), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT46), .ZN(new_n772));
  AOI22_X1  g586(.A1(new_n771), .A2(new_n772), .B1(new_n514), .B2(new_n504), .ZN(new_n773));
  OAI211_X1 g587(.A(KEYINPUT46), .B(new_n765), .C1(new_n768), .C2(new_n770), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n452), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n763), .A2(new_n775), .A3(new_n671), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G137), .ZN(G39));
  NAND2_X1  g591(.A1(new_n438), .A2(new_n448), .ZN(new_n778));
  INV_X1    g592(.A(new_n734), .ZN(new_n779));
  NOR4_X1   g593(.A1(new_n778), .A2(new_n779), .A3(new_n363), .A4(new_n695), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n775), .A2(KEYINPUT47), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT47), .ZN(new_n782));
  AOI211_X1 g596(.A(new_n782), .B(new_n452), .C1(new_n773), .C2(new_n774), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n780), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G140), .ZN(G42));
  NAND3_X1  g599(.A1(new_n363), .A2(new_n308), .A3(new_n451), .ZN(new_n786));
  AOI211_X1 g600(.A(new_n753), .B(new_n786), .C1(new_n701), .C2(KEYINPUT49), .ZN(new_n787));
  OR2_X1    g601(.A1(new_n701), .A2(KEYINPUT49), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n680), .A2(new_n787), .A3(new_n688), .A4(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT53), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n624), .A2(new_n660), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n703), .A2(new_n706), .A3(new_n709), .A4(new_n720), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n568), .A2(new_n569), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n612), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n621), .B1(new_n640), .B2(new_n794), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n314), .A2(new_n631), .A3(new_n795), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n791), .A2(new_n792), .A3(new_n796), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n613), .A2(new_n793), .A3(new_n664), .ZN(new_n798));
  XOR2_X1   g612(.A(new_n798), .B(KEYINPUT105), .Z(new_n799));
  NAND4_X1  g613(.A1(new_n694), .A2(new_n516), .A3(new_n734), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n736), .A2(new_n723), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n751), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n802), .B1(new_n746), .B2(new_n748), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n655), .B(new_n665), .C1(new_n656), .C2(new_n357), .ZN(new_n804));
  AOI211_X1 g618(.A(new_n452), .B(new_n804), .C1(new_n515), .C2(new_n731), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n805), .A2(new_n687), .A3(new_n715), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n697), .A2(new_n669), .A3(new_n724), .A4(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(KEYINPUT52), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n797), .A2(new_n803), .A3(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT106), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n807), .A2(new_n810), .ZN(new_n811));
  AOI22_X1  g625(.A1(new_n668), .A2(new_n667), .B1(new_n708), .B2(new_n723), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n812), .A2(KEYINPUT106), .A3(new_n697), .A4(new_n806), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT52), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n790), .B1(new_n809), .B2(new_n814), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n811), .A2(KEYINPUT52), .A3(new_n813), .ZN(new_n816));
  OAI21_X1  g630(.A(KEYINPUT107), .B1(new_n816), .B2(new_n814), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n811), .A2(new_n813), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT52), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT107), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n811), .A2(KEYINPUT52), .A3(new_n813), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n797), .A2(new_n803), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n817), .A2(new_n823), .A3(new_n825), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n815), .B1(new_n826), .B2(new_n790), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(KEYINPUT54), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n826), .A2(new_n790), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n809), .A2(new_n790), .A3(new_n814), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n828), .B1(KEYINPUT54), .B2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT108), .ZN(new_n834));
  INV_X1    g648(.A(new_n702), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n835), .A2(new_n617), .A3(new_n779), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n836), .A2(new_n363), .A3(new_n688), .ZN(new_n837));
  OR3_X1    g651(.A1(new_n837), .A2(new_n613), .A3(new_n639), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n755), .A2(new_n757), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n719), .A2(new_n618), .A3(new_n839), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n841), .A2(new_n835), .A3(new_n308), .ZN(new_n842));
  AOI21_X1  g656(.A(KEYINPUT50), .B1(new_n842), .B2(new_n680), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n842), .A2(KEYINPUT50), .A3(new_n680), .ZN(new_n844));
  OAI221_X1 g658(.A(new_n838), .B1(new_n722), .B2(new_n840), .C1(new_n843), .C2(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n781), .A2(new_n783), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n515), .A2(new_n452), .A3(new_n700), .ZN(new_n847));
  AOI211_X1 g661(.A(new_n779), .B(new_n841), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n834), .B1(new_n845), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n849), .A2(KEYINPUT51), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n849), .A2(KEYINPUT51), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n836), .A2(new_n739), .A3(new_n839), .ZN(new_n852));
  XOR2_X1   g666(.A(new_n852), .B(KEYINPUT48), .Z(new_n853));
  INV_X1    g667(.A(new_n708), .ZN(new_n854));
  OAI221_X1 g668(.A(new_n614), .B1(new_n854), .B2(new_n841), .C1(new_n837), .C2(new_n640), .ZN(new_n855));
  OR2_X1    g669(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  NOR4_X1   g670(.A1(new_n833), .A2(new_n850), .A3(new_n851), .A4(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(G952), .A2(G953), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n789), .B1(new_n857), .B2(new_n858), .ZN(G75));
  NOR2_X1   g673(.A1(new_n348), .A2(G952), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT112), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n316), .A2(new_n303), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n832), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n250), .A2(new_n252), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT109), .ZN(new_n866));
  XOR2_X1   g680(.A(new_n281), .B(KEYINPUT55), .Z(new_n867));
  XNOR2_X1  g681(.A(new_n866), .B(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n868), .A2(KEYINPUT56), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n862), .B1(new_n864), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n830), .B1(new_n826), .B2(new_n790), .ZN(new_n871));
  INV_X1    g685(.A(new_n863), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n862), .B(new_n869), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n861), .B1(new_n870), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n820), .A2(new_n822), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n824), .B1(new_n876), .B2(KEYINPUT107), .ZN(new_n877));
  AOI21_X1  g691(.A(KEYINPUT53), .B1(new_n877), .B2(new_n823), .ZN(new_n878));
  OAI211_X1 g692(.A(KEYINPUT110), .B(new_n863), .C1(new_n878), .C2(new_n830), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT110), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n880), .B1(new_n871), .B2(new_n872), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT56), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n879), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(new_n868), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(KEYINPUT111), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT111), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n883), .A2(new_n886), .A3(new_n868), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n875), .B1(new_n885), .B2(new_n887), .ZN(G51));
  XNOR2_X1  g702(.A(new_n512), .B(KEYINPUT113), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n871), .B(KEYINPUT54), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n764), .B(KEYINPUT57), .Z(new_n891));
  OAI21_X1  g705(.A(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n768), .A2(new_n770), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT114), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n832), .A2(new_n562), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n860), .B1(new_n892), .B2(new_n895), .ZN(G54));
  OR2_X1    g710(.A1(new_n596), .A2(new_n605), .ZN(new_n897));
  AND2_X1   g711(.A1(KEYINPUT58), .A2(G475), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n832), .A2(new_n562), .A3(new_n897), .A4(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT115), .ZN(new_n900));
  OR2_X1    g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n899), .A2(new_n900), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n832), .A2(new_n562), .A3(new_n898), .ZN(new_n903));
  INV_X1    g717(.A(new_n897), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n860), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n901), .A2(new_n902), .A3(new_n905), .ZN(G60));
  AND2_X1   g720(.A1(new_n635), .A2(new_n636), .ZN(new_n907));
  XNOR2_X1  g721(.A(KEYINPUT116), .B(KEYINPUT59), .ZN(new_n908));
  NAND2_X1  g722(.A1(G478), .A2(G902), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n908), .B(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n861), .B1(new_n890), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n907), .B1(new_n833), .B2(new_n910), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n912), .A2(new_n913), .ZN(G63));
  INV_X1    g728(.A(new_n359), .ZN(new_n915));
  NAND2_X1  g729(.A1(G217), .A2(G902), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT60), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n915), .B1(new_n871), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(new_n861), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT117), .ZN(new_n920));
  INV_X1    g734(.A(new_n917), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n832), .A2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(new_n654), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n920), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NOR4_X1   g738(.A1(new_n871), .A2(new_n920), .A3(new_n923), .A4(new_n917), .ZN(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n919), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n922), .A2(KEYINPUT118), .A3(new_n915), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT118), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n918), .A2(new_n929), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n928), .A2(new_n930), .A3(KEYINPUT61), .A4(new_n861), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n871), .A2(new_n917), .ZN(new_n932));
  AOI21_X1  g746(.A(KEYINPUT117), .B1(new_n932), .B2(new_n654), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n933), .A2(new_n925), .ZN(new_n934));
  OAI22_X1  g748(.A1(new_n927), .A2(KEYINPUT61), .B1(new_n931), .B2(new_n934), .ZN(G66));
  OAI21_X1  g749(.A(G953), .B1(new_n620), .B2(new_n279), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT119), .ZN(new_n937));
  INV_X1    g751(.A(new_n797), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n937), .B1(new_n938), .B2(new_n348), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n866), .B1(G898), .B2(new_n348), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT120), .Z(new_n941));
  XNOR2_X1  g755(.A(new_n939), .B(new_n941), .ZN(G69));
  INV_X1    g756(.A(new_n784), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT123), .ZN(new_n944));
  INV_X1    g758(.A(new_n776), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n640), .A2(new_n794), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n449), .A2(new_n734), .A3(new_n946), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n673), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n944), .B1(new_n945), .B2(new_n948), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n776), .B(KEYINPUT123), .C1(new_n673), .C2(new_n947), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n943), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n812), .A2(new_n697), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n692), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(KEYINPUT122), .B1(new_n954), .B2(KEYINPUT62), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT122), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT62), .ZN(new_n957));
  AOI211_X1 g771(.A(new_n956), .B(new_n957), .C1(new_n692), .C2(new_n953), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n951), .B1(new_n955), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n692), .A2(new_n953), .A3(new_n957), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT121), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n960), .B(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n348), .B1(new_n959), .B2(new_n962), .ZN(new_n963));
  OR2_X1    g777(.A1(new_n408), .A2(new_n409), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(new_n601), .Z(new_n965));
  NAND2_X1  g779(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n776), .A2(new_n953), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT124), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n967), .B(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n751), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n775), .A2(new_n671), .ZN(new_n971));
  AND2_X1   g785(.A1(new_n715), .A2(new_n739), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n970), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n973), .A2(new_n784), .A3(new_n749), .ZN(new_n974));
  OAI21_X1  g788(.A(KEYINPUT125), .B1(new_n969), .B2(new_n974), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n967), .B(KEYINPUT124), .ZN(new_n976));
  AND3_X1   g790(.A1(new_n973), .A2(new_n784), .A3(new_n749), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT125), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n976), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n975), .A2(new_n979), .A3(new_n348), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n965), .B1(G900), .B2(G953), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT126), .ZN(new_n983));
  AND3_X1   g797(.A1(new_n966), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n983), .B1(new_n966), .B2(new_n982), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n348), .B1(G227), .B2(G900), .ZN(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(new_n987));
  NOR3_X1   g801(.A1(new_n984), .A2(new_n985), .A3(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(new_n982), .ZN(new_n989));
  INV_X1    g803(.A(new_n965), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n954), .A2(KEYINPUT62), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n991), .A2(new_n956), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n954), .A2(KEYINPUT122), .A3(KEYINPUT62), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n960), .B(KEYINPUT121), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n994), .A2(new_n995), .A3(new_n951), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n990), .B1(new_n996), .B2(new_n348), .ZN(new_n997));
  OAI21_X1  g811(.A(KEYINPUT126), .B1(new_n989), .B2(new_n997), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n966), .A2(new_n982), .A3(new_n983), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n986), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n988), .A2(new_n1000), .ZN(G72));
  NAND2_X1  g815(.A1(G472), .A2(G902), .ZN(new_n1002));
  XOR2_X1   g816(.A(new_n1002), .B(KEYINPUT63), .Z(new_n1003));
  NAND4_X1  g817(.A1(new_n827), .A2(new_n440), .A3(new_n682), .A4(new_n1003), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n975), .A2(new_n979), .A3(new_n797), .ZN(new_n1005));
  AND2_X1   g819(.A1(new_n1005), .A2(new_n1003), .ZN(new_n1006));
  OAI211_X1 g820(.A(new_n861), .B(new_n1004), .C1(new_n1006), .C2(new_n440), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1003), .B1(new_n996), .B2(new_n938), .ZN(new_n1008));
  INV_X1    g822(.A(KEYINPUT127), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n1010), .A2(new_n682), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1007), .B1(new_n1011), .B2(new_n1012), .ZN(G57));
endmodule


