//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 0 0 1 1 1 1 1 0 1 1 0 1 0 1 1 0 0 0 1 1 0 0 0 1 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 1 1 0 1 0 0 0 1 0 1 1 1 1 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:23 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1310, new_n1311, new_n1312, new_n1313, new_n1314,
    new_n1316, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1372, new_n1373, new_n1374, new_n1375, new_n1376;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(new_n204));
  XOR2_X1   g0004(.A(new_n204), .B(KEYINPUT64), .Z(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT65), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  AND2_X1   g0014(.A1(KEYINPUT66), .A2(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(KEYINPUT66), .A2(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G58), .ZN(new_n220));
  INV_X1    g0020(.A(G68), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(G50), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n219), .A2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(KEYINPUT67), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  AOI22_X1  g0030(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n231));
  AOI22_X1  g0031(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n232));
  NAND3_X1  g0032(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n228), .A2(new_n229), .ZN(new_n234));
  OAI21_X1  g0034(.A(new_n211), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  OAI211_X1 g0035(.A(new_n214), .B(new_n225), .C1(KEYINPUT1), .C2(new_n235), .ZN(new_n236));
  AOI21_X1  g0036(.A(new_n236), .B1(KEYINPUT1), .B2(new_n235), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XOR2_X1   g0039(.A(KEYINPUT2), .B(G226), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G264), .B(G270), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n241), .B(new_n245), .ZN(G358));
  XNOR2_X1  g0046(.A(G50), .B(G68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n247), .B(new_n248), .Z(new_n249));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XOR2_X1   g0050(.A(G107), .B(G116), .Z(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n249), .B(new_n252), .Z(G351));
  INV_X1    g0053(.A(G13), .ZN(new_n254));
  INV_X1    g0054(.A(G20), .ZN(new_n255));
  NOR3_X1   g0055(.A1(new_n254), .A2(new_n255), .A3(G1), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n256), .A2(G116), .ZN(new_n257));
  INV_X1    g0057(.A(new_n256), .ZN(new_n258));
  NAND3_X1  g0058(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(new_n218), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G1), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G33), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n258), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n257), .B1(new_n264), .B2(G116), .ZN(new_n265));
  NAND2_X1  g0065(.A1(G33), .A2(G283), .ZN(new_n266));
  INV_X1    g0066(.A(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G97), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n217), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT89), .ZN(new_n270));
  INV_X1    g0070(.A(G116), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G20), .ZN(new_n272));
  AND3_X1   g0072(.A1(new_n260), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n270), .B1(new_n260), .B2(new_n272), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n269), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT20), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  OAI211_X1 g0077(.A(KEYINPUT20), .B(new_n269), .C1(new_n273), .C2(new_n274), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n265), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT3), .B(G33), .ZN(new_n280));
  NOR2_X1   g0080(.A1(G257), .A2(G1698), .ZN(new_n281));
  INV_X1    g0081(.A(G1698), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(G264), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n280), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n218), .B1(G33), .B2(G41), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n267), .A2(KEYINPUT3), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT3), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G303), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n284), .A2(new_n285), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(G33), .A2(G41), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n218), .B1(KEYINPUT69), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT69), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n295), .A2(G33), .A3(G41), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g0097(.A(KEYINPUT5), .B(G41), .ZN(new_n298));
  INV_X1    g0098(.A(G45), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n299), .A2(G1), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n297), .A2(new_n301), .A3(G270), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n300), .A2(G274), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n297), .A2(new_n304), .A3(new_n298), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n292), .A2(new_n302), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G169), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(KEYINPUT21), .ZN(new_n309));
  AND3_X1   g0109(.A1(new_n292), .A2(new_n302), .A3(new_n305), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(G179), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n279), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n310), .A2(G190), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n306), .A2(G200), .ZN(new_n314));
  AND3_X1   g0114(.A1(new_n279), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n265), .ZN(new_n316));
  INV_X1    g0116(.A(new_n274), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n260), .A2(new_n270), .A3(new_n272), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(KEYINPUT20), .B1(new_n319), .B2(new_n269), .ZN(new_n320));
  INV_X1    g0120(.A(new_n278), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n316), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT90), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n322), .A2(new_n308), .A3(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(KEYINPUT90), .B1(new_n279), .B2(new_n307), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT21), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT91), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n324), .A2(new_n325), .A3(KEYINPUT91), .A4(new_n326), .ZN(new_n330));
  AOI211_X1 g0130(.A(new_n312), .B(new_n315), .C1(new_n329), .C2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n220), .A2(KEYINPUT8), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT8), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(G58), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n332), .A2(new_n334), .A3(KEYINPUT72), .ZN(new_n335));
  OR3_X1    g0135(.A1(new_n333), .A2(KEYINPUT72), .A3(G58), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(KEYINPUT73), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT73), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n335), .A2(new_n336), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n217), .A2(G33), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n338), .A2(new_n340), .A3(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT74), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n255), .A2(new_n267), .ZN(new_n345));
  INV_X1    g0145(.A(G150), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n343), .A2(new_n344), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n203), .A2(G20), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n344), .B1(new_n343), .B2(new_n348), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n260), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n258), .A2(G50), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n260), .B1(new_n262), .B2(G20), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n354), .B1(G50), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT71), .ZN(new_n358));
  INV_X1    g0158(.A(new_n285), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n280), .A2(G222), .A3(new_n282), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT70), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n280), .A2(KEYINPUT70), .A3(G222), .A4(new_n282), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n289), .A2(new_n282), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n365), .A2(G223), .B1(G77), .B2(new_n289), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n359), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(G41), .ZN(new_n368));
  AOI21_X1  g0168(.A(G1), .B1(new_n368), .B2(new_n299), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n369), .B1(new_n294), .B2(new_n296), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(G226), .ZN(new_n371));
  INV_X1    g0171(.A(G274), .ZN(new_n372));
  AOI211_X1 g0172(.A(G1), .B(new_n372), .C1(new_n368), .C2(new_n299), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n297), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n358), .B1(new_n367), .B2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n375), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n280), .A2(G1698), .ZN(new_n378));
  INV_X1    g0178(.A(G223), .ZN(new_n379));
  INV_X1    g0179(.A(G77), .ZN(new_n380));
  OAI22_X1  g0180(.A1(new_n378), .A2(new_n379), .B1(new_n380), .B2(new_n280), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n381), .B1(new_n362), .B2(new_n363), .ZN(new_n382));
  OAI211_X1 g0182(.A(KEYINPUT71), .B(new_n377), .C1(new_n382), .C2(new_n359), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n376), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n357), .B1(G169), .B2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(G179), .ZN(new_n386));
  AOI22_X1  g0186(.A1(new_n385), .A2(KEYINPUT75), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT75), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n357), .B(new_n388), .C1(G169), .C2(new_n384), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT10), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT9), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n392), .B1(new_n353), .B2(new_n356), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n353), .A2(new_n392), .A3(new_n356), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(G190), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n397), .B1(new_n376), .B2(new_n383), .ZN(new_n398));
  INV_X1    g0198(.A(new_n384), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n398), .B1(new_n399), .B2(G200), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n391), .B1(new_n396), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n395), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n400), .B(new_n391), .C1(new_n402), .C2(new_n393), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n390), .B1(new_n401), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(KEYINPUT7), .B1(new_n280), .B2(G20), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT7), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n289), .A2(new_n217), .A3(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n406), .A2(new_n408), .A3(G68), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT81), .ZN(new_n410));
  NAND2_X1  g0210(.A1(G58), .A2(G68), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n255), .B1(new_n222), .B2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(G159), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n345), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n410), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  AND2_X1   g0215(.A1(G58), .A2(G68), .ZN(new_n416));
  OAI21_X1  g0216(.A(G20), .B1(new_n416), .B2(new_n201), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n417), .B(KEYINPUT81), .C1(new_n413), .C2(new_n345), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n409), .A2(KEYINPUT16), .A3(new_n415), .A4(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n415), .A2(new_n418), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT82), .ZN(new_n421));
  AOI21_X1  g0221(.A(G20), .B1(new_n286), .B2(new_n288), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n421), .B1(new_n422), .B2(KEYINPUT7), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n289), .A2(new_n217), .A3(KEYINPUT7), .ZN(new_n424));
  OAI211_X1 g0224(.A(KEYINPUT82), .B(new_n407), .C1(new_n280), .C2(G20), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n420), .B1(new_n426), .B2(G68), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n260), .B(new_n419), .C1(new_n427), .C2(KEYINPUT16), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n338), .A2(new_n340), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n258), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n430), .B1(new_n429), .B2(new_n355), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n286), .A2(new_n288), .A3(G223), .A4(new_n282), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n286), .A2(new_n288), .A3(G226), .A4(G1698), .ZN(new_n433));
  INV_X1    g0233(.A(G87), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n432), .B(new_n433), .C1(new_n267), .C2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n285), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n370), .A2(G232), .B1(new_n297), .B2(new_n373), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n436), .A2(new_n437), .A3(new_n397), .ZN(new_n438));
  AND2_X1   g0238(.A1(new_n436), .A2(new_n437), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n438), .B1(new_n439), .B2(G200), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n428), .A2(new_n431), .A3(new_n440), .ZN(new_n441));
  XNOR2_X1  g0241(.A(new_n441), .B(KEYINPUT17), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n425), .A2(new_n424), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n287), .A2(G33), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n267), .A2(KEYINPUT3), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n255), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(KEYINPUT82), .B1(new_n446), .B2(new_n407), .ZN(new_n447));
  OAI21_X1  g0247(.A(G68), .B1(new_n443), .B2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n420), .ZN(new_n449));
  AOI21_X1  g0249(.A(KEYINPUT16), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n419), .A2(new_n260), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n431), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT18), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n439), .A2(G179), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n436), .A2(new_n437), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(G169), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  AND3_X1   g0257(.A1(new_n452), .A2(new_n453), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n453), .B1(new_n452), .B2(new_n457), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AND2_X1   g0260(.A1(new_n442), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n280), .A2(G232), .A3(G1698), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n280), .A2(G226), .A3(new_n282), .ZN(new_n463));
  NAND2_X1  g0263(.A1(G33), .A2(G97), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(new_n285), .ZN(new_n466));
  AOI22_X1  g0266(.A1(new_n374), .A2(KEYINPUT79), .B1(new_n370), .B2(G238), .ZN(new_n467));
  AND2_X1   g0267(.A1(new_n297), .A2(new_n373), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT79), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n466), .A2(new_n467), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(KEYINPUT13), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT13), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n466), .A2(new_n467), .A3(new_n470), .A4(new_n473), .ZN(new_n474));
  AND2_X1   g0274(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(G169), .ZN(new_n476));
  OAI21_X1  g0276(.A(KEYINPUT14), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n475), .A2(G179), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n472), .A2(new_n474), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT14), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n479), .A2(new_n480), .A3(G169), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n477), .A2(new_n478), .A3(new_n481), .ZN(new_n482));
  OAI22_X1  g0282(.A1(new_n341), .A2(new_n380), .B1(new_n255), .B2(G68), .ZN(new_n483));
  OAI22_X1  g0283(.A1(new_n483), .A2(KEYINPUT80), .B1(new_n202), .B2(new_n345), .ZN(new_n484));
  AND2_X1   g0284(.A1(new_n483), .A2(KEYINPUT80), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n260), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT11), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI211_X1 g0288(.A(KEYINPUT11), .B(new_n260), .C1(new_n484), .C2(new_n485), .ZN(new_n489));
  OR3_X1    g0289(.A1(new_n258), .A2(KEYINPUT12), .A3(G68), .ZN(new_n490));
  OAI21_X1  g0290(.A(KEYINPUT12), .B1(new_n258), .B2(G68), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n490), .A2(new_n491), .B1(G68), .B2(new_n355), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n488), .A2(new_n489), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n482), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n479), .A2(new_n397), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n495), .A2(new_n493), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n479), .A2(G200), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n280), .A2(G232), .A3(new_n282), .ZN(new_n499));
  INV_X1    g0299(.A(G238), .ZN(new_n500));
  OAI221_X1 g0300(.A(new_n499), .B1(new_n207), .B2(new_n280), .C1(new_n378), .C2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n285), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n468), .B1(G244), .B2(new_n370), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n386), .ZN(new_n506));
  INV_X1    g0306(.A(new_n217), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(G77), .ZN(new_n508));
  XNOR2_X1  g0308(.A(KEYINPUT15), .B(G87), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n332), .A2(new_n334), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT77), .ZN(new_n511));
  XNOR2_X1  g0311(.A(new_n510), .B(new_n511), .ZN(new_n512));
  OAI221_X1 g0312(.A(new_n508), .B1(new_n341), .B2(new_n509), .C1(new_n512), .C2(new_n345), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n260), .ZN(new_n514));
  OR3_X1    g0314(.A1(new_n258), .A2(KEYINPUT78), .A3(G77), .ZN(new_n515));
  OAI21_X1  g0315(.A(KEYINPUT78), .B1(new_n258), .B2(G77), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n515), .A2(new_n516), .B1(G77), .B2(new_n355), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n504), .A2(new_n476), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n506), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n505), .A2(KEYINPUT76), .A3(G190), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT76), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n523), .B1(new_n504), .B2(new_n397), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n518), .B1(G200), .B2(new_n504), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n521), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n461), .A2(new_n494), .A3(new_n498), .A4(new_n527), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n405), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n256), .A2(new_n206), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n530), .B1(new_n264), .B2(new_n206), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT84), .ZN(new_n532));
  AND2_X1   g0332(.A1(G97), .A2(G107), .ZN(new_n533));
  NOR2_X1   g0333(.A1(G97), .A2(G107), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT83), .ZN(new_n535));
  OAI22_X1  g0335(.A1(new_n533), .A2(new_n534), .B1(new_n535), .B2(KEYINPUT6), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n535), .A2(KEYINPUT6), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT6), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n538), .A2(G97), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(G97), .A2(G107), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n208), .A2(new_n541), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n532), .B(new_n536), .C1(new_n540), .C2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n208), .B(new_n541), .C1(new_n537), .C2(new_n539), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n532), .B1(new_n545), .B2(new_n536), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n507), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n426), .A2(G107), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n255), .A2(new_n267), .A3(G77), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n531), .B1(new_n550), .B2(new_n260), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n286), .A2(new_n288), .A3(G244), .A4(new_n282), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT4), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(KEYINPUT85), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n280), .A2(KEYINPUT4), .A3(G244), .A4(new_n282), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(KEYINPUT86), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT85), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n552), .A2(new_n558), .A3(new_n553), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n555), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n280), .A2(G250), .A3(G1698), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n266), .B(new_n561), .C1(new_n556), .C2(KEYINPUT86), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n285), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n296), .A2(new_n294), .B1(new_n298), .B2(new_n300), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(G257), .ZN(new_n565));
  AND2_X1   g0365(.A1(new_n565), .A2(new_n305), .ZN(new_n566));
  AND3_X1   g0366(.A1(new_n563), .A2(new_n386), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(G169), .B1(new_n563), .B2(new_n566), .ZN(new_n568));
  NOR3_X1   g0368(.A1(new_n551), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  AND3_X1   g0369(.A1(new_n563), .A2(new_n397), .A3(new_n566), .ZN(new_n570));
  AOI21_X1  g0370(.A(G200), .B1(new_n563), .B2(new_n566), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n551), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(KEYINPUT87), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT87), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n551), .B(new_n574), .C1(new_n570), .C2(new_n571), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n569), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT24), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n217), .A2(new_n280), .A3(G87), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(KEYINPUT22), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT22), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n217), .A2(new_n280), .A3(new_n580), .A4(G87), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g0382(.A1(KEYINPUT23), .A2(G107), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(new_n215), .B2(new_n216), .ZN(new_n584));
  NAND2_X1  g0384(.A1(G33), .A2(G116), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT23), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n255), .ZN(new_n588));
  NAND2_X1  g0388(.A1(KEYINPUT23), .A2(G107), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n584), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n577), .B1(new_n582), .B2(new_n591), .ZN(new_n592));
  AOI211_X1 g0392(.A(KEYINPUT24), .B(new_n590), .C1(new_n579), .C2(new_n581), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n260), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(new_n264), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT25), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(new_n258), .B2(G107), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n256), .A2(KEYINPUT25), .A3(new_n207), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n595), .A2(G107), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n594), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n280), .A2(G257), .A3(G1698), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n286), .A2(new_n288), .A3(G250), .A4(new_n282), .ZN(new_n602));
  NAND2_X1  g0402(.A1(G33), .A2(G294), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n285), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n564), .A2(G264), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n605), .A2(new_n606), .A3(new_n305), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(G169), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n608), .B(KEYINPUT92), .C1(new_n386), .C2(new_n607), .ZN(new_n609));
  OR3_X1    g0409(.A1(new_n607), .A2(KEYINPUT92), .A3(new_n386), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n600), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  OR2_X1    g0412(.A1(KEYINPUT66), .A2(G20), .ZN(new_n613));
  NAND2_X1  g0413(.A1(KEYINPUT66), .A2(G20), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n613), .A2(G33), .A3(G97), .A4(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT19), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n217), .A2(new_n280), .A3(G68), .ZN(new_n618));
  NAND3_X1  g0418(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n613), .A2(new_n614), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n534), .A2(new_n434), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n617), .A2(new_n618), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n260), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n595), .A2(G87), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n509), .A2(new_n256), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n286), .A2(new_n288), .A3(G244), .A4(G1698), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n286), .A2(new_n288), .A3(G238), .A4(new_n282), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n628), .A2(new_n629), .A3(new_n585), .ZN(new_n630));
  INV_X1    g0430(.A(G250), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n303), .B1(new_n300), .B2(new_n631), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n630), .A2(new_n285), .B1(new_n632), .B2(new_n297), .ZN(new_n633));
  INV_X1    g0433(.A(G200), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n627), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n633), .A2(KEYINPUT88), .A3(G190), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n633), .A2(G190), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT88), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n636), .A2(new_n637), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n630), .A2(new_n285), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n632), .A2(new_n297), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n642), .A2(new_n386), .A3(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(G169), .B1(new_n642), .B2(new_n643), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n624), .B(new_n626), .C1(new_n264), .C2(new_n509), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n641), .A2(new_n648), .ZN(new_n649));
  AOI22_X1  g0449(.A1(new_n604), .A2(new_n285), .B1(new_n564), .B2(G264), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n650), .A2(G190), .A3(new_n305), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n607), .A2(G200), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n594), .A2(new_n599), .A3(new_n651), .A4(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NOR3_X1   g0454(.A1(new_n612), .A2(new_n649), .A3(new_n654), .ZN(new_n655));
  AND4_X1   g0455(.A1(new_n331), .A2(new_n529), .A3(new_n576), .A4(new_n655), .ZN(G372));
  INV_X1    g0456(.A(new_n312), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n277), .A2(new_n278), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n307), .B1(new_n658), .B2(new_n316), .ZN(new_n659));
  AOI21_X1  g0459(.A(KEYINPUT21), .B1(new_n659), .B2(new_n323), .ZN(new_n660));
  AOI21_X1  g0460(.A(KEYINPUT91), .B1(new_n660), .B2(new_n325), .ZN(new_n661));
  AND4_X1   g0461(.A1(KEYINPUT91), .A2(new_n324), .A3(new_n325), .A4(new_n326), .ZN(new_n662));
  OAI211_X1 g0462(.A(new_n657), .B(new_n611), .C1(new_n661), .C2(new_n662), .ZN(new_n663));
  AOI22_X1  g0463(.A1(new_n636), .A2(new_n638), .B1(new_n646), .B2(new_n647), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n653), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n663), .A2(new_n576), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n550), .A2(new_n260), .ZN(new_n668));
  INV_X1    g0468(.A(new_n531), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n563), .A2(new_n386), .A3(new_n566), .ZN(new_n671));
  INV_X1    g0471(.A(new_n568), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(KEYINPUT26), .B1(new_n673), .B2(new_n649), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n551), .A2(new_n568), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT26), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n675), .A2(new_n676), .A3(new_n671), .A4(new_n664), .ZN(new_n677));
  AND3_X1   g0477(.A1(new_n674), .A2(new_n648), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n667), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n529), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g0480(.A(new_n680), .B(KEYINPUT93), .Z(new_n681));
  INV_X1    g0481(.A(KEYINPUT94), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n682), .B1(new_n458), .B2(new_n459), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n452), .A2(new_n457), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(KEYINPUT18), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n452), .A2(new_n453), .A3(new_n457), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(KEYINPUT94), .A3(new_n686), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  AOI22_X1  g0488(.A1(new_n498), .A2(new_n521), .B1(new_n482), .B2(new_n493), .ZN(new_n689));
  INV_X1    g0489(.A(new_n442), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n688), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n400), .B1(new_n402), .B2(new_n393), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(KEYINPUT10), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n403), .ZN(new_n694));
  AOI22_X1  g0494(.A1(new_n691), .A2(new_n694), .B1(new_n389), .B2(new_n387), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n681), .A2(new_n695), .ZN(G369));
  NAND3_X1  g0496(.A1(new_n217), .A2(new_n262), .A3(G13), .ZN(new_n697));
  OR2_X1    g0497(.A1(new_n697), .A2(KEYINPUT27), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(KEYINPUT27), .ZN(new_n699));
  AND3_X1   g0499(.A1(new_n698), .A2(G213), .A3(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(G343), .ZN(new_n702));
  OAI21_X1  g0502(.A(KEYINPUT95), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT95), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n700), .A2(new_n704), .A3(G343), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(new_n322), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n312), .B1(new_n329), .B2(new_n330), .ZN(new_n709));
  INV_X1    g0509(.A(new_n315), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT96), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n708), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n331), .A2(KEYINPUT96), .ZN(new_n714));
  AOI22_X1  g0514(.A1(new_n713), .A2(new_n714), .B1(new_n709), .B2(new_n708), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n706), .A2(new_n600), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n611), .B1(new_n716), .B2(new_n654), .ZN(new_n717));
  INV_X1    g0517(.A(new_n706), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n612), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n715), .A2(G330), .A3(new_n721), .ZN(new_n722));
  OR3_X1    g0522(.A1(new_n709), .A2(KEYINPUT97), .A3(new_n706), .ZN(new_n723));
  OAI21_X1  g0523(.A(KEYINPUT97), .B1(new_n709), .B2(new_n706), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n720), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n719), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n722), .A2(new_n727), .ZN(G399));
  INV_X1    g0528(.A(new_n212), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(G41), .ZN(new_n730));
  NOR4_X1   g0530(.A1(new_n730), .A2(new_n262), .A3(G116), .A4(new_n621), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n731), .B1(new_n224), .B2(new_n730), .ZN(new_n732));
  XOR2_X1   g0532(.A(new_n732), .B(KEYINPUT28), .Z(new_n733));
  INV_X1    g0533(.A(G330), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n331), .A2(new_n576), .A3(new_n655), .A4(new_n718), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT31), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n563), .A2(new_n566), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n310), .A2(new_n650), .A3(G179), .A4(new_n633), .ZN(new_n738));
  OAI21_X1  g0538(.A(KEYINPUT98), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n633), .ZN(new_n740));
  AND4_X1   g0540(.A1(new_n386), .A2(new_n607), .A3(new_n306), .A4(new_n740), .ZN(new_n741));
  AOI22_X1  g0541(.A1(new_n739), .A2(KEYINPUT30), .B1(new_n737), .B2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT30), .ZN(new_n743));
  OAI211_X1 g0543(.A(KEYINPUT98), .B(new_n743), .C1(new_n737), .C2(new_n738), .ZN(new_n744));
  AOI211_X1 g0544(.A(new_n736), .B(new_n718), .C1(new_n742), .C2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n739), .A2(KEYINPUT30), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n741), .A2(new_n737), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n746), .A2(new_n744), .A3(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(KEYINPUT31), .B1(new_n748), .B2(new_n706), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n734), .B1(new_n735), .B2(new_n750), .ZN(new_n751));
  XNOR2_X1  g0551(.A(KEYINPUT99), .B(KEYINPUT29), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n674), .A2(new_n648), .A3(new_n677), .ZN(new_n753));
  AOI211_X1 g0553(.A(new_n665), .B(new_n569), .C1(new_n573), .C2(new_n575), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n753), .B1(new_n754), .B2(new_n663), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n752), .B1(new_n755), .B2(new_n706), .ZN(new_n756));
  AND3_X1   g0556(.A1(new_n663), .A2(new_n576), .A3(new_n666), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n569), .A2(new_n676), .A3(new_n648), .A4(new_n641), .ZN(new_n758));
  INV_X1    g0558(.A(new_n664), .ZN(new_n759));
  OAI21_X1  g0559(.A(KEYINPUT26), .B1(new_n673), .B2(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n758), .A2(new_n760), .A3(new_n648), .ZN(new_n761));
  OAI211_X1 g0561(.A(KEYINPUT29), .B(new_n718), .C1(new_n757), .C2(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n751), .B1(new_n756), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n733), .B1(new_n763), .B2(G1), .ZN(G364));
  NOR2_X1   g0564(.A1(new_n507), .A2(new_n254), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G45), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G1), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n730), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n768), .B1(new_n715), .B2(G330), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n715), .A2(G330), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n715), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G13), .A2(G33), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(G20), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n212), .A2(new_n280), .ZN(new_n777));
  INV_X1    g0577(.A(G355), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n777), .A2(new_n778), .B1(G116), .B2(new_n212), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n729), .A2(new_n280), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n781), .B1(new_n299), .B2(new_n224), .ZN(new_n782));
  OR2_X1    g0582(.A1(new_n249), .A2(new_n299), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n779), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n218), .B1(G20), .B2(new_n476), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n786), .B1(G20), .B2(new_n774), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n768), .B1(new_n784), .B2(new_n787), .ZN(new_n788));
  NOR3_X1   g0588(.A1(G179), .A2(G190), .A3(G200), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n507), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n413), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT32), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR3_X1   g0593(.A1(new_n397), .A2(G179), .A3(G200), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n217), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(G97), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n793), .A2(new_n280), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n507), .A2(G179), .ZN(new_n799));
  NOR3_X1   g0599(.A1(new_n799), .A2(new_n397), .A3(G200), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n801), .A2(new_n220), .B1(new_n792), .B2(new_n791), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n386), .A2(G200), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n803), .B(KEYINPUT102), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(new_n397), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n805), .A2(new_n217), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n798), .B(new_n802), .C1(G107), .C2(new_n806), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n804), .A2(G20), .A3(G190), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT103), .ZN(new_n809));
  OR2_X1    g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n808), .A2(new_n809), .ZN(new_n811));
  AND2_X1   g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n507), .A2(G179), .A3(new_n397), .A4(new_n634), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n813), .A2(KEYINPUT100), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n813), .A2(KEYINPUT100), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  AOI22_X1  g0617(.A1(G87), .A2(new_n812), .B1(new_n817), .B2(G77), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT101), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(new_n799), .B2(new_n634), .ZN(new_n820));
  NAND4_X1  g0620(.A1(new_n507), .A2(KEYINPUT101), .A3(G179), .A4(G200), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n822), .A2(new_n397), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n822), .A2(G190), .ZN(new_n824));
  AOI22_X1  g0624(.A1(G50), .A2(new_n823), .B1(new_n824), .B2(G68), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n807), .A2(new_n818), .A3(new_n825), .ZN(new_n826));
  AOI22_X1  g0626(.A1(G303), .A2(new_n812), .B1(new_n817), .B2(G311), .ZN(new_n827));
  INV_X1    g0627(.A(new_n790), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(G329), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n280), .B1(new_n796), .B2(G294), .ZN(new_n830));
  INV_X1    g0630(.A(G322), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n829), .B(new_n830), .C1(new_n801), .C2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n832), .B1(G283), .B2(new_n806), .ZN(new_n833));
  XNOR2_X1  g0633(.A(KEYINPUT33), .B(G317), .ZN(new_n834));
  AOI22_X1  g0634(.A1(G326), .A2(new_n823), .B1(new_n824), .B2(new_n834), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n827), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n826), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n788), .B1(new_n837), .B2(new_n785), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n769), .A2(new_n771), .B1(new_n776), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(G396));
  AOI21_X1  g0640(.A(new_n706), .B1(new_n667), .B2(new_n678), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n520), .A2(new_n706), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n526), .A2(new_n525), .B1(new_n518), .B2(new_n706), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n843), .B1(new_n844), .B2(new_n521), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n841), .B(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n751), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  XOR2_X1   g0649(.A(new_n849), .B(KEYINPUT106), .Z(new_n850));
  AOI21_X1  g0650(.A(new_n768), .B1(new_n847), .B2(new_n848), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n785), .A2(new_n773), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n768), .B1(G77), .B2(new_n854), .ZN(new_n855));
  XOR2_X1   g0655(.A(new_n855), .B(KEYINPUT104), .Z(new_n856));
  INV_X1    g0656(.A(new_n806), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n857), .A2(new_n434), .ZN(new_n858));
  INV_X1    g0658(.A(G311), .ZN(new_n859));
  INV_X1    g0659(.A(G294), .ZN(new_n860));
  OAI221_X1 g0660(.A(new_n797), .B1(new_n859), .B2(new_n790), .C1(new_n801), .C2(new_n860), .ZN(new_n861));
  AOI211_X1 g0661(.A(new_n858), .B(new_n861), .C1(G116), .C2(new_n817), .ZN(new_n862));
  INV_X1    g0662(.A(G283), .ZN(new_n863));
  INV_X1    g0663(.A(new_n824), .ZN(new_n864));
  INV_X1    g0664(.A(new_n823), .ZN(new_n865));
  OAI221_X1 g0665(.A(new_n862), .B1(new_n863), .B2(new_n864), .C1(new_n290), .C2(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n280), .B1(new_n812), .B2(G107), .ZN(new_n867));
  XOR2_X1   g0667(.A(new_n867), .B(KEYINPUT105), .Z(new_n868));
  NOR2_X1   g0668(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  AOI22_X1  g0669(.A1(new_n817), .A2(G159), .B1(G143), .B2(new_n800), .ZN(new_n870));
  INV_X1    g0670(.A(G137), .ZN(new_n871));
  OAI221_X1 g0671(.A(new_n870), .B1(new_n871), .B2(new_n865), .C1(new_n346), .C2(new_n864), .ZN(new_n872));
  XNOR2_X1  g0672(.A(new_n872), .B(KEYINPUT34), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n806), .A2(G68), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n289), .B1(new_n796), .B2(G58), .ZN(new_n875));
  INV_X1    g0675(.A(G132), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n874), .B(new_n875), .C1(new_n876), .C2(new_n790), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n877), .B1(G50), .B2(new_n812), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n869), .B1(new_n873), .B2(new_n878), .ZN(new_n879));
  OAI221_X1 g0679(.A(new_n856), .B1(new_n846), .B2(new_n774), .C1(new_n786), .C2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n852), .A2(new_n880), .ZN(G384));
  NOR2_X1   g0681(.A1(new_n544), .A2(new_n546), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  OR2_X1    g0683(.A1(new_n883), .A2(KEYINPUT35), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(KEYINPUT35), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n884), .A2(new_n885), .A3(G116), .A4(new_n219), .ZN(new_n886));
  XOR2_X1   g0686(.A(new_n886), .B(KEYINPUT36), .Z(new_n887));
  NAND3_X1  g0687(.A1(new_n224), .A2(G77), .A3(new_n411), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n202), .A2(G68), .ZN(new_n889));
  AOI211_X1 g0689(.A(new_n262), .B(G13), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n735), .A2(new_n750), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n493), .A2(new_n706), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n494), .A2(new_n498), .A3(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n482), .A2(new_n493), .A3(new_n706), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n845), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n892), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT37), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT16), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n449), .A2(new_n409), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n451), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n431), .ZN(new_n902));
  OAI22_X1  g0702(.A1(new_n901), .A2(new_n902), .B1(new_n457), .B2(new_n700), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n898), .B1(new_n903), .B2(new_n441), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  AND3_X1   g0705(.A1(new_n428), .A2(new_n431), .A3(new_n440), .ZN(new_n906));
  AOI22_X1  g0706(.A1(new_n428), .A2(new_n431), .B1(new_n456), .B2(new_n454), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(KEYINPUT37), .B1(new_n452), .B2(new_n700), .ZN(new_n909));
  AOI21_X1  g0709(.A(KEYINPUT107), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n909), .A2(KEYINPUT107), .A3(new_n684), .A4(new_n441), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n905), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n442), .A2(new_n460), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n700), .B1(new_n901), .B2(new_n902), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n913), .A2(new_n917), .A3(KEYINPUT38), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT38), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n452), .A2(new_n700), .ZN(new_n920));
  NAND4_X1  g0720(.A1(new_n684), .A2(new_n920), .A3(new_n898), .A4(new_n441), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT107), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n904), .B1(new_n923), .B2(new_n911), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n915), .B1(new_n442), .B2(new_n460), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n919), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT108), .ZN(new_n927));
  AND3_X1   g0727(.A1(new_n918), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n927), .B1(new_n918), .B2(new_n926), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n897), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT40), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n892), .A2(new_n896), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n442), .A2(new_n683), .A3(new_n687), .ZN(new_n934));
  INV_X1    g0734(.A(new_n920), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n684), .A2(new_n441), .ZN(new_n937));
  OAI21_X1  g0737(.A(KEYINPUT37), .B1(new_n937), .B2(new_n935), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n910), .B2(new_n912), .ZN(new_n939));
  AOI21_X1  g0739(.A(KEYINPUT38), .B1(new_n936), .B2(new_n939), .ZN(new_n940));
  NOR3_X1   g0740(.A1(new_n924), .A2(new_n925), .A3(new_n919), .ZN(new_n941));
  OAI21_X1  g0741(.A(KEYINPUT40), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n932), .B1(new_n933), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n529), .A2(new_n892), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(G330), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n946), .B1(new_n943), .B2(new_n944), .ZN(new_n947));
  AOI21_X1  g0747(.A(KEYINPUT38), .B1(new_n913), .B2(new_n917), .ZN(new_n948));
  OAI21_X1  g0748(.A(KEYINPUT108), .B1(new_n948), .B2(new_n941), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n918), .A2(new_n926), .A3(new_n927), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n894), .A2(new_n895), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n841), .A2(new_n846), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n953), .B1(new_n954), .B2(new_n843), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n951), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT39), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n940), .B2(new_n941), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT109), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n494), .B2(new_n706), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n482), .A2(KEYINPUT109), .A3(new_n493), .A4(new_n718), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n918), .A2(new_n926), .A3(KEYINPUT39), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n958), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n688), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n701), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n956), .A2(new_n964), .A3(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n756), .A2(new_n529), .A3(new_n762), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n695), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n967), .B(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n947), .A2(new_n971), .B1(new_n262), .B2(new_n765), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n947), .A2(new_n971), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n891), .B1(new_n972), .B2(new_n973), .ZN(G367));
  NAND2_X1  g0774(.A1(new_n723), .A2(new_n724), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n721), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n723), .A2(new_n720), .A3(new_n724), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n772), .B2(new_n734), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n976), .A2(new_n715), .A3(G330), .A4(new_n977), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n979), .A2(new_n763), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n976), .A2(new_n719), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n706), .A2(new_n670), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n576), .A2(new_n983), .B1(new_n569), .B2(new_n706), .ZN(new_n984));
  AOI21_X1  g0784(.A(KEYINPUT44), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  OAI211_X1 g0785(.A(KEYINPUT44), .B(new_n984), .C1(new_n725), .C2(new_n726), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n984), .ZN(new_n988));
  AOI21_X1  g0788(.A(KEYINPUT45), .B1(new_n727), .B2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT45), .ZN(new_n990));
  NOR4_X1   g0790(.A1(new_n725), .A2(new_n990), .A3(new_n726), .A4(new_n984), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n985), .A2(new_n987), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n722), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n981), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n722), .B1(new_n989), .B2(new_n991), .C1(new_n985), .C2(new_n987), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n763), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n730), .B(KEYINPUT41), .Z(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n767), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  OR3_X1    g0800(.A1(new_n722), .A2(KEYINPUT110), .A3(new_n984), .ZN(new_n1001));
  OAI21_X1  g0801(.A(KEYINPUT110), .B1(new_n722), .B2(new_n984), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n706), .A2(new_n627), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n1004), .A2(new_n648), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n664), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1007), .A2(KEYINPUT43), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1003), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1001), .A2(new_n1008), .A3(new_n1002), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n573), .A2(new_n575), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(new_n612), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n706), .B1(new_n1014), .B2(new_n673), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n725), .A2(new_n988), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1015), .B1(new_n1016), .B2(KEYINPUT42), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(KEYINPUT42), .B2(new_n1016), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1007), .A2(KEYINPUT43), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1012), .A2(new_n1020), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1010), .A2(new_n1019), .A3(new_n1018), .A4(new_n1011), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n823), .A2(G143), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n805), .A2(new_n508), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n1025), .A2(new_n289), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT111), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n796), .A2(G68), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n871), .B2(new_n790), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(G150), .B2(new_n800), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1024), .A2(new_n1028), .A3(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(G159), .B2(new_n824), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(G58), .A2(new_n812), .B1(new_n817), .B2(G50), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n1033), .B(new_n1034), .C1(new_n1027), .C2(new_n1026), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n812), .A2(G116), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT46), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n857), .A2(new_n206), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n280), .B1(new_n828), .B2(G317), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1039), .B1(new_n207), .B2(new_n795), .C1(new_n801), .C2(new_n290), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n1038), .B(new_n1040), .C1(G283), .C2(new_n817), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(G294), .A2(new_n824), .B1(new_n823), .B2(G311), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1037), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  AND2_X1   g0843(.A1(new_n1035), .A2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n785), .B1(new_n1044), .B2(KEYINPUT47), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(KEYINPUT47), .B2(new_n1044), .ZN(new_n1046));
  AND2_X1   g0846(.A1(new_n245), .A2(new_n780), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n786), .B1(G20), .B2(new_n774), .C1(new_n212), .C2(new_n509), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n775), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n768), .B1(new_n1047), .B2(new_n1048), .C1(new_n1007), .C2(new_n1049), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n1000), .A2(new_n1023), .B1(new_n1046), .B2(new_n1050), .ZN(G387));
  NAND2_X1  g0851(.A1(new_n979), .A2(new_n980), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n763), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  OR2_X1    g0854(.A1(new_n1054), .A2(KEYINPUT113), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1054), .A2(KEYINPUT113), .ZN(new_n1056));
  NAND4_X1  g0856(.A1(new_n1055), .A2(new_n730), .A3(new_n981), .A4(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n767), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1052), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n812), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n1060), .A2(new_n860), .B1(new_n863), .B2(new_n795), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n817), .A2(G303), .B1(G317), .B2(new_n800), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1062), .B1(new_n859), .B2(new_n864), .C1(new_n831), .C2(new_n865), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT48), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1061), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n1064), .B2(new_n1063), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT49), .ZN(new_n1067));
  OR2_X1    g0867(.A1(new_n1067), .A2(KEYINPUT112), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n280), .B1(new_n828), .B2(G326), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n857), .B2(new_n271), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n1067), .B2(KEYINPUT112), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n812), .A2(G77), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n817), .A2(G68), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n801), .A2(new_n202), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n280), .B1(new_n795), .B2(new_n509), .C1(new_n790), .C2(new_n346), .ZN(new_n1076));
  NOR4_X1   g0876(.A1(new_n1074), .A2(new_n1038), .A3(new_n1075), .A4(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n429), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(G159), .A2(new_n823), .B1(new_n824), .B2(new_n1078), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n1068), .A2(new_n1071), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1080));
  OR2_X1    g0880(.A1(new_n1080), .A2(new_n786), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n621), .A2(G116), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n777), .A2(new_n1082), .B1(G107), .B2(new_n212), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n512), .A2(G50), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT50), .ZN(new_n1085));
  AOI21_X1  g0885(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1085), .A2(new_n1082), .A3(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n781), .B1(new_n241), .B2(G45), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1083), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n768), .B1(new_n1089), .B2(new_n787), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(new_n720), .B2(new_n775), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1059), .B1(new_n1081), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1057), .A2(new_n1092), .ZN(G393));
  NAND2_X1  g0893(.A1(new_n992), .A2(new_n993), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT114), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1094), .A2(new_n995), .A3(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n992), .A2(KEYINPUT114), .A3(new_n993), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1096), .A2(new_n981), .A3(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1098), .A2(new_n730), .A3(new_n996), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n780), .A2(new_n252), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n787), .B1(new_n729), .B2(G97), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  AND2_X1   g0902(.A1(new_n828), .A2(G143), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n795), .A2(new_n380), .ZN(new_n1104));
  NOR4_X1   g0904(.A1(new_n858), .A2(new_n289), .A3(new_n1103), .A4(new_n1104), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n1105), .B1(new_n221), .B2(new_n1060), .C1(new_n512), .C2(new_n816), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(G50), .B2(new_n824), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n823), .A2(G150), .B1(G159), .B2(new_n800), .ZN(new_n1108));
  XOR2_X1   g0908(.A(new_n1108), .B(KEYINPUT51), .Z(new_n1109));
  AOI22_X1  g0909(.A1(new_n823), .A2(G317), .B1(G311), .B2(new_n800), .ZN(new_n1110));
  XOR2_X1   g0910(.A(new_n1110), .B(KEYINPUT52), .Z(new_n1111));
  OAI221_X1 g0911(.A(new_n289), .B1(new_n795), .B2(new_n271), .C1(new_n790), .C2(new_n831), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(G107), .B2(new_n806), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n1113), .B1(new_n860), .B2(new_n816), .C1(new_n1060), .C2(new_n863), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(G303), .B2(new_n824), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n1107), .A2(new_n1109), .B1(new_n1111), .B2(new_n1115), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n768), .B(new_n1102), .C1(new_n1116), .C2(new_n786), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(new_n984), .B2(new_n775), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1118), .B1(new_n1119), .B2(new_n767), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1099), .A2(new_n1120), .ZN(G390));
  NAND2_X1  g0921(.A1(new_n529), .A2(new_n751), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n968), .A2(new_n695), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(KEYINPUT115), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT115), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n968), .A2(new_n695), .A3(new_n1125), .A4(new_n1122), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  AND4_X1   g0927(.A1(G330), .A2(new_n892), .A3(new_n846), .A4(new_n952), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n706), .B(new_n845), .C1(new_n667), .C2(new_n678), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n952), .B1(new_n1129), .B2(new_n842), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n962), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n1130), .A2(new_n1131), .B1(new_n958), .B2(new_n963), .ZN(new_n1132));
  OR2_X1    g0932(.A1(new_n844), .A2(new_n521), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n718), .B(new_n1133), .C1(new_n757), .C2(new_n761), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n953), .B1(new_n1134), .B2(new_n843), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1131), .B1(new_n940), .B2(new_n941), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1128), .B1(new_n1132), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n842), .B1(new_n841), .B2(new_n846), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1131), .B1(new_n1139), .B2(new_n953), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n958), .A2(new_n963), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n751), .A2(new_n846), .A3(new_n952), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n936), .A2(new_n939), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n919), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n962), .B1(new_n1145), .B2(new_n918), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n761), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n706), .B1(new_n1147), .B2(new_n667), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n842), .B1(new_n1148), .B2(new_n1133), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1146), .B1(new_n953), .B2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1142), .A2(new_n1143), .A3(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1139), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n952), .B1(new_n751), .B2(new_n846), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1152), .B1(new_n1128), .B2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n892), .A2(G330), .A3(new_n846), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(new_n953), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1156), .A2(new_n1143), .A3(new_n1149), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1154), .A2(new_n1157), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1127), .A2(new_n1138), .A3(new_n1151), .A4(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1158), .A2(new_n1126), .A3(new_n1124), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1143), .B1(new_n1142), .B2(new_n1150), .ZN(new_n1161));
  NOR3_X1   g0961(.A1(new_n1132), .A2(new_n1137), .A3(new_n1128), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1160), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1159), .A2(new_n1163), .A3(new_n730), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1141), .A2(new_n773), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n768), .B1(new_n1078), .B2(new_n854), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n864), .A2(new_n207), .B1(new_n206), .B2(new_n816), .ZN(new_n1167));
  OR2_X1    g0967(.A1(new_n1167), .A2(KEYINPUT117), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(KEYINPUT117), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n823), .A2(G283), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n280), .B(new_n1104), .C1(G294), .C2(new_n828), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1171), .B(new_n874), .C1(new_n271), .C2(new_n801), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(G87), .B2(new_n812), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .A4(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n812), .A2(G150), .ZN(new_n1175));
  XOR2_X1   g0975(.A(new_n1175), .B(KEYINPUT53), .Z(new_n1176));
  XNOR2_X1  g0976(.A(KEYINPUT54), .B(G143), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n817), .A2(new_n1178), .B1(new_n824), .B2(G137), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(KEYINPUT116), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n857), .A2(new_n202), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n289), .B1(new_n828), .B2(G125), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n1182), .B1(new_n413), .B2(new_n795), .C1(new_n801), .C2(new_n876), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n1181), .B(new_n1183), .C1(G128), .C2(new_n823), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1176), .A2(new_n1180), .A3(new_n1184), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1179), .A2(KEYINPUT116), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1174), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT118), .ZN(new_n1188));
  OR2_X1    g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n786), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1166), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1165), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1138), .A2(new_n1151), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1192), .B1(new_n1193), .B2(new_n1058), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  AND3_X1   g0995(.A1(new_n1164), .A2(new_n1195), .A3(KEYINPUT119), .ZN(new_n1196));
  AOI21_X1  g0996(.A(KEYINPUT119), .B1(new_n1164), .B2(new_n1195), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1196), .A2(new_n1197), .ZN(G378));
  NOR2_X1   g0998(.A1(new_n280), .A2(G41), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(G33), .A2(G41), .ZN(new_n1200));
  NOR3_X1   g1000(.A1(new_n1199), .A2(G50), .A3(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n806), .A2(G58), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1029), .B(new_n1199), .C1(new_n863), .C2(new_n790), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(G107), .B2(new_n800), .ZN(new_n1204));
  AND3_X1   g1004(.A1(new_n1072), .A2(new_n1202), .A3(new_n1204), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n864), .A2(new_n206), .B1(new_n509), .B2(new_n816), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT120), .ZN(new_n1207));
  AND2_X1   g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1205), .B1(new_n271), .B2(new_n865), .C1(new_n1208), .C2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT58), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1201), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1212), .B1(new_n1211), .B2(new_n1210), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n812), .A2(new_n1178), .ZN(new_n1214));
  XOR2_X1   g1014(.A(new_n1214), .B(KEYINPUT121), .Z(new_n1215));
  INV_X1    g1015(.A(KEYINPUT59), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n823), .A2(G125), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n800), .A2(G128), .B1(G150), .B2(new_n796), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n1217), .B(new_n1218), .C1(new_n871), .C2(new_n816), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(G132), .B2(new_n824), .ZN(new_n1220));
  AND3_X1   g1020(.A1(new_n1215), .A2(new_n1216), .A3(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1216), .B1(new_n1215), .B2(new_n1220), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n828), .A2(G124), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1200), .B(new_n1223), .C1(new_n857), .C2(new_n413), .ZN(new_n1224));
  NOR3_X1   g1024(.A1(new_n1221), .A2(new_n1222), .A3(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n785), .B1(new_n1213), .B2(new_n1225), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(new_n1226), .B(KEYINPUT122), .ZN(new_n1227));
  XOR2_X1   g1027(.A(KEYINPUT123), .B(KEYINPUT56), .Z(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n357), .A2(new_n700), .ZN(new_n1230));
  OR2_X1    g1030(.A1(new_n1230), .A2(KEYINPUT55), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(KEYINPUT55), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n694), .A2(new_n390), .A3(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1233), .B1(new_n694), .B2(new_n390), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1229), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1236), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1238), .A2(new_n1228), .A3(new_n1234), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1237), .A2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(new_n773), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n853), .A2(new_n202), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1227), .A2(new_n1241), .A3(new_n768), .A4(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT124), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n951), .A2(new_n955), .B1(new_n965), .B2(new_n701), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1245), .B1(new_n1246), .B2(new_n964), .ZN(new_n1247));
  AOI21_X1  g1047(.A(KEYINPUT40), .B1(new_n951), .B2(new_n897), .ZN(new_n1248));
  OAI21_X1  g1048(.A(G330), .B1(new_n942), .B2(new_n933), .ZN(new_n1249));
  NOR3_X1   g1049(.A1(new_n1248), .A2(new_n1249), .A3(new_n1240), .ZN(new_n1250));
  AND2_X1   g1050(.A1(new_n1237), .A2(new_n1239), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n931), .B1(new_n1145), .B2(new_n918), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n734), .B1(new_n1252), .B2(new_n897), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1251), .B1(new_n932), .B2(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1247), .B1(new_n1250), .B2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n967), .A2(KEYINPUT124), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n932), .A2(new_n1253), .A3(new_n1251), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1240), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1256), .A2(new_n1257), .A3(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1255), .A2(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1244), .B1(new_n1260), .B2(new_n767), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n967), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1262), .B1(new_n1250), .B2(new_n1254), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1258), .A2(new_n1257), .A3(new_n967), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1263), .A2(KEYINPUT57), .A3(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1162), .A2(new_n1161), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1266), .B1(new_n1267), .B2(new_n1158), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n730), .B1(new_n1265), .B2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1158), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1127), .B1(new_n1193), .B2(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(KEYINPUT57), .B1(new_n1260), .B2(new_n1271), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1261), .B1(new_n1269), .B2(new_n1272), .ZN(G375));
  NAND2_X1  g1073(.A1(new_n953), .A2(new_n773), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n768), .B1(G68), .B2(new_n854), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n790), .A2(new_n290), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n795), .A2(new_n509), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1278), .B1(new_n801), .B2(new_n863), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1279), .B1(new_n817), .B2(G107), .ZN(new_n1280));
  OAI221_X1 g1080(.A(new_n1280), .B1(new_n271), .B2(new_n864), .C1(new_n860), .C2(new_n865), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1025), .A2(new_n280), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(KEYINPUT125), .ZN(new_n1283));
  OR2_X1    g1083(.A1(new_n1282), .A2(KEYINPUT125), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1283), .B(new_n1284), .C1(new_n1060), .C2(new_n206), .ZN(new_n1285));
  AOI22_X1  g1085(.A1(new_n812), .A2(G159), .B1(G150), .B2(new_n817), .ZN(new_n1286));
  INV_X1    g1086(.A(G128), .ZN(new_n1287));
  OAI221_X1 g1087(.A(new_n280), .B1(new_n795), .B2(new_n202), .C1(new_n790), .C2(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1288), .B1(G137), .B2(new_n800), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1286), .A2(new_n1202), .A3(new_n1289), .ZN(new_n1290));
  OAI22_X1  g1090(.A1(new_n865), .A2(new_n876), .B1(new_n864), .B2(new_n1177), .ZN(new_n1291));
  OAI22_X1  g1091(.A1(new_n1281), .A2(new_n1285), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1275), .B1(new_n1292), .B2(new_n785), .ZN(new_n1293));
  AOI22_X1  g1093(.A1(new_n1158), .A2(new_n767), .B1(new_n1274), .B2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1160), .A2(new_n999), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1158), .B1(new_n1126), .B2(new_n1124), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1294), .B1(new_n1295), .B2(new_n1296), .ZN(G381));
  NOR4_X1   g1097(.A1(G393), .A2(G384), .A3(G381), .A4(G396), .ZN(new_n1298));
  AND2_X1   g1098(.A1(new_n1099), .A2(new_n1120), .ZN(new_n1299));
  AND2_X1   g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1046), .A2(new_n1050), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1023), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1053), .B1(new_n994), .B2(new_n995), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1058), .B1(new_n1303), .B2(new_n998), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1301), .B1(new_n1302), .B2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n730), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1306), .B1(new_n1193), .B2(new_n1160), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1194), .B1(new_n1159), .B2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1260), .A2(new_n767), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(new_n1243), .ZN(new_n1310));
  AND3_X1   g1110(.A1(new_n1263), .A2(KEYINPUT57), .A3(new_n1264), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1306), .B1(new_n1311), .B2(new_n1271), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1272), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1310), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1300), .A2(new_n1305), .A3(new_n1308), .A4(new_n1314), .ZN(G407));
  NAND3_X1  g1115(.A1(new_n1314), .A2(new_n702), .A3(new_n1308), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(G407), .A2(G213), .A3(new_n1316), .ZN(G409));
  NAND3_X1  g1117(.A1(new_n1260), .A2(new_n999), .A3(new_n1271), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1318), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1263), .A2(new_n767), .A3(new_n1264), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(new_n1243), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1308), .B1(new_n1319), .B2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1164), .A2(new_n1195), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT119), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1308), .A2(KEYINPUT119), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1322), .B1(new_n1327), .B2(G375), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1296), .B1(KEYINPUT60), .B2(new_n1160), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1270), .A2(new_n1266), .A3(KEYINPUT60), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1330), .A2(new_n730), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1294), .B1(new_n1329), .B2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(G384), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1332), .A2(new_n1333), .ZN(new_n1334));
  OAI211_X1 g1134(.A(G384), .B(new_n1294), .C1(new_n1329), .C2(new_n1331), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(G213), .ZN(new_n1338));
  NOR2_X1   g1138(.A1(new_n1338), .A2(G343), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1339), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1328), .A2(new_n1337), .A3(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1341), .A2(KEYINPUT62), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT61), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1339), .A2(G2897), .ZN(new_n1344));
  AND3_X1   g1144(.A1(new_n1334), .A2(new_n1335), .A3(new_n1344), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n1344), .B1(new_n1334), .B2(new_n1335), .ZN(new_n1346));
  NOR2_X1   g1146(.A1(new_n1345), .A2(new_n1346), .ZN(new_n1347));
  INV_X1    g1147(.A(new_n1321), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1323), .B1(new_n1348), .B2(new_n1318), .ZN(new_n1349));
  AOI21_X1  g1149(.A(new_n1349), .B1(new_n1314), .B2(G378), .ZN(new_n1350));
  OAI21_X1  g1150(.A(new_n1347), .B1(new_n1350), .B2(new_n1339), .ZN(new_n1351));
  INV_X1    g1151(.A(KEYINPUT62), .ZN(new_n1352));
  NAND4_X1  g1152(.A1(new_n1328), .A2(new_n1352), .A3(new_n1337), .A4(new_n1340), .ZN(new_n1353));
  NAND4_X1  g1153(.A1(new_n1342), .A2(new_n1343), .A3(new_n1351), .A4(new_n1353), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(G387), .A2(new_n1299), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1305), .A2(G390), .ZN(new_n1356));
  XNOR2_X1  g1156(.A(G393), .B(new_n839), .ZN(new_n1357));
  AND4_X1   g1157(.A1(KEYINPUT127), .A2(new_n1355), .A3(new_n1356), .A4(new_n1357), .ZN(new_n1358));
  INV_X1    g1158(.A(KEYINPUT127), .ZN(new_n1359));
  OAI21_X1  g1159(.A(new_n1359), .B1(new_n1305), .B2(G390), .ZN(new_n1360));
  AOI22_X1  g1160(.A1(new_n1360), .A2(new_n1357), .B1(new_n1355), .B2(new_n1356), .ZN(new_n1361));
  OR2_X1    g1161(.A1(new_n1358), .A2(new_n1361), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1354), .A2(new_n1362), .ZN(new_n1363));
  NOR2_X1   g1163(.A1(new_n1358), .A2(new_n1361), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1328), .A2(new_n1340), .ZN(new_n1365));
  AOI21_X1  g1165(.A(KEYINPUT61), .B1(new_n1365), .B2(new_n1347), .ZN(new_n1366));
  XOR2_X1   g1166(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n1367));
  NAND2_X1  g1167(.A1(new_n1341), .A2(new_n1367), .ZN(new_n1368));
  NAND4_X1  g1168(.A1(new_n1328), .A2(KEYINPUT63), .A3(new_n1337), .A4(new_n1340), .ZN(new_n1369));
  NAND4_X1  g1169(.A1(new_n1364), .A2(new_n1366), .A3(new_n1368), .A4(new_n1369), .ZN(new_n1370));
  NAND2_X1  g1170(.A1(new_n1363), .A2(new_n1370), .ZN(G405));
  NAND2_X1  g1171(.A1(new_n1314), .A2(G378), .ZN(new_n1372));
  NAND2_X1  g1172(.A1(G375), .A2(new_n1308), .ZN(new_n1373));
  AND3_X1   g1173(.A1(new_n1372), .A2(new_n1336), .A3(new_n1373), .ZN(new_n1374));
  AOI21_X1  g1174(.A(new_n1336), .B1(new_n1372), .B2(new_n1373), .ZN(new_n1375));
  NOR2_X1   g1175(.A1(new_n1374), .A2(new_n1375), .ZN(new_n1376));
  XNOR2_X1  g1176(.A(new_n1376), .B(new_n1364), .ZN(G402));
endmodule


