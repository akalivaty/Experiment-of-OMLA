//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 1 1 1 0 1 0 0 0 1 1 1 0 0 1 1 0 0 0 1 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 1 0 1 0 1 0 0 1 1 1 1 1 1 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:33 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1263, new_n1264, new_n1266, new_n1267,
    new_n1268, new_n1269, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  AND2_X1   g0012(.A1(KEYINPUT64), .A2(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(KEYINPUT64), .A2(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(G50), .B1(G58), .B2(G68), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n209), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n212), .B(new_n220), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XOR2_X1   g0029(.A(G238), .B(G244), .Z(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT65), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT66), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n234), .B(new_n238), .Z(G358));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G351));
  OAI21_X1  g0046(.A(KEYINPUT70), .B1(new_n207), .B2(G1), .ZN(new_n247));
  INV_X1    g0047(.A(KEYINPUT70), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n248), .A2(new_n206), .A3(G20), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n251), .A2(new_n202), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(new_n216), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  AOI22_X1  g0057(.A1(new_n252), .A2(new_n257), .B1(new_n202), .B2(new_n254), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  AOI22_X1  g0059(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n259), .ZN(new_n260));
  OR2_X1    g0060(.A1(KEYINPUT64), .A2(G20), .ZN(new_n261));
  NAND2_X1  g0061(.A1(KEYINPUT64), .A2(G20), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n261), .A2(G33), .A3(new_n262), .ZN(new_n263));
  XNOR2_X1  g0063(.A(KEYINPUT8), .B(G58), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n260), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(new_n256), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n258), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G33), .A2(G41), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT67), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n216), .ZN(new_n272));
  NAND3_X1  g0072(.A1(KEYINPUT67), .A2(G33), .A3(G41), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G41), .ZN(new_n275));
  INV_X1    g0075(.A(G45), .ZN(new_n276));
  AOI21_X1  g0076(.A(G1), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n274), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(KEYINPUT69), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT69), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n274), .A2(new_n278), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G226), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n274), .A2(G274), .A3(new_n277), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT68), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND4_X1  g0087(.A1(new_n274), .A2(KEYINPUT68), .A3(G274), .A4(new_n277), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G1698), .ZN(new_n290));
  OR2_X1    g0090(.A1(KEYINPUT3), .A2(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(KEYINPUT3), .A2(G33), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n290), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  AND2_X1   g0093(.A1(KEYINPUT3), .A2(G33), .ZN(new_n294));
  NOR2_X1   g0094(.A1(KEYINPUT3), .A2(G33), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AOI22_X1  g0096(.A1(new_n293), .A2(G223), .B1(new_n296), .B2(G77), .ZN(new_n297));
  AOI21_X1  g0097(.A(G1698), .B1(new_n291), .B2(new_n292), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G222), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n272), .A2(new_n269), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n284), .A2(new_n289), .A3(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G169), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n268), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n306), .B1(G179), .B2(new_n304), .ZN(new_n307));
  XNOR2_X1  g0107(.A(new_n307), .B(KEYINPUT71), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT75), .ZN(new_n309));
  OAI211_X1 g0109(.A(G232), .B(new_n290), .C1(new_n294), .C2(new_n295), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT72), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g0112(.A(KEYINPUT3), .B(G33), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n313), .A2(KEYINPUT72), .A3(G232), .A4(new_n290), .ZN(new_n314));
  INV_X1    g0114(.A(G107), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT73), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT73), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(G107), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(new_n296), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n313), .A2(G238), .A3(G1698), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n312), .A2(new_n314), .A3(new_n320), .A4(new_n321), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n322), .A2(new_n302), .B1(new_n287), .B2(new_n288), .ZN(new_n323));
  AND3_X1   g0123(.A1(new_n274), .A2(new_n281), .A3(new_n278), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n281), .B1(new_n274), .B2(new_n278), .ZN(new_n325));
  OAI21_X1  g0125(.A(G244), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(G169), .B1(new_n323), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G77), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n254), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n250), .A2(G77), .ZN(new_n330));
  AND2_X1   g0130(.A1(new_n255), .A2(new_n216), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n253), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n329), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  XOR2_X1   g0133(.A(KEYINPUT8), .B(G58), .Z(new_n334));
  NAND2_X1  g0134(.A1(new_n261), .A2(new_n262), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n334), .A2(new_n259), .B1(new_n335), .B2(G77), .ZN(new_n336));
  XOR2_X1   g0136(.A(KEYINPUT15), .B(G87), .Z(new_n337));
  NAND4_X1  g0137(.A1(new_n337), .A2(KEYINPUT74), .A3(G33), .A4(new_n215), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT74), .ZN(new_n339));
  XNOR2_X1  g0139(.A(KEYINPUT15), .B(G87), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n339), .B1(new_n263), .B2(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n336), .A2(new_n338), .A3(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n333), .B1(new_n342), .B2(new_n256), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n309), .B1(new_n327), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n322), .A2(new_n302), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n345), .A2(new_n289), .A3(new_n326), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n305), .ZN(new_n347));
  INV_X1    g0147(.A(new_n343), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n347), .A2(KEYINPUT75), .A3(new_n348), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n346), .A2(G179), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n344), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n346), .A2(G200), .ZN(new_n353));
  INV_X1    g0153(.A(G190), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n353), .B(new_n343), .C1(new_n354), .C2(new_n346), .ZN(new_n355));
  AND3_X1   g0155(.A1(new_n308), .A2(new_n352), .A3(new_n355), .ZN(new_n356));
  XNOR2_X1  g0156(.A(new_n267), .B(KEYINPUT9), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n357), .B1(new_n304), .B2(new_n354), .ZN(new_n358));
  INV_X1    g0158(.A(new_n304), .ZN(new_n359));
  INV_X1    g0159(.A(G200), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT76), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n362), .A2(new_n363), .A3(KEYINPUT10), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(KEYINPUT10), .ZN(new_n365));
  OR2_X1    g0165(.A1(new_n363), .A2(KEYINPUT10), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n365), .B(new_n366), .C1(new_n358), .C2(new_n361), .ZN(new_n367));
  AND2_X1   g0167(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT83), .ZN(new_n369));
  OR2_X1    g0169(.A1(G223), .A2(G1698), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n370), .B1(G226), .B2(new_n290), .ZN(new_n371));
  INV_X1    g0171(.A(G33), .ZN(new_n372));
  INV_X1    g0172(.A(G87), .ZN(new_n373));
  OAI22_X1  g0173(.A1(new_n371), .A2(new_n296), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n216), .B1(new_n270), .B2(new_n269), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n277), .B1(new_n375), .B2(new_n273), .ZN(new_n376));
  AOI22_X1  g0176(.A1(new_n374), .A2(new_n302), .B1(new_n376), .B2(G232), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n305), .B1(new_n289), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n289), .A2(new_n377), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n378), .B1(new_n380), .B2(G179), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n251), .A2(new_n264), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n382), .A2(new_n257), .B1(new_n254), .B2(new_n264), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  XNOR2_X1  g0184(.A(G58), .B(G68), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(G20), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n259), .A2(G159), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT7), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n215), .A2(new_n296), .A3(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(G68), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n291), .A2(new_n207), .A3(new_n292), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n391), .B1(new_n392), .B2(KEYINPUT7), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n388), .B1(new_n390), .B2(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n331), .B1(new_n394), .B2(KEYINPUT16), .ZN(new_n395));
  OAI21_X1  g0195(.A(KEYINPUT7), .B1(new_n335), .B2(new_n313), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n296), .A2(new_n389), .A3(new_n207), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n396), .A2(G68), .A3(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n388), .ZN(new_n399));
  AOI21_X1  g0199(.A(KEYINPUT16), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n384), .B1(new_n395), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g0202(.A(KEYINPUT18), .B1(new_n381), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n379), .A2(G169), .ZN(new_n404));
  INV_X1    g0204(.A(G179), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n404), .B1(new_n405), .B2(new_n379), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT18), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n393), .A2(new_n390), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n399), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT16), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n256), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n383), .B1(new_n411), .B2(new_n400), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n406), .A2(new_n407), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n369), .B1(new_n403), .B2(new_n413), .ZN(new_n414));
  NOR2_X1   g0214(.A1(KEYINPUT83), .A2(KEYINPUT18), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(new_n381), .B2(new_n402), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT17), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n379), .A2(G200), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n289), .A2(new_n377), .A3(G190), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n417), .B1(new_n412), .B2(new_n420), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n402), .A2(KEYINPUT17), .A3(new_n419), .A4(new_n418), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n416), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n414), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n356), .A2(new_n368), .A3(new_n424), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n253), .A2(G68), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT80), .ZN(new_n427));
  OAI21_X1  g0227(.A(KEYINPUT79), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT12), .ZN(new_n429));
  OR2_X1    g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n428), .B(new_n429), .C1(KEYINPUT79), .C2(new_n426), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n257), .A2(G68), .A3(new_n250), .ZN(new_n432));
  AND3_X1   g0232(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  AOI22_X1  g0233(.A1(new_n259), .A2(G50), .B1(G20), .B2(new_n391), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n434), .B1(new_n263), .B2(new_n328), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n256), .ZN(new_n436));
  XNOR2_X1  g0236(.A(new_n436), .B(KEYINPUT11), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n433), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n283), .A2(G238), .B1(new_n287), .B2(new_n288), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT13), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT78), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n442), .A2(G33), .A3(G97), .ZN(new_n443));
  INV_X1    g0243(.A(G97), .ZN(new_n444));
  OAI21_X1  g0244(.A(KEYINPUT78), .B1(new_n372), .B2(new_n444), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n298), .A2(G226), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(KEYINPUT77), .B1(new_n293), .B2(G232), .ZN(new_n447));
  OAI211_X1 g0247(.A(G232), .B(G1698), .C1(new_n294), .C2(new_n295), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT77), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n446), .B1(new_n447), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(new_n302), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n440), .A2(new_n441), .A3(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(G238), .B1(new_n324), .B2(new_n325), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(new_n289), .ZN(new_n455));
  XNOR2_X1  g0255(.A(new_n448), .B(new_n449), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n301), .B1(new_n456), .B2(new_n446), .ZN(new_n457));
  OAI21_X1  g0257(.A(KEYINPUT13), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n453), .A2(new_n458), .A3(G190), .ZN(new_n459));
  NOR3_X1   g0259(.A1(new_n455), .A2(new_n457), .A3(KEYINPUT13), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n441), .B1(new_n440), .B2(new_n452), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n439), .B(new_n459), .C1(new_n462), .C2(new_n360), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT14), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n464), .B(G169), .C1(new_n460), .C2(new_n461), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n453), .A2(new_n458), .A3(G179), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI211_X1 g0267(.A(KEYINPUT81), .B(KEYINPUT14), .C1(new_n462), .C2(new_n305), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT81), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n305), .B1(new_n453), .B2(new_n458), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n469), .B1(new_n470), .B2(new_n464), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n467), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n438), .A2(KEYINPUT82), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT82), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n433), .A2(new_n437), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n463), .B1(new_n472), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n425), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  OAI211_X1 g0279(.A(G250), .B(G1698), .C1(new_n294), .C2(new_n295), .ZN(new_n480));
  NAND2_X1  g0280(.A1(G33), .A2(G283), .ZN(new_n481));
  OAI211_X1 g0281(.A(G244), .B(new_n290), .C1(new_n294), .C2(new_n295), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT4), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n480), .B(new_n481), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(KEYINPUT4), .B1(new_n298), .B2(G244), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n302), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(KEYINPUT5), .A2(G41), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  NOR2_X1   g0288(.A1(KEYINPUT5), .A2(G41), .ZN(new_n489));
  OR2_X1    g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n276), .A2(G1), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n490), .A2(new_n274), .A3(G274), .A4(new_n491), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n491), .B1(new_n488), .B2(new_n489), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n274), .A2(new_n493), .A3(G257), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n486), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n305), .ZN(new_n496));
  AND3_X1   g0296(.A1(new_n396), .A2(new_n319), .A3(new_n397), .ZN(new_n497));
  AND3_X1   g0297(.A1(new_n259), .A2(KEYINPUT84), .A3(G77), .ZN(new_n498));
  AOI21_X1  g0298(.A(KEYINPUT84), .B1(new_n259), .B2(G77), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT6), .ZN(new_n501));
  NOR3_X1   g0301(.A1(new_n501), .A2(new_n444), .A3(G107), .ZN(new_n502));
  XNOR2_X1  g0302(.A(G97), .B(G107), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n502), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n500), .B1(new_n504), .B2(new_n215), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n256), .B1(new_n497), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n253), .A2(G97), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n257), .B1(G1), .B2(new_n372), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n508), .B1(new_n509), .B2(new_n444), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n506), .A2(new_n511), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n486), .A2(new_n405), .A3(new_n492), .A4(new_n494), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n496), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n495), .A2(G200), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n396), .A2(new_n319), .A3(new_n397), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n503), .A2(new_n501), .ZN(new_n517));
  INV_X1    g0317(.A(new_n502), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n335), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n516), .A2(new_n520), .A3(new_n500), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n510), .B1(new_n521), .B2(new_n256), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n486), .A2(G190), .A3(new_n492), .A4(new_n494), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n515), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n514), .A2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT85), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n313), .A2(G238), .A3(new_n290), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT86), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n298), .A2(KEYINPUT86), .A3(G238), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n293), .A2(G244), .ZN(new_n533));
  NAND2_X1  g0333(.A1(G33), .A2(G116), .ZN(new_n534));
  AND2_X1   g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n301), .B1(new_n532), .B2(new_n535), .ZN(new_n536));
  OR2_X1    g0336(.A1(new_n491), .A2(G250), .ZN(new_n537));
  OR3_X1    g0337(.A1(new_n276), .A2(G1), .A3(G274), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n537), .A2(new_n274), .A3(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  OAI21_X1  g0340(.A(G200), .B1(new_n536), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n445), .A2(new_n443), .A3(KEYINPUT19), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n215), .ZN(new_n543));
  XNOR2_X1  g0343(.A(KEYINPUT73), .B(G107), .ZN(new_n544));
  NOR2_X1   g0344(.A1(G87), .A2(G97), .ZN(new_n545));
  AND3_X1   g0345(.A1(new_n544), .A2(KEYINPUT87), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(KEYINPUT87), .B1(new_n544), .B2(new_n545), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n543), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n215), .A2(new_n313), .A3(G68), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT19), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n550), .B1(new_n263), .B2(new_n444), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n548), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n552), .A2(new_n256), .B1(new_n254), .B2(new_n340), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n533), .A2(new_n534), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n554), .B1(new_n530), .B2(new_n531), .ZN(new_n555));
  OAI211_X1 g0355(.A(G190), .B(new_n539), .C1(new_n555), .C2(new_n301), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n332), .B1(new_n206), .B2(G33), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(G87), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n541), .A2(new_n553), .A3(new_n556), .A4(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n544), .A2(new_n545), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT87), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n544), .A2(KEYINPUT87), .A3(new_n545), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n562), .A2(new_n563), .B1(new_n215), .B2(new_n542), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n551), .A2(new_n549), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n256), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n340), .A2(new_n254), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n557), .A2(new_n337), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n305), .B1(new_n536), .B2(new_n540), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n405), .B(new_n539), .C1(new_n555), .C2(new_n301), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  AND2_X1   g0372(.A1(new_n559), .A2(new_n572), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n298), .A2(G250), .B1(G33), .B2(G294), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n313), .A2(G257), .A3(G1698), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n301), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n274), .A2(new_n493), .A3(G264), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n492), .A2(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n405), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT91), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT23), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n315), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n581), .B1(new_n215), .B2(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n335), .A2(KEYINPUT91), .A3(new_n582), .A4(new_n315), .ZN(new_n585));
  OAI21_X1  g0385(.A(KEYINPUT23), .B1(new_n319), .B2(new_n207), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n207), .A2(G33), .A3(G116), .ZN(new_n587));
  AND4_X1   g0387(.A1(new_n584), .A2(new_n585), .A3(new_n586), .A4(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT24), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n373), .A2(KEYINPUT90), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n215), .A2(new_n313), .A3(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT22), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n215), .A2(new_n313), .A3(KEYINPUT22), .A4(new_n590), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n588), .A2(new_n589), .A3(new_n593), .A4(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n593), .A2(new_n594), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n585), .A2(new_n586), .A3(new_n584), .A4(new_n587), .ZN(new_n597));
  OAI21_X1  g0397(.A(KEYINPUT24), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n331), .B1(new_n595), .B2(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(KEYINPUT25), .B1(new_n254), .B2(new_n315), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n254), .A2(KEYINPUT25), .A3(new_n315), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n557), .A2(G107), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  OAI221_X1 g0404(.A(new_n580), .B1(G169), .B2(new_n579), .C1(new_n599), .C2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n595), .A2(new_n598), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n256), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n579), .A2(new_n354), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n360), .B1(new_n576), .B2(new_n578), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n607), .A2(new_n610), .A3(new_n603), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n527), .A2(new_n573), .A3(new_n605), .A4(new_n611), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n253), .A2(G116), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n613), .B1(new_n557), .B2(G116), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n256), .B1(new_n207), .B2(G116), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n372), .A2(G97), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n481), .ZN(new_n617));
  OAI21_X1  g0417(.A(KEYINPUT89), .B1(new_n335), .B2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT89), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n215), .A2(new_n619), .A3(new_n481), .A4(new_n616), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n615), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n621), .A2(KEYINPUT20), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT20), .ZN(new_n623));
  AOI211_X1 g0423(.A(new_n623), .B(new_n615), .C1(new_n618), .C2(new_n620), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n614), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n274), .A2(new_n493), .A3(G270), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n492), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n313), .A2(G264), .A3(G1698), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n313), .A2(G257), .A3(new_n290), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n296), .A2(G303), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT88), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n629), .A2(new_n630), .A3(KEYINPUT88), .A4(new_n631), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n302), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n628), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n625), .B1(G200), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n638), .B1(new_n354), .B2(new_n637), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n625), .A2(new_n637), .A3(KEYINPUT21), .A4(G169), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n635), .A2(new_n302), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n632), .A2(new_n633), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n627), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n643), .A2(new_n625), .A3(G179), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n625), .A2(new_n637), .A3(G169), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT21), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n514), .A2(new_n524), .A3(KEYINPUT85), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n639), .A2(new_n645), .A3(new_n648), .A4(new_n649), .ZN(new_n650));
  NOR3_X1   g0450(.A1(new_n479), .A2(new_n612), .A3(new_n650), .ZN(G372));
  NAND3_X1  g0451(.A1(new_n605), .A2(new_n645), .A3(new_n648), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n514), .A2(new_n524), .ZN(new_n653));
  AND2_X1   g0453(.A1(new_n611), .A2(new_n559), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT26), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n559), .A2(new_n572), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n656), .B1(new_n657), .B2(new_n514), .ZN(new_n658));
  INV_X1    g0458(.A(new_n514), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n659), .A2(new_n559), .A3(new_n572), .A4(KEYINPUT26), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n655), .A2(new_n572), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n478), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n308), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n403), .A2(new_n413), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n472), .ZN(new_n667));
  INV_X1    g0467(.A(new_n476), .ZN(new_n668));
  INV_X1    g0468(.A(new_n352), .ZN(new_n669));
  AOI22_X1  g0469(.A1(new_n667), .A2(new_n668), .B1(new_n463), .B2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n420), .ZN(new_n671));
  AOI21_X1  g0471(.A(KEYINPUT17), .B1(new_n671), .B2(new_n402), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n412), .A2(new_n420), .A3(new_n417), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n666), .B1(new_n670), .B2(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n664), .B1(new_n676), .B2(new_n368), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n663), .A2(new_n677), .ZN(G369));
  NAND2_X1  g0478(.A1(new_n645), .A2(new_n648), .ZN(new_n679));
  INV_X1    g0479(.A(G13), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(G1), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n215), .A2(new_n681), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(G213), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(G343), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n625), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n679), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n645), .A2(new_n648), .A3(new_n639), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n689), .B1(new_n690), .B2(new_n688), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n691), .A2(G330), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n605), .A2(new_n611), .ZN(new_n693));
  INV_X1    g0493(.A(new_n687), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n694), .B1(new_n607), .B2(new_n603), .ZN(new_n695));
  OAI22_X1  g0495(.A1(new_n693), .A2(new_n695), .B1(new_n605), .B2(new_n694), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n692), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n687), .B1(new_n645), .B2(new_n648), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n698), .A2(new_n605), .A3(new_n611), .ZN(new_n699));
  OR2_X1    g0499(.A1(new_n605), .A2(new_n687), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n697), .A2(new_n702), .ZN(G399));
  NOR2_X1   g0503(.A1(new_n546), .A2(new_n547), .ZN(new_n704));
  INV_X1    g0504(.A(G116), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n210), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(G41), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(new_n206), .ZN(new_n710));
  AOI22_X1  g0510(.A1(new_n707), .A2(new_n710), .B1(new_n219), .B2(new_n709), .ZN(new_n711));
  XOR2_X1   g0511(.A(new_n711), .B(KEYINPUT28), .Z(new_n712));
  INV_X1    g0512(.A(new_n572), .ZN(new_n713));
  AND3_X1   g0513(.A1(new_n653), .A2(new_n559), .A3(new_n611), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n713), .B1(new_n714), .B2(new_n652), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n687), .B1(new_n715), .B2(new_n661), .ZN(new_n716));
  OAI21_X1  g0516(.A(KEYINPUT93), .B1(new_n716), .B2(KEYINPUT29), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n662), .A2(new_n694), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT93), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT29), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n718), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n658), .A2(KEYINPUT94), .A3(new_n660), .ZN(new_n722));
  OR2_X1    g0522(.A1(new_n660), .A2(KEYINPUT94), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n715), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n724), .A2(KEYINPUT29), .A3(new_n694), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n717), .A2(new_n721), .A3(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(G330), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n536), .A2(new_n540), .ZN(new_n728));
  AND2_X1   g0528(.A1(new_n486), .A2(new_n494), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n728), .A2(new_n729), .A3(new_n579), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n643), .A2(G179), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT30), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n730), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n728), .A2(G179), .A3(new_n579), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n735), .A2(new_n495), .A3(new_n637), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n732), .B1(new_n730), .B2(new_n731), .ZN(new_n737));
  AND2_X1   g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n734), .B1(new_n738), .B2(KEYINPUT92), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n736), .A2(new_n737), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT92), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  OAI211_X1 g0542(.A(KEYINPUT31), .B(new_n687), .C1(new_n739), .C2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(KEYINPUT31), .B1(new_n612), .B2(new_n650), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT31), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n734), .A2(new_n745), .A3(new_n737), .A4(new_n736), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(new_n687), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n727), .B1(new_n743), .B2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  AND2_X1   g0550(.A1(new_n726), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n712), .B1(new_n751), .B2(G1), .ZN(G364));
  NOR2_X1   g0552(.A1(new_n335), .A2(new_n680), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G45), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n710), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n692), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n757), .B1(G330), .B2(new_n691), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n708), .A2(new_n296), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G355), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n760), .B1(G116), .B2(new_n210), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n708), .A2(new_n313), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n763), .B1(new_n276), .B2(new_n219), .ZN(new_n764));
  OR2_X1    g0564(.A1(new_n242), .A2(new_n276), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n761), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G13), .A2(G33), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(G20), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n216), .B1(G20), .B2(new_n305), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  XOR2_X1   g0571(.A(new_n771), .B(KEYINPUT95), .Z(new_n772));
  OAI21_X1  g0572(.A(new_n756), .B1(new_n766), .B2(new_n772), .ZN(new_n773));
  NOR4_X1   g0573(.A1(new_n215), .A2(G179), .A3(G190), .A4(new_n360), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(G283), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n296), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NOR4_X1   g0577(.A1(new_n207), .A2(new_n354), .A3(new_n360), .A4(G179), .ZN(new_n778));
  XOR2_X1   g0578(.A(new_n778), .B(KEYINPUT101), .Z(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(G303), .ZN(new_n781));
  INV_X1    g0581(.A(G311), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n215), .A2(new_n405), .ZN(new_n783));
  NOR2_X1   g0583(.A1(G190), .A2(G200), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n780), .A2(new_n781), .B1(new_n782), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n354), .A2(G200), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n335), .B1(new_n788), .B2(G179), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n777), .B(new_n786), .C1(G294), .C2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n783), .ZN(new_n791));
  NOR3_X1   g0591(.A1(new_n791), .A2(KEYINPUT96), .A3(new_n788), .ZN(new_n792));
  INV_X1    g0592(.A(KEYINPUT96), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n793), .B1(new_n783), .B2(new_n787), .ZN(new_n794));
  OR2_X1    g0594(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G322), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n335), .A2(new_n405), .A3(new_n784), .ZN(new_n797));
  OR2_X1    g0597(.A1(new_n797), .A2(KEYINPUT98), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(KEYINPUT98), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(G329), .ZN(new_n802));
  OR3_X1    g0602(.A1(new_n791), .A2(KEYINPUT97), .A3(new_n360), .ZN(new_n803));
  OAI21_X1  g0603(.A(KEYINPUT97), .B1(new_n791), .B2(new_n360), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n803), .A2(G190), .A3(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n803), .A2(new_n354), .A3(new_n804), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  XNOR2_X1  g0608(.A(KEYINPUT33), .B(G317), .ZN(new_n809));
  AOI22_X1  g0609(.A1(G326), .A2(new_n806), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n790), .A2(new_n796), .A3(new_n802), .A4(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n789), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(new_n444), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n813), .B1(new_n808), .B2(G68), .ZN(new_n814));
  XOR2_X1   g0614(.A(new_n814), .B(KEYINPUT100), .Z(new_n815));
  INV_X1    g0615(.A(G159), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n800), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g0617(.A(KEYINPUT99), .B(KEYINPUT32), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n817), .B(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n296), .B1(new_n778), .B2(G87), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n820), .B1(new_n785), .B2(new_n328), .C1(new_n775), .C2(new_n315), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n821), .B1(new_n795), .B2(G58), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n819), .B(new_n822), .C1(new_n202), .C2(new_n805), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n811), .B1(new_n815), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n773), .B1(new_n824), .B2(new_n770), .ZN(new_n825));
  INV_X1    g0625(.A(new_n769), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n825), .B1(new_n691), .B2(new_n826), .ZN(new_n827));
  AND2_X1   g0627(.A1(new_n758), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(G396));
  AND4_X1   g0629(.A1(KEYINPUT103), .A2(new_n344), .A3(new_n351), .A4(new_n349), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n343), .B1(new_n346), .B2(new_n305), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n350), .B1(new_n831), .B2(KEYINPUT75), .ZN(new_n832));
  AOI21_X1  g0632(.A(KEYINPUT103), .B1(new_n832), .B2(new_n344), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n348), .A2(new_n687), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n355), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(KEYINPUT104), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT103), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n352), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n832), .A2(KEYINPUT103), .A3(new_n344), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n839), .A2(KEYINPUT104), .A3(new_n840), .A4(new_n836), .ZN(new_n841));
  OR2_X1    g0641(.A1(new_n352), .A2(new_n835), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(KEYINPUT105), .B1(new_n837), .B2(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n839), .A2(new_n840), .A3(new_n836), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT104), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT105), .ZN(new_n848));
  NAND4_X1  g0648(.A1(new_n847), .A2(new_n848), .A3(new_n842), .A4(new_n841), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n844), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(new_n718), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n850), .A2(new_n716), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n756), .B1(new_n854), .B2(new_n750), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(new_n750), .B2(new_n854), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n770), .A2(new_n767), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n756), .B1(G77), .B2(new_n858), .ZN(new_n859));
  OAI22_X1  g0659(.A1(new_n780), .A2(new_n315), .B1(new_n705), .B2(new_n785), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n775), .A2(new_n373), .ZN(new_n861));
  NOR4_X1   g0661(.A1(new_n860), .A2(new_n313), .A3(new_n813), .A4(new_n861), .ZN(new_n862));
  AOI22_X1  g0662(.A1(G283), .A2(new_n808), .B1(new_n806), .B2(G303), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n795), .A2(G294), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n801), .A2(G311), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n862), .A2(new_n863), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n785), .ZN(new_n867));
  AOI22_X1  g0667(.A1(new_n795), .A2(G143), .B1(G159), .B2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(G137), .ZN(new_n869));
  INV_X1    g0669(.A(G150), .ZN(new_n870));
  OAI221_X1 g0670(.A(new_n868), .B1(new_n869), .B2(new_n805), .C1(new_n870), .C2(new_n807), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n871), .B(KEYINPUT102), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT34), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n775), .A2(new_n391), .ZN(new_n875));
  AOI211_X1 g0675(.A(new_n296), .B(new_n875), .C1(G58), .C2(new_n789), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n876), .B1(new_n202), .B2(new_n780), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n877), .B1(G132), .B2(new_n801), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n872), .A2(new_n873), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n866), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n859), .B1(new_n881), .B2(new_n770), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n882), .B1(new_n768), .B2(new_n850), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT106), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n883), .B(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n856), .A2(new_n885), .ZN(G384));
  OR2_X1    g0686(.A1(new_n519), .A2(KEYINPUT35), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n519), .A2(KEYINPUT35), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n887), .A2(G116), .A3(new_n217), .A4(new_n888), .ZN(new_n889));
  XOR2_X1   g0689(.A(new_n889), .B(KEYINPUT36), .Z(new_n890));
  INV_X1    g0690(.A(G58), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n219), .B(G77), .C1(new_n891), .C2(new_n391), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n202), .A2(G68), .ZN(new_n893));
  AOI211_X1 g0693(.A(new_n206), .B(G13), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n890), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n473), .A2(new_n475), .A3(new_n687), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n896), .B(KEYINPUT107), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n463), .B(new_n897), .C1(new_n472), .C2(new_n476), .ZN(new_n898));
  INV_X1    g0698(.A(new_n467), .ZN(new_n899));
  INV_X1    g0699(.A(new_n471), .ZN(new_n900));
  NOR3_X1   g0700(.A1(new_n470), .A2(new_n469), .A3(new_n464), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n899), .B(new_n463), .C1(new_n900), .C2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n896), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n898), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n834), .A2(new_n687), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n906), .B1(new_n853), .B2(new_n908), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n394), .A2(KEYINPUT16), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n383), .B1(new_n411), .B2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n685), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(new_n414), .B2(new_n423), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n671), .A2(new_n402), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n406), .A2(new_n412), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT37), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n412), .A2(new_n912), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n916), .A2(new_n917), .A3(new_n918), .A4(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n381), .A2(new_n685), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n921), .A2(new_n911), .B1(new_n671), .B2(new_n402), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n920), .B1(new_n922), .B2(new_n918), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT38), .B1(new_n915), .B2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n915), .A2(KEYINPUT38), .A3(new_n923), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n909), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n665), .A2(new_n685), .ZN(new_n929));
  AND3_X1   g0729(.A1(new_n915), .A2(KEYINPUT38), .A3(new_n923), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT39), .ZN(new_n931));
  NOR3_X1   g0731(.A1(new_n930), .A2(new_n924), .A3(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT108), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(new_n672), .B2(new_n673), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n421), .A2(new_n422), .A3(KEYINPUT108), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n935), .A2(new_n666), .A3(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n919), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n916), .A2(new_n917), .A3(new_n919), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(KEYINPUT37), .ZN(new_n940));
  AOI22_X1  g0740(.A1(new_n937), .A2(new_n938), .B1(new_n920), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n926), .B1(new_n941), .B2(KEYINPUT38), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n931), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n667), .A2(new_n668), .A3(new_n694), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n933), .A2(new_n943), .A3(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n928), .A2(new_n929), .A3(new_n946), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n478), .A2(new_n717), .A3(new_n725), .A4(new_n721), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n677), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n947), .B(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  OAI211_X1 g0751(.A(KEYINPUT31), .B(new_n687), .C1(new_n740), .C2(new_n733), .ZN(new_n952));
  AOI22_X1  g0752(.A1(new_n748), .A2(new_n952), .B1(new_n898), .B2(new_n904), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n850), .A2(new_n953), .A3(new_n942), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(KEYINPUT40), .ZN(new_n955));
  AOI21_X1  g0755(.A(KEYINPUT40), .B1(new_n925), .B2(new_n926), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n956), .A2(new_n850), .A3(new_n953), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n479), .B1(new_n748), .B2(new_n952), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n958), .A2(new_n959), .ZN(new_n962));
  NOR3_X1   g0762(.A1(new_n961), .A2(new_n962), .A3(new_n727), .ZN(new_n963));
  OAI22_X1  g0763(.A1(new_n951), .A2(new_n963), .B1(new_n206), .B2(new_n753), .ZN(new_n964));
  AND2_X1   g0764(.A1(new_n951), .A2(new_n963), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n895), .B1(new_n964), .B2(new_n965), .ZN(G367));
  OAI21_X1  g0766(.A(new_n653), .B1(new_n522), .B2(new_n694), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n514), .B1(new_n967), .B2(new_n605), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT111), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n968), .A2(new_n969), .ZN(new_n971));
  AND3_X1   g0771(.A1(new_n970), .A2(new_n694), .A3(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n694), .B1(new_n553), .B2(new_n558), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT109), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n713), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n657), .B2(new_n975), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT110), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(KEYINPUT43), .B1(new_n977), .B2(new_n978), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n659), .A2(new_n687), .ZN(new_n982));
  AND2_X1   g0782(.A1(new_n967), .A2(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n983), .A2(new_n699), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT112), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n984), .B(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(KEYINPUT42), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n986), .A2(KEYINPUT42), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n973), .B(new_n981), .C1(new_n988), .C2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n989), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n972), .B1(new_n991), .B2(new_n987), .ZN(new_n992));
  AND2_X1   g0792(.A1(new_n977), .A2(KEYINPUT43), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n981), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n990), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n697), .A2(new_n983), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n996), .B(new_n990), .C1(new_n992), .C2(new_n994), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n709), .B(KEYINPUT41), .Z(new_n1000));
  OAI21_X1  g0800(.A(new_n699), .B1(new_n696), .B2(new_n698), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n692), .B(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n751), .A2(KEYINPUT115), .A3(new_n1002), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n726), .A2(new_n1002), .A3(new_n750), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT115), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT44), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n967), .A2(new_n982), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1008), .B1(new_n702), .B2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n701), .A2(KEYINPUT44), .A3(new_n983), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT113), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n699), .A2(new_n700), .A3(new_n1009), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT45), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1014), .B(new_n1015), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1012), .A2(new_n1013), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(KEYINPUT114), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n697), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT114), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1013), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1012), .A2(new_n1016), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1020), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1007), .A2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1000), .B1(new_n1026), .B2(new_n751), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n754), .A2(G1), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n998), .B(new_n999), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n772), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n210), .B2(new_n340), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n238), .A2(new_n763), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n756), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n774), .A2(G97), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n778), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1035), .A2(new_n705), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1034), .B(new_n296), .C1(new_n1036), .C2(KEYINPUT46), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(G317), .B2(new_n801), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n779), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n867), .A2(G283), .B1(new_n319), .B2(new_n789), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(G303), .B2(new_n795), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(G294), .A2(new_n808), .B1(new_n806), .B2(G311), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n801), .A2(G137), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n789), .A2(G68), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n867), .A2(G50), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n313), .B1(new_n1035), .B2(new_n891), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(G77), .B2(new_n774), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .A4(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(G150), .B2(new_n795), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(G143), .A2(new_n806), .B1(new_n808), .B2(G159), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n1042), .A2(new_n1043), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT47), .Z(new_n1053));
  AOI21_X1  g0853(.A(new_n1033), .B1(new_n1053), .B2(new_n770), .ZN(new_n1054));
  OR2_X1    g0854(.A1(new_n977), .A2(new_n826), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1029), .A2(new_n1056), .ZN(G387));
  NAND2_X1  g0857(.A1(new_n1002), .A2(new_n1028), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n770), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n806), .A2(G322), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n795), .A2(G317), .B1(G303), .B2(new_n867), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1060), .B(new_n1061), .C1(new_n782), .C2(new_n807), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT48), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n789), .A2(G283), .B1(new_n778), .B2(G294), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT49), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n801), .A2(G326), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n313), .B1(new_n774), .B2(G116), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .A4(new_n1072), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(G159), .A2(new_n806), .B1(new_n808), .B2(new_n334), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n812), .A2(new_n340), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n296), .B1(new_n778), .B2(G77), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1034), .B(new_n1076), .C1(new_n391), .C2(new_n785), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n1075), .B(new_n1077), .C1(G150), .C2(new_n801), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n795), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1074), .B(new_n1078), .C1(new_n202), .C2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1059), .B1(new_n1073), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n763), .B1(new_n234), .B2(G45), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(new_n706), .B2(new_n759), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n264), .A2(G50), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT50), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n276), .B1(new_n391), .B2(new_n328), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n1086), .B(new_n706), .C1(new_n1085), .C2(new_n1084), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n1083), .A2(new_n1087), .B1(G107), .B2(new_n210), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n755), .B1(new_n1088), .B2(new_n1030), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n696), .B2(new_n826), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n751), .A2(new_n1002), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1004), .A2(new_n709), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n1058), .B1(new_n1081), .B2(new_n1090), .C1(new_n1091), .C2(new_n1092), .ZN(G393));
  INV_X1    g0893(.A(G294), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n785), .A2(new_n1094), .B1(new_n812), .B2(new_n705), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n296), .B1(new_n776), .B2(new_n1035), .C1(new_n775), .C2(new_n315), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(new_n801), .B2(G322), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT118), .Z(new_n1098));
  AOI211_X1 g0898(.A(new_n1095), .B(new_n1098), .C1(G303), .C2(new_n808), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n806), .A2(G317), .B1(G311), .B2(new_n795), .ZN(new_n1100));
  XOR2_X1   g0900(.A(new_n1100), .B(KEYINPUT52), .Z(new_n1101));
  INV_X1    g0901(.A(KEYINPUT117), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n1079), .A2(new_n816), .B1(new_n870), .B2(new_n805), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT51), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n867), .A2(new_n334), .B1(G77), .B2(new_n789), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1105), .B1(new_n807), .B2(new_n202), .ZN(new_n1106));
  XOR2_X1   g0906(.A(new_n1106), .B(KEYINPUT116), .Z(new_n1107));
  OAI21_X1  g0907(.A(new_n313), .B1(new_n1035), .B2(new_n391), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n1108), .B(new_n861), .C1(new_n801), .C2(G143), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1104), .A2(new_n1107), .A3(new_n1109), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n1099), .A2(new_n1101), .B1(new_n1102), .B2(new_n1110), .ZN(new_n1111));
  OR2_X1    g0911(.A1(new_n1110), .A2(new_n1102), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1059), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  AND2_X1   g0913(.A1(new_n762), .A2(new_n245), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1030), .B1(new_n444), .B2(new_n210), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n756), .B1(new_n1114), .B2(new_n1115), .C1(new_n1009), .C2(new_n826), .ZN(new_n1116));
  OR2_X1    g0916(.A1(new_n1113), .A2(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1023), .B(new_n1019), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1028), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1117), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  AOI211_X1 g0920(.A(G41), .B(new_n708), .C1(new_n1118), .C2(new_n1004), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1120), .B1(new_n1121), .B2(new_n1026), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(G390));
  AOI21_X1  g0923(.A(new_n932), .B1(new_n931), .B2(new_n942), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(new_n909), .B2(new_n945), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n850), .A2(new_n749), .A3(new_n905), .ZN(new_n1127));
  AND2_X1   g0927(.A1(new_n724), .A2(new_n694), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n907), .B1(new_n850), .B2(new_n1128), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n944), .B(new_n942), .C1(new_n1129), .C2(new_n906), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1126), .A2(new_n1127), .A3(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n727), .B1(new_n748), .B2(new_n952), .ZN(new_n1132));
  AND3_X1   g0932(.A1(new_n850), .A2(new_n905), .A3(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n942), .A2(new_n944), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n850), .A2(new_n1128), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n908), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1134), .B1(new_n1136), .B2(new_n905), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n718), .B1(new_n844), .B2(new_n849), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n905), .B1(new_n1138), .B2(new_n907), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1124), .B1(new_n1139), .B2(new_n944), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1133), .B1(new_n1137), .B2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1131), .A2(new_n1141), .A3(new_n1028), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(KEYINPUT119), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT119), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1131), .A2(new_n1141), .A3(new_n1144), .A4(new_n1028), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n478), .A2(new_n1132), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n948), .A2(new_n677), .A3(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n905), .B1(new_n850), .B2(new_n749), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n1133), .A2(new_n1149), .B1(new_n1138), .B2(new_n907), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n850), .A2(new_n1132), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1127), .B(new_n1129), .C1(new_n1151), .C2(new_n905), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1148), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1127), .ZN(new_n1155));
  NOR3_X1   g0955(.A1(new_n1137), .A2(new_n1140), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1133), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(new_n1126), .B2(new_n1130), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1154), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1131), .A2(new_n1141), .A3(new_n1153), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1159), .A2(new_n709), .A3(new_n1160), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n756), .B1(new_n334), .B2(new_n858), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n313), .B(new_n875), .C1(G77), .C2(new_n789), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n779), .A2(G87), .B1(G97), .B2(new_n867), .ZN(new_n1164));
  AND2_X1   g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n1165), .B1(new_n705), .B2(new_n1079), .C1(new_n1094), .C2(new_n800), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n776), .A2(new_n805), .B1(new_n807), .B2(new_n544), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(KEYINPUT54), .B(G143), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1168), .B(KEYINPUT120), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1170), .A2(new_n785), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n313), .B1(new_n812), .B2(new_n816), .C1(new_n775), .C2(new_n202), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT53), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n1035), .B2(new_n870), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n778), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n1171), .B(new_n1172), .C1(new_n1174), .C2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(G125), .ZN(new_n1177));
  INV_X1    g0977(.A(G132), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n1176), .B1(new_n1177), .B2(new_n800), .C1(new_n1178), .C2(new_n1079), .ZN(new_n1179));
  INV_X1    g0979(.A(G128), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n1180), .A2(new_n805), .B1(new_n807), .B2(new_n869), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n1166), .A2(new_n1167), .B1(new_n1179), .B2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1162), .B1(new_n1182), .B2(new_n770), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1183), .B1(new_n1124), .B2(new_n768), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1146), .A2(new_n1161), .A3(new_n1184), .ZN(G378));
  AOI22_X1  g0985(.A1(G97), .A2(new_n808), .B1(new_n806), .B2(G116), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n775), .A2(new_n891), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n867), .A2(new_n337), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n296), .A2(new_n275), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(G77), .B2(new_n778), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1188), .A2(new_n1045), .A3(new_n1189), .A4(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(G283), .B2(new_n801), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1186), .B(new_n1193), .C1(new_n315), .C2(new_n1079), .ZN(new_n1194));
  XOR2_X1   g0994(.A(new_n1194), .B(KEYINPUT121), .Z(new_n1195));
  AOI21_X1  g0995(.A(G50), .B1(new_n372), .B2(new_n275), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n1195), .A2(KEYINPUT58), .B1(new_n1190), .B2(new_n1196), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n1169), .A2(new_n778), .B1(G150), .B2(new_n789), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1198), .B1(new_n1079), .B2(new_n1180), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n807), .A2(new_n1178), .B1(new_n869), .B2(new_n785), .ZN(new_n1200));
  XOR2_X1   g1000(.A(new_n1200), .B(KEYINPUT122), .Z(new_n1201));
  AOI211_X1 g1001(.A(new_n1199), .B(new_n1201), .C1(G125), .C2(new_n806), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1203), .A2(KEYINPUT59), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n372), .B(new_n275), .C1(new_n775), .C2(new_n816), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(new_n801), .B2(G124), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT59), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1206), .B1(new_n1202), .B2(new_n1207), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1197), .B1(KEYINPUT58), .B2(new_n1195), .C1(new_n1204), .C2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(new_n770), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n364), .A2(new_n307), .A3(new_n367), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n268), .A2(new_n685), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1212), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n364), .A2(new_n307), .A3(new_n367), .A4(new_n1214), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n1213), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1216), .B1(new_n1213), .B2(new_n1215), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(new_n767), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n857), .A2(new_n202), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1210), .A2(new_n756), .A3(new_n1220), .A4(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1219), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(new_n958), .B2(G330), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n727), .B(new_n1219), .C1(new_n955), .C2(new_n957), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n947), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  AND2_X1   g1027(.A1(new_n850), .A2(new_n953), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n1228), .A2(new_n956), .B1(new_n954), .B2(KEYINPUT40), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1219), .B1(new_n1229), .B2(new_n727), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n946), .A2(new_n929), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(new_n927), .B2(new_n909), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n958), .A2(G330), .A3(new_n1224), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1230), .A2(new_n1232), .A3(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1227), .A2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1223), .B1(new_n1235), .B2(new_n1028), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1148), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1160), .A2(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1238), .A2(new_n1235), .A3(KEYINPUT57), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1239), .A2(new_n709), .ZN(new_n1240));
  AOI21_X1  g1040(.A(KEYINPUT57), .B1(new_n1238), .B2(new_n1235), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1236), .B1(new_n1240), .B2(new_n1241), .ZN(G375));
  INV_X1    g1042(.A(new_n1000), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1150), .A2(new_n1152), .A3(new_n1148), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1154), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1119), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n906), .A2(new_n767), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n756), .B1(G68), .B2(new_n858), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n780), .A2(new_n816), .B1(new_n870), .B2(new_n785), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1188), .B(new_n313), .C1(new_n202), .C2(new_n812), .ZN(new_n1250));
  AOI211_X1 g1050(.A(new_n1249), .B(new_n1250), .C1(G128), .C2(new_n801), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1251), .B1(new_n869), .B2(new_n1079), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n1178), .A2(new_n805), .B1(new_n807), .B2(new_n1170), .ZN(new_n1253));
  AOI211_X1 g1053(.A(new_n313), .B(new_n1075), .C1(G77), .C2(new_n774), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n779), .A2(G97), .B1(new_n319), .B2(new_n867), .ZN(new_n1255));
  AND2_X1   g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  OAI221_X1 g1056(.A(new_n1256), .B1(new_n776), .B2(new_n1079), .C1(new_n781), .C2(new_n800), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n705), .A2(new_n807), .B1(new_n805), .B2(new_n1094), .ZN(new_n1258));
  OAI22_X1  g1058(.A1(new_n1252), .A2(new_n1253), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1248), .B1(new_n1259), .B2(new_n770), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1246), .B1(new_n1247), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1245), .A2(new_n1261), .ZN(G381));
  NOR3_X1   g1062(.A1(G384), .A2(G393), .A3(G396), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1263), .A2(new_n1122), .A3(new_n1261), .A4(new_n1245), .ZN(new_n1264));
  OR4_X1    g1064(.A1(G387), .A2(G375), .A3(new_n1264), .A4(G378), .ZN(G407));
  AND3_X1   g1065(.A1(new_n1146), .A2(new_n1161), .A3(new_n1184), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n686), .A2(G213), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1266), .A2(new_n1268), .ZN(new_n1269));
  OAI211_X1 g1069(.A(G407), .B(G213), .C1(G375), .C2(new_n1269), .ZN(G409));
  INV_X1    g1070(.A(KEYINPUT60), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1244), .B1(new_n1153), .B2(new_n1271), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1150), .A2(new_n1152), .A3(new_n1148), .A4(KEYINPUT60), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1272), .A2(new_n709), .A3(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(G384), .B1(new_n1274), .B2(new_n1261), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1274), .A2(G384), .A3(new_n1261), .ZN(new_n1277));
  AOI22_X1  g1077(.A1(new_n1276), .A2(new_n1277), .B1(G2897), .B2(new_n1268), .ZN(new_n1278));
  AND3_X1   g1078(.A1(new_n1274), .A2(G384), .A3(new_n1261), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1268), .A2(G2897), .ZN(new_n1280));
  NOR3_X1   g1080(.A1(new_n1279), .A2(new_n1275), .A3(new_n1280), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1278), .A2(new_n1281), .ZN(new_n1282));
  OAI211_X1 g1082(.A(G378), .B(new_n1236), .C1(new_n1240), .C2(new_n1241), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1238), .A2(new_n1235), .A3(new_n1243), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1227), .A2(new_n1234), .A3(KEYINPUT123), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(new_n1028), .ZN(new_n1286));
  AOI21_X1  g1086(.A(KEYINPUT123), .B1(new_n1227), .B2(new_n1234), .ZN(new_n1287));
  OAI211_X1 g1087(.A(new_n1284), .B(new_n1222), .C1(new_n1286), .C2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(new_n1266), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1268), .B1(new_n1283), .B2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT124), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1282), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1283), .A2(new_n1289), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(new_n1267), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(KEYINPUT124), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1292), .A2(new_n1295), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1279), .A2(new_n1275), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1290), .A2(KEYINPUT63), .A3(new_n1297), .ZN(new_n1298));
  XNOR2_X1  g1098(.A(G393), .B(new_n828), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(G390), .B1(new_n1029), .B2(new_n1056), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n998), .A2(new_n999), .ZN(new_n1302));
  AOI22_X1  g1102(.A1(new_n1003), .A2(new_n1006), .B1(new_n1020), .B2(new_n1024), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n751), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1243), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1302), .B1(new_n1305), .B2(new_n1119), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1056), .ZN(new_n1307));
  NOR3_X1   g1107(.A1(new_n1306), .A2(new_n1307), .A3(new_n1122), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1300), .B1(new_n1301), .B2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT61), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1122), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1029), .A2(new_n1056), .A3(G390), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1311), .A2(new_n1312), .A3(new_n1299), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1309), .A2(new_n1310), .A3(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1293), .A2(new_n1267), .A3(new_n1297), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT63), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1314), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1296), .A2(new_n1298), .A3(new_n1317), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1315), .A2(KEYINPUT62), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1310), .B1(new_n1290), .B2(new_n1282), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT62), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1321), .B1(new_n1290), .B2(new_n1297), .ZN(new_n1322));
  NOR3_X1   g1122(.A1(new_n1319), .A2(new_n1320), .A3(new_n1322), .ZN(new_n1323));
  AND2_X1   g1123(.A1(new_n1309), .A2(new_n1313), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1318), .B1(new_n1323), .B2(new_n1324), .ZN(G405));
  NAND2_X1  g1125(.A1(G375), .A2(new_n1266), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT126), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1297), .A2(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT125), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1329), .A2(new_n1283), .A3(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1331), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1329), .B1(new_n1283), .B2(new_n1330), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1327), .B1(new_n1332), .B2(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1283), .A2(new_n1330), .ZN(new_n1335));
  NOR3_X1   g1135(.A1(new_n1279), .A2(new_n1275), .A3(KEYINPUT126), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1337), .A2(new_n1331), .A3(new_n1326), .ZN(new_n1338));
  AND3_X1   g1138(.A1(new_n1334), .A2(new_n1324), .A3(new_n1338), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1324), .B1(new_n1334), .B2(new_n1338), .ZN(new_n1340));
  NOR2_X1   g1140(.A1(new_n1339), .A2(new_n1340), .ZN(G402));
endmodule


