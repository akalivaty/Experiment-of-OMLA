//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 0 0 1 0 0 0 0 0 1 0 0 1 0 1 1 0 0 0 0 0 1 1 1 1 0 0 0 1 1 1 1 1 0 1 1 1 1 0 0 1 1 1 1 0 0 1 0 1 0 1 1 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:38 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1218, new_n1219,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI211_X1 g0005(.A(G50), .B(G77), .C1(new_n203), .C2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT0), .Z(new_n211));
  AOI22_X1  g0011(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n208), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT1), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  INV_X1    g0020(.A(G20), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n203), .A2(new_n205), .ZN(new_n223));
  INV_X1    g0023(.A(G50), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AOI211_X1 g0025(.A(new_n211), .B(new_n219), .C1(new_n222), .C2(new_n225), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(G232), .ZN(new_n228));
  XOR2_X1   g0028(.A(KEYINPUT2), .B(G226), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G270), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT65), .B(G264), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n230), .B(new_n234), .Z(G358));
  XOR2_X1   g0035(.A(G87), .B(G97), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT66), .ZN(new_n237));
  XOR2_X1   g0037(.A(G107), .B(G116), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G351));
  NAND3_X1  g0043(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(new_n220), .ZN(new_n245));
  XOR2_X1   g0045(.A(KEYINPUT8), .B(G58), .Z(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n221), .A2(G33), .ZN(new_n248));
  INV_X1    g0048(.A(G150), .ZN(new_n249));
  NOR2_X1   g0049(.A1(G20), .A2(G33), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  OAI22_X1  g0051(.A1(new_n247), .A2(new_n248), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n221), .B1(new_n223), .B2(new_n224), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n245), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G1), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(G13), .A3(G20), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT67), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND4_X1  g0058(.A1(new_n255), .A2(KEYINPUT67), .A3(G13), .A4(G20), .ZN(new_n259));
  AND2_X1   g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(new_n224), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n258), .A2(new_n259), .ZN(new_n262));
  INV_X1    g0062(.A(new_n245), .ZN(new_n263));
  OAI211_X1 g0063(.A(new_n262), .B(new_n263), .C1(G1), .C2(new_n221), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n254), .B(new_n261), .C1(new_n224), .C2(new_n264), .ZN(new_n265));
  XNOR2_X1  g0065(.A(new_n265), .B(KEYINPUT9), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT3), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G33), .ZN(new_n268));
  INV_X1    g0068(.A(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT3), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n271), .A2(G1698), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G222), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT3), .B(G33), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n274), .A2(G223), .A3(G1698), .ZN(new_n275));
  INV_X1    g0075(.A(G77), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n273), .B(new_n275), .C1(new_n276), .C2(new_n274), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n220), .B1(G33), .B2(G41), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n255), .B1(G41), .B2(G45), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G274), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G41), .ZN(new_n284));
  OAI211_X1 g0084(.A(G1), .B(G13), .C1(new_n269), .C2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(new_n280), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n283), .B1(new_n287), .B2(G226), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n279), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G200), .ZN(new_n290));
  INV_X1    g0090(.A(G190), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n266), .B(new_n290), .C1(new_n291), .C2(new_n289), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT10), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n293), .B1(new_n290), .B2(KEYINPUT70), .ZN(new_n294));
  AND2_X1   g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n292), .A2(new_n294), .ZN(new_n296));
  OR2_X1    g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n247), .A2(new_n262), .ZN(new_n298));
  INV_X1    g0098(.A(new_n264), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n298), .B1(new_n299), .B2(new_n247), .ZN(new_n300));
  OAI21_X1  g0100(.A(KEYINPUT75), .B1(new_n267), .B2(G33), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT75), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n302), .A2(new_n269), .A3(KEYINPUT3), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n301), .A2(new_n303), .A3(new_n268), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT76), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT7), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n306), .A2(G20), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n304), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n306), .B1(new_n274), .B2(G20), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n305), .B1(new_n304), .B2(new_n307), .ZN(new_n311));
  OAI21_X1  g0111(.A(G68), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n203), .B(new_n205), .C1(new_n201), .C2(new_n202), .ZN(new_n313));
  AOI22_X1  g0113(.A1(new_n313), .A2(G20), .B1(G159), .B2(new_n250), .ZN(new_n314));
  AOI21_X1  g0114(.A(KEYINPUT16), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n271), .A2(new_n307), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n309), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(G68), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n318), .A2(KEYINPUT16), .A3(new_n314), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(new_n245), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n300), .B1(new_n315), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n285), .A2(G232), .A3(new_n280), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n282), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n274), .A2(G226), .A3(G1698), .ZN(new_n324));
  INV_X1    g0124(.A(G1698), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n274), .A2(G223), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(G33), .A2(G87), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n324), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n323), .B1(new_n328), .B2(new_n278), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(G179), .ZN(new_n330));
  INV_X1    g0130(.A(G169), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n330), .B1(new_n331), .B2(new_n329), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n321), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT18), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(KEYINPUT18), .B1(new_n321), .B2(new_n332), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AOI211_X1 g0137(.A(new_n291), .B(new_n323), .C1(new_n328), .C2(new_n278), .ZN(new_n338));
  INV_X1    g0138(.A(G200), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n328), .A2(new_n278), .ZN(new_n340));
  INV_X1    g0140(.A(new_n323), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n339), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n338), .A2(new_n342), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n343), .B(new_n300), .C1(new_n315), .C2(new_n320), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT17), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n344), .B(new_n345), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n337), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n289), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n265), .B1(new_n348), .B2(G169), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT68), .ZN(new_n350));
  INV_X1    g0150(.A(G179), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n349), .A2(new_n350), .B1(new_n351), .B2(new_n348), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n352), .B1(new_n350), .B2(new_n349), .ZN(new_n353));
  AND2_X1   g0153(.A1(new_n287), .A2(G244), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n272), .A2(G232), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n274), .A2(G238), .A3(G1698), .ZN(new_n356));
  XNOR2_X1  g0156(.A(KEYINPUT69), .B(G107), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n355), .B(new_n356), .C1(new_n274), .C2(new_n357), .ZN(new_n358));
  AOI211_X1 g0158(.A(new_n283), .B(new_n354), .C1(new_n358), .C2(new_n278), .ZN(new_n359));
  AND2_X1   g0159(.A1(new_n359), .A2(new_n351), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n246), .A2(new_n250), .B1(G20), .B2(G77), .ZN(new_n361));
  XNOR2_X1  g0161(.A(KEYINPUT15), .B(G87), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n361), .B1(new_n248), .B2(new_n362), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n363), .A2(new_n245), .B1(new_n276), .B2(new_n260), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(new_n276), .B2(new_n264), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n365), .B1(new_n359), .B2(G169), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n360), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n365), .B1(new_n359), .B2(G190), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n369), .B1(new_n339), .B2(new_n359), .ZN(new_n370));
  AND2_X1   g0170(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n297), .A2(new_n347), .A3(new_n353), .A4(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n202), .A2(G20), .ZN(new_n373));
  OAI221_X1 g0173(.A(new_n373), .B1(new_n248), .B2(new_n276), .C1(new_n251), .C2(new_n224), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n245), .ZN(new_n375));
  XNOR2_X1  g0175(.A(new_n375), .B(KEYINPUT11), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n299), .A2(G68), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n262), .A2(G68), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT12), .ZN(new_n379));
  XNOR2_X1  g0179(.A(new_n378), .B(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n376), .A2(new_n377), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(KEYINPUT73), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT73), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n376), .A2(new_n380), .A3(new_n383), .A4(new_n377), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(G238), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n282), .B1(new_n286), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT72), .ZN(new_n389));
  XNOR2_X1  g0189(.A(new_n388), .B(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n274), .A2(G232), .A3(G1698), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n274), .A2(G226), .A3(new_n325), .ZN(new_n392));
  NAND2_X1  g0192(.A1(G33), .A2(G97), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(KEYINPUT71), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT71), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n391), .A2(new_n392), .A3(new_n396), .A4(new_n393), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n395), .A2(new_n397), .A3(new_n278), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n390), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(KEYINPUT13), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT13), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n390), .A2(new_n398), .A3(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n331), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT14), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n400), .A2(new_n402), .ZN(new_n405));
  OAI22_X1  g0205(.A1(new_n403), .A2(new_n404), .B1(new_n405), .B2(new_n351), .ZN(new_n406));
  AND3_X1   g0206(.A1(new_n390), .A2(new_n398), .A3(new_n401), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n401), .B1(new_n390), .B2(new_n398), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n404), .B(G169), .C1(new_n407), .C2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n386), .B1(new_n406), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(G200), .B1(new_n407), .B2(new_n408), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n400), .A2(G190), .A3(new_n402), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n385), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT74), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT74), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n385), .A2(new_n412), .A3(new_n413), .A4(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n411), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n372), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n255), .B(G45), .C1(new_n284), .C2(KEYINPUT5), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT5), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n423), .A2(G41), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(KEYINPUT78), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT78), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(new_n423), .B2(G41), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n422), .A2(new_n425), .A3(G274), .A4(new_n427), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n285), .B(G270), .C1(new_n421), .C2(new_n424), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n268), .A2(new_n270), .A3(G257), .A4(new_n325), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n268), .A2(new_n270), .A3(G264), .A4(G1698), .ZN(new_n433));
  INV_X1    g0233(.A(G303), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n432), .B(new_n433), .C1(new_n434), .C2(new_n274), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n278), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n431), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT79), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n255), .A2(G33), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n262), .A2(new_n263), .A3(G116), .A4(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(G116), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n258), .A2(new_n441), .A3(new_n259), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  AOI22_X1  g0243(.A1(new_n244), .A2(new_n220), .B1(G20), .B2(new_n441), .ZN(new_n444));
  NAND2_X1  g0244(.A1(G33), .A2(G283), .ZN(new_n445));
  INV_X1    g0245(.A(G97), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n445), .B(new_n221), .C1(G33), .C2(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n444), .A2(KEYINPUT20), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(KEYINPUT20), .B1(new_n444), .B2(new_n447), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n438), .B1(new_n443), .B2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n450), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n448), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n454), .A2(KEYINPUT79), .A3(new_n440), .A4(new_n442), .ZN(new_n455));
  AOI211_X1 g0255(.A(new_n351), .B(new_n437), .C1(new_n452), .C2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n437), .A2(G200), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n431), .A2(G190), .A3(new_n436), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n458), .A2(new_n452), .A3(new_n455), .A4(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n452), .A2(new_n455), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n331), .B1(new_n431), .B2(new_n436), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT80), .ZN(new_n464));
  AOI21_X1  g0264(.A(KEYINPUT21), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT21), .ZN(new_n466));
  AOI211_X1 g0266(.A(KEYINPUT80), .B(new_n466), .C1(new_n461), .C2(new_n462), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n457), .B(new_n460), .C1(new_n465), .C2(new_n467), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n268), .A2(new_n270), .A3(new_n221), .A4(G68), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n248), .A2(new_n446), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n469), .B1(KEYINPUT19), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(G87), .A2(G97), .ZN(new_n472));
  NAND3_X1  g0272(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n357), .A2(new_n472), .B1(new_n221), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n245), .B1(new_n471), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n260), .A2(new_n362), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n262), .A2(new_n263), .A3(G87), .A4(new_n439), .ZN(new_n477));
  AND3_X1   g0277(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n255), .A2(G45), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(G250), .ZN(new_n480));
  INV_X1    g0280(.A(G274), .ZN(new_n481));
  OAI22_X1  g0281(.A1(new_n278), .A2(new_n480), .B1(new_n481), .B2(new_n479), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n268), .A2(new_n270), .A3(G244), .A4(G1698), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n268), .A2(new_n270), .A3(G238), .A4(new_n325), .ZN(new_n484));
  NAND2_X1  g0284(.A1(G33), .A2(G116), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n482), .B1(new_n486), .B2(new_n278), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(G190), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n486), .A2(new_n278), .ZN(new_n489));
  INV_X1    g0289(.A(new_n482), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(G200), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n478), .A2(new_n488), .A3(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n262), .A2(new_n263), .A3(new_n439), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n475), .B(new_n476), .C1(new_n362), .C2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n491), .A2(new_n331), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n487), .A2(new_n351), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n268), .A2(new_n270), .A3(G250), .A4(new_n325), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n268), .A2(new_n270), .A3(G257), .A4(G1698), .ZN(new_n501));
  NAND2_X1  g0301(.A1(G33), .A2(G294), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n278), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n285), .B(G264), .C1(new_n421), .C2(new_n424), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n504), .A2(new_n428), .A3(new_n505), .ZN(new_n506));
  OR2_X1    g0306(.A1(new_n506), .A2(G190), .ZN(new_n507));
  INV_X1    g0307(.A(new_n428), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n504), .A2(new_n505), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT83), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n504), .A2(KEYINPUT83), .A3(new_n505), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n508), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n507), .B1(new_n513), .B2(G200), .ZN(new_n514));
  INV_X1    g0314(.A(G107), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n258), .A2(KEYINPUT25), .A3(new_n515), .A4(new_n259), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT81), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n262), .A2(G107), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n518), .B1(new_n519), .B2(KEYINPUT25), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n516), .A2(new_n517), .ZN(new_n521));
  OAI22_X1  g0321(.A1(new_n520), .A2(new_n521), .B1(new_n515), .B2(new_n494), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n485), .A2(G20), .ZN(new_n523));
  NOR3_X1   g0323(.A1(new_n221), .A2(KEYINPUT23), .A3(G107), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n357), .A2(G20), .ZN(new_n525));
  AOI211_X1 g0325(.A(new_n523), .B(new_n524), .C1(new_n525), .C2(KEYINPUT23), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n274), .A2(new_n221), .A3(G87), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(KEYINPUT22), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT22), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n274), .A2(new_n529), .A3(new_n221), .A4(G87), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(KEYINPUT24), .B1(new_n526), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n532), .A2(new_n263), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n526), .A2(new_n531), .A3(KEYINPUT24), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n522), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n499), .B1(new_n514), .B2(new_n535), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n285), .B(G257), .C1(new_n421), .C2(new_n424), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n428), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n274), .A2(G244), .A3(new_n325), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT4), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n274), .A2(KEYINPUT4), .A3(G244), .A4(new_n325), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n274), .A2(G250), .A3(G1698), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n541), .A2(new_n445), .A3(new_n542), .A4(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n538), .B1(new_n544), .B2(new_n278), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(G179), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n546), .B1(new_n331), .B2(new_n545), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n515), .A2(KEYINPUT6), .A3(G97), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n446), .A2(new_n515), .ZN(new_n549));
  NOR2_X1   g0349(.A1(G97), .A2(G107), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n548), .B1(new_n551), .B2(KEYINPUT6), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n552), .A2(G20), .B1(G77), .B2(new_n250), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n357), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n555), .B1(new_n310), .B2(new_n311), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n554), .B1(new_n556), .B2(KEYINPUT77), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT77), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n558), .B(new_n555), .C1(new_n310), .C2(new_n311), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n263), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n262), .A2(G97), .ZN(new_n561));
  INV_X1    g0361(.A(new_n494), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n561), .B1(new_n562), .B2(G97), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n547), .B1(new_n560), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n533), .A2(new_n534), .ZN(new_n566));
  INV_X1    g0366(.A(new_n522), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(new_n512), .ZN(new_n569));
  AOI21_X1  g0369(.A(KEYINPUT83), .B1(new_n504), .B2(new_n505), .ZN(new_n570));
  OAI211_X1 g0370(.A(G179), .B(new_n428), .C1(new_n569), .C2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n506), .A2(G169), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(KEYINPUT82), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT82), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n506), .A2(new_n574), .A3(G169), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n571), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n568), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n556), .A2(KEYINPUT77), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n578), .A2(new_n559), .A3(new_n553), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n245), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n545), .A2(new_n291), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n581), .B1(G200), .B2(new_n545), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n580), .A2(new_n563), .A3(new_n582), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n536), .A2(new_n565), .A3(new_n577), .A4(new_n583), .ZN(new_n584));
  NOR3_X1   g0384(.A1(new_n420), .A2(new_n468), .A3(new_n584), .ZN(G372));
  XNOR2_X1  g0385(.A(new_n333), .B(new_n334), .ZN(new_n586));
  INV_X1    g0386(.A(new_n411), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n587), .B1(new_n414), .B2(new_n367), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n586), .B1(new_n588), .B2(new_n346), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n297), .ZN(new_n590));
  AND2_X1   g0390(.A1(new_n590), .A2(new_n353), .ZN(new_n591));
  XNOR2_X1  g0391(.A(new_n498), .B(KEYINPUT84), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n536), .A2(new_n565), .A3(new_n583), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n435), .A2(new_n278), .ZN(new_n595));
  OAI21_X1  g0395(.A(G169), .B1(new_n595), .B2(new_n430), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n596), .B1(new_n452), .B2(new_n455), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n466), .B1(new_n597), .B2(KEYINPUT80), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n463), .A2(new_n464), .A3(KEYINPUT21), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n456), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n577), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n593), .B1(new_n594), .B2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT85), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n546), .B(new_n603), .C1(new_n331), .C2(new_n545), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n544), .A2(new_n278), .ZN(new_n605));
  INV_X1    g0405(.A(new_n538), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n331), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  AOI211_X1 g0407(.A(new_n351), .B(new_n538), .C1(new_n544), .C2(new_n278), .ZN(new_n608));
  OAI21_X1  g0408(.A(KEYINPUT85), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n604), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT26), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n580), .A2(new_n563), .ZN(new_n612));
  INV_X1    g0412(.A(new_n499), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n610), .A2(new_n611), .A3(new_n612), .A4(new_n613), .ZN(new_n614));
  OAI21_X1  g0414(.A(KEYINPUT26), .B1(new_n565), .B2(new_n499), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n602), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n419), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n591), .A2(new_n619), .ZN(G369));
  INV_X1    g0420(.A(G13), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n621), .A2(G20), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n255), .ZN(new_n623));
  OR2_X1    g0423(.A1(new_n623), .A2(KEYINPUT27), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(KEYINPUT27), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n624), .A2(G213), .A3(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(G343), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n461), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g0429(.A(new_n629), .B(KEYINPUT86), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n630), .B1(new_n468), .B2(KEYINPUT87), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n631), .B1(KEYINPUT87), .B2(new_n468), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n600), .A2(new_n630), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n632), .A2(G330), .A3(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n577), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n628), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n514), .A2(new_n535), .ZN(new_n638));
  INV_X1    g0438(.A(new_n628), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n577), .B(new_n638), .C1(new_n535), .C2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n635), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n600), .A2(new_n628), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n577), .A2(new_n638), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n645), .B1(new_n636), .B2(new_n639), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n642), .A2(new_n646), .ZN(G399));
  INV_X1    g0447(.A(KEYINPUT88), .ZN(new_n648));
  INV_X1    g0448(.A(new_n209), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n648), .B1(new_n649), .B2(G41), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n209), .A2(KEYINPUT88), .A3(new_n284), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  AND2_X1   g0453(.A1(new_n357), .A2(new_n472), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n441), .ZN(new_n655));
  NOR3_X1   g0455(.A1(new_n653), .A2(new_n255), .A3(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n656), .B1(new_n225), .B2(new_n653), .ZN(new_n657));
  XOR2_X1   g0457(.A(new_n657), .B(KEYINPUT28), .Z(new_n658));
  AOI21_X1  g0458(.A(new_n628), .B1(new_n602), .B2(new_n617), .ZN(new_n659));
  XNOR2_X1  g0459(.A(KEYINPUT90), .B(KEYINPUT29), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n598), .A2(new_n599), .ZN(new_n662));
  AND3_X1   g0462(.A1(new_n662), .A2(new_n457), .A3(new_n577), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n536), .A2(new_n565), .A3(new_n583), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n592), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n610), .A2(new_n612), .A3(new_n613), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(KEYINPUT26), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n612), .A2(new_n611), .A3(new_n547), .A4(new_n613), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OAI211_X1 g0469(.A(KEYINPUT29), .B(new_n639), .C1(new_n665), .C2(new_n669), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n670), .A2(KEYINPUT91), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(KEYINPUT91), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n661), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT30), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n511), .A2(new_n512), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n437), .A2(new_n491), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n674), .B1(new_n677), .B2(new_n546), .ZN(new_n678));
  INV_X1    g0478(.A(new_n545), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n679), .A2(new_n351), .A3(new_n437), .A4(new_n491), .ZN(new_n680));
  OAI22_X1  g0480(.A1(new_n678), .A2(KEYINPUT89), .B1(new_n513), .B2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n608), .A2(new_n675), .A3(new_n676), .A4(KEYINPUT30), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT89), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(new_n678), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n639), .B1(new_n682), .B2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n460), .ZN(new_n688));
  AOI211_X1 g0488(.A(new_n456), .B(new_n688), .C1(new_n598), .C2(new_n599), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n594), .A2(new_n689), .A3(new_n577), .A4(new_n639), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n687), .B1(new_n690), .B2(KEYINPUT31), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT31), .ZN(new_n692));
  INV_X1    g0492(.A(new_n678), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n680), .A2(new_n513), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AOI211_X1 g0495(.A(new_n692), .B(new_n639), .C1(new_n695), .C2(new_n683), .ZN(new_n696));
  OAI21_X1  g0496(.A(G330), .B1(new_n691), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n673), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT92), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n673), .A2(KEYINPUT92), .A3(new_n697), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n658), .B1(new_n702), .B2(G1), .ZN(G364));
  AOI21_X1  g0503(.A(new_n255), .B1(new_n622), .B2(G45), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n653), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n635), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(G330), .B1(new_n632), .B2(new_n633), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n632), .A2(new_n633), .ZN(new_n710));
  NOR2_X1   g0510(.A1(G13), .A2(G33), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(G20), .ZN(new_n713));
  XNOR2_X1  g0513(.A(new_n713), .B(KEYINPUT98), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n710), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n274), .A2(new_n209), .ZN(new_n716));
  INV_X1    g0516(.A(G355), .ZN(new_n717));
  OAI22_X1  g0517(.A1(new_n716), .A2(new_n717), .B1(G116), .B2(new_n209), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n649), .A2(new_n274), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(G45), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n720), .B1(new_n225), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n242), .A2(G45), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n718), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n220), .B1(G20), .B2(new_n331), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n713), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n706), .B1(new_n724), .B2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(G179), .A2(G200), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n729), .A2(G20), .A3(new_n291), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(G159), .ZN(new_n732));
  XNOR2_X1  g0532(.A(new_n732), .B(KEYINPUT94), .ZN(new_n733));
  XNOR2_X1  g0533(.A(new_n733), .B(KEYINPUT32), .ZN(new_n734));
  NAND2_X1  g0534(.A1(G20), .A2(G179), .ZN(new_n735));
  XOR2_X1   g0535(.A(new_n735), .B(KEYINPUT93), .Z(new_n736));
  NOR2_X1   g0536(.A1(new_n291), .A2(new_n339), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n221), .A2(G179), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n271), .B1(new_n742), .B2(G87), .ZN(new_n743));
  AOI22_X1  g0543(.A1(new_n739), .A2(G50), .B1(KEYINPUT95), .B2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n291), .A2(G200), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n736), .A2(new_n745), .ZN(new_n746));
  OAI211_X1 g0546(.A(new_n734), .B(new_n744), .C1(new_n201), .C2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n743), .A2(KEYINPUT95), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n221), .B1(new_n729), .B2(G190), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(new_n446), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n740), .A2(new_n291), .A3(G200), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(new_n515), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n748), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n736), .A2(new_n291), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n339), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n754), .A2(G200), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  OAI221_X1 g0558(.A(new_n753), .B1(new_n202), .B2(new_n756), .C1(new_n276), .C2(new_n758), .ZN(new_n759));
  AND2_X1   g0559(.A1(new_n731), .A2(KEYINPUT97), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n731), .A2(KEYINPUT97), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI22_X1  g0563(.A1(new_n763), .A2(G329), .B1(G326), .B2(new_n739), .ZN(new_n764));
  INV_X1    g0564(.A(G322), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n764), .B1(new_n765), .B2(new_n746), .ZN(new_n766));
  INV_X1    g0566(.A(G294), .ZN(new_n767));
  INV_X1    g0567(.A(G283), .ZN(new_n768));
  OAI221_X1 g0568(.A(new_n271), .B1(new_n749), .B2(new_n767), .C1(new_n751), .C2(new_n768), .ZN(new_n769));
  AND2_X1   g0569(.A1(new_n741), .A2(KEYINPUT96), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n741), .A2(KEYINPUT96), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n769), .B1(new_n773), .B2(G303), .ZN(new_n774));
  INV_X1    g0574(.A(G311), .ZN(new_n775));
  XOR2_X1   g0575(.A(KEYINPUT33), .B(G317), .Z(new_n776));
  OAI221_X1 g0576(.A(new_n774), .B1(new_n775), .B2(new_n758), .C1(new_n756), .C2(new_n776), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n747), .A2(new_n759), .B1(new_n766), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n728), .B1(new_n778), .B2(new_n725), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n707), .A2(new_n709), .B1(new_n715), .B2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(G396));
  OAI21_X1  g0581(.A(new_n274), .B1(new_n751), .B2(new_n202), .ZN(new_n782));
  INV_X1    g0582(.A(new_n749), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n782), .B1(G58), .B2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(G132), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n784), .B1(new_n762), .B2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n746), .ZN(new_n787));
  AOI22_X1  g0587(.A1(G137), .A2(new_n739), .B1(new_n787), .B2(G143), .ZN(new_n788));
  INV_X1    g0588(.A(G159), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n788), .B1(new_n756), .B2(new_n249), .C1(new_n789), .C2(new_n758), .ZN(new_n790));
  XOR2_X1   g0590(.A(new_n790), .B(KEYINPUT34), .Z(new_n791));
  AOI211_X1 g0591(.A(new_n786), .B(new_n791), .C1(G50), .C2(new_n773), .ZN(new_n792));
  INV_X1    g0592(.A(new_n751), .ZN(new_n793));
  AOI211_X1 g0593(.A(new_n274), .B(new_n750), .C1(G87), .C2(new_n793), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n794), .B1(new_n775), .B2(new_n762), .C1(new_n756), .C2(new_n768), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n773), .A2(G107), .B1(G303), .B2(new_n739), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(new_n767), .B2(new_n746), .ZN(new_n797));
  AOI211_X1 g0597(.A(new_n795), .B(new_n797), .C1(G116), .C2(new_n757), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n725), .B1(new_n792), .B2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n725), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(new_n712), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n799), .B1(G77), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n368), .A2(new_n628), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n365), .A2(new_n628), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n370), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n803), .B1(new_n368), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(new_n712), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n706), .B1(new_n802), .B2(new_n807), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n639), .B(new_n806), .C1(new_n665), .C2(new_n616), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n806), .B(KEYINPUT99), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n809), .B1(new_n810), .B2(new_n659), .ZN(new_n811));
  INV_X1    g0611(.A(new_n697), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n811), .A2(new_n812), .B1(new_n653), .B2(new_n705), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n811), .A2(new_n812), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n808), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  XOR2_X1   g0615(.A(new_n815), .B(KEYINPUT100), .Z(G384));
  NOR2_X1   g0616(.A1(new_n622), .A2(new_n255), .ZN(new_n817));
  INV_X1    g0617(.A(G330), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT102), .ZN(new_n819));
  INV_X1    g0619(.A(new_n686), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n628), .B1(new_n820), .B2(new_n681), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(new_n692), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n819), .B1(new_n691), .B2(new_n822), .ZN(new_n823));
  NOR3_X1   g0623(.A1(new_n584), .A2(new_n468), .A3(new_n628), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n821), .B1(new_n824), .B2(new_n692), .ZN(new_n825));
  INV_X1    g0625(.A(new_n822), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n825), .A2(KEYINPUT102), .A3(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n818), .B1(new_n823), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n419), .ZN(new_n829));
  AOI21_X1  g0629(.A(KEYINPUT16), .B1(new_n318), .B2(new_n314), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n300), .B1(new_n320), .B2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n626), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n831), .B1(new_n332), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(new_n344), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n834), .A2(KEYINPUT37), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT101), .ZN(new_n836));
  AND3_X1   g0636(.A1(new_n321), .A2(new_n836), .A3(new_n832), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n836), .B1(new_n321), .B2(new_n832), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n333), .B(new_n344), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n835), .B1(new_n839), .B2(KEYINPUT37), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n831), .A2(new_n832), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(new_n337), .B2(new_n346), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n840), .A2(new_n842), .A3(KEYINPUT38), .ZN(new_n843));
  OR2_X1    g0643(.A1(new_n837), .A2(new_n838), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT37), .ZN(new_n845));
  AND2_X1   g0645(.A1(new_n333), .A2(new_n344), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n839), .A2(KEYINPUT37), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n344), .B(KEYINPUT17), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n586), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n844), .ZN(new_n851));
  AOI22_X1  g0651(.A1(new_n847), .A2(new_n848), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n843), .B1(new_n852), .B2(KEYINPUT38), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n385), .A2(new_n639), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  AND2_X1   g0655(.A1(new_n855), .A2(new_n414), .ZN(new_n856));
  AOI22_X1  g0656(.A1(new_n418), .A2(new_n854), .B1(new_n411), .B2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n806), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NOR3_X1   g0659(.A1(new_n691), .A2(new_n819), .A3(new_n822), .ZN(new_n860));
  AOI21_X1  g0660(.A(KEYINPUT102), .B1(new_n825), .B2(new_n826), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n853), .B(new_n859), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n415), .A2(new_n417), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n855), .B1(new_n863), .B2(new_n411), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n856), .A2(new_n411), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n806), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n866), .B1(new_n823), .B2(new_n827), .ZN(new_n867));
  AND3_X1   g0667(.A1(new_n840), .A2(new_n842), .A3(KEYINPUT38), .ZN(new_n868));
  AOI21_X1  g0668(.A(KEYINPUT38), .B1(new_n840), .B2(new_n842), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n870), .A2(KEYINPUT40), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n862), .A2(KEYINPUT40), .B1(new_n867), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n829), .B1(new_n872), .B2(new_n818), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n419), .B1(new_n860), .B2(new_n861), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n873), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n591), .B1(new_n673), .B2(new_n420), .ZN(new_n876));
  XOR2_X1   g0676(.A(new_n875), .B(new_n876), .Z(new_n877));
  OAI21_X1  g0677(.A(KEYINPUT39), .B1(new_n868), .B2(new_n869), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT39), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n879), .B(new_n843), .C1(new_n852), .C2(KEYINPUT38), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n411), .A2(new_n628), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n803), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n857), .B1(new_n809), .B2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  OAI22_X1  g0687(.A1(new_n887), .A2(new_n870), .B1(new_n586), .B2(new_n832), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n817), .B1(new_n877), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n890), .B1(new_n889), .B2(new_n877), .ZN(new_n891));
  OAI211_X1 g0691(.A(G116), .B(new_n222), .C1(new_n552), .C2(KEYINPUT35), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n892), .B1(KEYINPUT35), .B2(new_n552), .ZN(new_n893));
  XOR2_X1   g0693(.A(new_n893), .B(KEYINPUT36), .Z(new_n894));
  OAI211_X1 g0694(.A(new_n225), .B(G77), .C1(new_n201), .C2(new_n202), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n895), .B1(G50), .B2(new_n202), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n896), .A2(G1), .A3(new_n621), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n891), .A2(new_n894), .A3(new_n897), .ZN(G367));
  OAI221_X1 g0698(.A(new_n726), .B1(new_n209), .B2(new_n362), .C1(new_n234), .C2(new_n720), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n706), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n751), .A2(new_n446), .ZN(new_n901));
  AOI211_X1 g0701(.A(new_n274), .B(new_n901), .C1(G317), .C2(new_n731), .ZN(new_n902));
  AOI21_X1  g0702(.A(KEYINPUT46), .B1(new_n742), .B2(G116), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n903), .B1(new_n555), .B2(new_n783), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  OAI221_X1 g0705(.A(new_n905), .B1(new_n768), .B2(new_n758), .C1(new_n767), .C2(new_n756), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n773), .A2(KEYINPUT46), .A3(G116), .ZN(new_n907));
  OAI22_X1  g0707(.A1(new_n434), .A2(new_n746), .B1(new_n738), .B2(new_n775), .ZN(new_n908));
  NOR3_X1   g0708(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  XOR2_X1   g0709(.A(new_n909), .B(KEYINPUT109), .Z(new_n910));
  AOI22_X1  g0710(.A1(new_n742), .A2(G58), .B1(new_n731), .B2(G137), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n911), .B(new_n274), .C1(new_n276), .C2(new_n751), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n758), .A2(new_n224), .ZN(new_n913));
  AOI211_X1 g0713(.A(new_n912), .B(new_n913), .C1(G143), .C2(new_n739), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(new_n789), .B2(new_n756), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n783), .A2(G68), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n746), .B2(new_n249), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n917), .B(KEYINPUT110), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n910), .B1(new_n915), .B2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT47), .ZN(new_n920));
  OR2_X1    g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n800), .B1(new_n919), .B2(new_n920), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n900), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT103), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n478), .A2(new_n639), .ZN(new_n925));
  OR2_X1    g0725(.A1(new_n592), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n613), .A2(new_n925), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n924), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n928), .B1(new_n924), .B2(new_n927), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(KEYINPUT104), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n714), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n923), .A2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT44), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n612), .A2(new_n628), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n934), .A2(new_n565), .A3(new_n583), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n610), .A2(new_n612), .A3(new_n628), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OR3_X1    g0737(.A1(new_n646), .A2(new_n933), .A3(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n933), .B1(new_n646), .B2(new_n937), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n646), .A2(new_n937), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT45), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n646), .A2(KEYINPUT45), .A3(new_n937), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AND3_X1   g0745(.A1(new_n940), .A2(new_n642), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n642), .B1(new_n940), .B2(new_n945), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OR3_X1    g0748(.A1(new_n641), .A2(KEYINPUT106), .A3(new_n643), .ZN(new_n949));
  OAI21_X1  g0749(.A(KEYINPUT106), .B1(new_n641), .B2(new_n643), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n645), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OR3_X1    g0751(.A1(new_n951), .A2(new_n634), .A3(KEYINPUT107), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n634), .A2(KEYINPUT107), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n634), .A2(KEYINPUT107), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n953), .A2(new_n954), .A3(new_n951), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n957), .B1(new_n700), .B2(new_n701), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n948), .B1(new_n958), .B2(KEYINPUT108), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT108), .ZN(new_n960));
  AOI211_X1 g0760(.A(new_n960), .B(new_n957), .C1(new_n700), .C2(new_n701), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n702), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n652), .B(KEYINPUT41), .Z(new_n963));
  AOI21_X1  g0763(.A(new_n705), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n645), .A2(new_n937), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(KEYINPUT42), .Z(new_n966));
  AOI22_X1  g0766(.A1(new_n937), .A2(new_n636), .B1(new_n547), .B2(new_n612), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n966), .B1(new_n628), .B2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT43), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n930), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n930), .A2(new_n969), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n971), .B(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n937), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n642), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT105), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n973), .A2(KEYINPUT105), .A3(new_n975), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n973), .A2(new_n975), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n932), .B1(new_n964), .B2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT111), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n982), .B(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(G387));
  NAND2_X1  g0785(.A1(new_n702), .A2(new_n956), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n700), .A2(new_n957), .A3(new_n701), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n986), .A2(new_n653), .A3(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n640), .A2(new_n637), .A3(new_n714), .ZN(new_n989));
  INV_X1    g0789(.A(new_n655), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n990), .A2(new_n716), .B1(G107), .B2(new_n209), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT112), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n990), .B(new_n721), .C1(new_n202), .C2(new_n276), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n246), .A2(new_n224), .ZN(new_n994));
  XOR2_X1   g0794(.A(KEYINPUT114), .B(KEYINPUT50), .Z(new_n995));
  XNOR2_X1  g0795(.A(new_n994), .B(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n719), .B1(new_n993), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n230), .A2(G45), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n997), .B1(new_n998), .B2(KEYINPUT113), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n998), .A2(KEYINPUT113), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n992), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n706), .B1(new_n1001), .B2(new_n727), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n901), .A2(new_n271), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n742), .A2(G77), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n1003), .B(new_n1004), .C1(new_n249), .C2(new_n730), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n224), .A2(new_n746), .B1(new_n738), .B2(new_n789), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n749), .A2(new_n362), .ZN(new_n1007));
  NOR3_X1   g0807(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n1008), .B1(new_n202), .B2(new_n758), .C1(new_n247), .C2(new_n756), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n274), .B1(new_n731), .B2(G326), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(G317), .A2(new_n787), .B1(new_n739), .B2(G322), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1011), .B1(new_n756), .B2(new_n775), .C1(new_n434), .C2(new_n758), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT48), .Z(new_n1013));
  OAI22_X1  g0813(.A1(new_n741), .A2(new_n767), .B1(new_n749), .B2(new_n768), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n1010), .B1(new_n441), .B2(new_n751), .C1(new_n1015), .C2(KEYINPUT49), .ZN(new_n1016));
  AND2_X1   g0816(.A1(new_n1015), .A2(KEYINPUT49), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1009), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1002), .B1(new_n1018), .B2(new_n725), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n956), .A2(new_n705), .B1(new_n989), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n988), .A2(new_n1020), .ZN(G393));
  NAND2_X1  g0821(.A1(new_n948), .A2(new_n705), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n974), .A2(new_n713), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n239), .A2(new_n720), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n726), .B1(new_n446), .B2(new_n209), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n706), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT115), .Z(new_n1027));
  AOI22_X1  g0827(.A1(G311), .A2(new_n787), .B1(new_n739), .B2(G317), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n1028), .B(KEYINPUT52), .Z(new_n1029));
  NOR2_X1   g0829(.A1(new_n749), .A2(new_n441), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n752), .A2(new_n274), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n1031), .B1(new_n768), .B2(new_n741), .C1(new_n765), .C2(new_n730), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n1030), .B(new_n1032), .C1(G294), .C2(new_n757), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1029), .B(new_n1033), .C1(new_n434), .C2(new_n756), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n1034), .A2(KEYINPUT116), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(KEYINPUT116), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n749), .A2(new_n276), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n742), .A2(G68), .B1(new_n731), .B2(G143), .ZN(new_n1038));
  INV_X1    g0838(.A(G87), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1038), .B(new_n274), .C1(new_n1039), .C2(new_n751), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n1037), .B(new_n1040), .C1(new_n246), .C2(new_n757), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n249), .A2(new_n738), .B1(new_n746), .B2(new_n789), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT51), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1041), .B(new_n1043), .C1(new_n224), .C2(new_n756), .ZN(new_n1044));
  AND3_X1   g0844(.A1(new_n1035), .A2(new_n1036), .A3(new_n1044), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1023), .B(new_n1027), .C1(new_n1045), .C2(new_n800), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1022), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT117), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n946), .A2(new_n947), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n986), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(KEYINPUT117), .B1(new_n958), .B2(new_n948), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n653), .B1(new_n959), .B2(new_n961), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1048), .B1(new_n1054), .B2(new_n1055), .ZN(G390));
  NAND2_X1  g0856(.A1(new_n867), .A2(G330), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n857), .B1(new_n697), .B2(new_n858), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n803), .B1(new_n659), .B2(new_n806), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n857), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n810), .ZN(new_n1064));
  OAI21_X1  g0864(.A(G330), .B1(new_n860), .B2(new_n861), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1064), .B1(new_n1065), .B2(KEYINPUT119), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT119), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n828), .A2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1063), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n812), .A2(new_n806), .A3(new_n1063), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n805), .A2(new_n368), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n639), .B(new_n1071), .C1(new_n665), .C2(new_n669), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n885), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1070), .A2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1062), .B1(new_n1069), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1057), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n878), .B(new_n880), .C1(new_n886), .C2(new_n882), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n847), .A2(new_n848), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n850), .A2(new_n851), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT38), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n882), .B1(new_n1083), .B2(new_n843), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1073), .A2(new_n1063), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1078), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1077), .A2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n883), .B1(new_n1060), .B2(new_n857), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n881), .A2(new_n1089), .B1(new_n1085), .B2(new_n1084), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n1088), .A2(KEYINPUT118), .B1(new_n1090), .B2(new_n1070), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT118), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1077), .A2(new_n1087), .A3(new_n1092), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n829), .B(new_n591), .C1(new_n420), .C2(new_n673), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n1076), .A2(new_n1091), .A3(new_n1093), .A4(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(KEYINPUT118), .B1(new_n1090), .B2(new_n1057), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1090), .A2(new_n1070), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1097), .A2(new_n1093), .A3(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1060), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n810), .B1(new_n828), .B2(new_n1067), .ZN(new_n1101));
  AOI211_X1 g0901(.A(KEYINPUT119), .B(new_n818), .C1(new_n823), .C2(new_n827), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n857), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1075), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1100), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1099), .B1(new_n1105), .B2(new_n1094), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1096), .A2(new_n1106), .A3(new_n653), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT120), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1099), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n881), .A2(new_n711), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n706), .B1(new_n246), .B2(new_n801), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n271), .B1(new_n751), .B2(new_n202), .ZN(new_n1112));
  AOI211_X1 g0912(.A(new_n1037), .B(new_n1112), .C1(new_n763), .C2(G294), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n1113), .B1(new_n446), .B2(new_n758), .C1(new_n357), .C2(new_n756), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n773), .A2(G87), .B1(G116), .B2(new_n787), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(new_n768), .B2(new_n738), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n274), .B1(new_n749), .B2(new_n789), .C1(new_n751), .C2(new_n224), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(G128), .B2(new_n739), .ZN(new_n1118));
  INV_X1    g0918(.A(G137), .ZN(new_n1119));
  XOR2_X1   g0919(.A(KEYINPUT54), .B(G143), .Z(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  OAI221_X1 g0921(.A(new_n1118), .B1(new_n756), .B2(new_n1119), .C1(new_n758), .C2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n741), .A2(new_n249), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1123), .B(KEYINPUT53), .ZN(new_n1124));
  INV_X1    g0924(.A(G125), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n1124), .B1(new_n785), .B2(new_n746), .C1(new_n1125), .C2(new_n762), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n1114), .A2(new_n1116), .B1(new_n1122), .B2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1111), .B1(new_n1127), .B2(new_n725), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n1109), .A2(new_n705), .B1(new_n1110), .B2(new_n1128), .ZN(new_n1129));
  AND3_X1   g0929(.A1(new_n1107), .A2(new_n1108), .A3(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1108), .B1(new_n1107), .B2(new_n1129), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(G378));
  INV_X1    g0933(.A(new_n889), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n265), .A2(new_n832), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n297), .A2(new_n353), .A3(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n353), .B1(new_n295), .B2(new_n296), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1137), .A2(new_n265), .A3(new_n832), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1139));
  AND3_X1   g0939(.A1(new_n1136), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1139), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n862), .A2(KEYINPUT40), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n867), .A2(new_n871), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1143), .B1(new_n1146), .B2(G330), .ZN(new_n1147));
  NOR3_X1   g0947(.A1(new_n872), .A2(new_n818), .A3(new_n1142), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1134), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1146), .A2(G330), .A3(new_n1143), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1142), .B1(new_n872), .B2(new_n818), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1150), .A2(new_n1151), .A3(new_n889), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1149), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1142), .A2(new_n711), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n706), .B1(G50), .B2(new_n801), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n793), .A2(G58), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1156), .B(KEYINPUT122), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n1157), .B1(new_n441), .B2(new_n738), .C1(new_n768), .C2(new_n762), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n274), .A2(G41), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1004), .A2(new_n916), .A3(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(G107), .B2(new_n787), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n362), .B2(new_n758), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n1158), .B(new_n1162), .C1(G97), .C2(new_n755), .ZN(new_n1163));
  OR2_X1    g0963(.A1(new_n1163), .A2(KEYINPUT58), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n785), .A2(new_n756), .B1(new_n758), .B2(new_n1119), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n742), .A2(new_n1120), .B1(new_n783), .B2(G150), .ZN(new_n1166));
  INV_X1    g0966(.A(G128), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n1166), .B1(new_n746), .B2(new_n1167), .C1(new_n1125), .C2(new_n738), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1165), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  OR2_X1    g0970(.A1(new_n1170), .A2(KEYINPUT59), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(KEYINPUT59), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n793), .A2(G159), .ZN(new_n1173));
  AOI211_X1 g0973(.A(G33), .B(G41), .C1(new_n731), .C2(G124), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .A4(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1163), .A2(KEYINPUT58), .ZN(new_n1176));
  AOI211_X1 g0976(.A(G50), .B(new_n1159), .C1(new_n269), .C2(new_n284), .ZN(new_n1177));
  XOR2_X1   g0977(.A(new_n1177), .B(KEYINPUT121), .Z(new_n1178));
  NAND4_X1  g0978(.A1(new_n1164), .A2(new_n1175), .A3(new_n1176), .A4(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1155), .B1(new_n1179), .B2(new_n725), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n1153), .A2(new_n705), .B1(new_n1154), .B2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1095), .B1(new_n1099), .B2(new_n1105), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1153), .A2(KEYINPUT57), .A3(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(new_n653), .ZN(new_n1184));
  AOI21_X1  g0984(.A(KEYINPUT57), .B1(new_n1153), .B2(new_n1182), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1181), .B1(new_n1184), .B2(new_n1185), .ZN(G375));
  NAND2_X1  g0986(.A1(new_n1065), .A2(KEYINPUT119), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1187), .A2(new_n1068), .A3(new_n810), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1075), .B1(new_n1188), .B2(new_n857), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1095), .B1(new_n1189), .B2(new_n1100), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1094), .B(new_n1062), .C1(new_n1069), .C2(new_n1075), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1190), .A2(new_n963), .A3(new_n1191), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n271), .B1(new_n751), .B2(new_n276), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n1007), .B(new_n1193), .C1(new_n763), .C2(G303), .ZN(new_n1194));
  OAI221_X1 g0994(.A(new_n1194), .B1(new_n441), .B2(new_n756), .C1(new_n357), .C2(new_n758), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n773), .A2(G97), .B1(G283), .B2(new_n787), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1196), .B1(new_n767), .B2(new_n738), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n271), .B1(new_n783), .B2(G50), .ZN(new_n1198));
  AND2_X1   g0998(.A1(new_n1157), .A2(new_n1198), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n1199), .B1(new_n249), .B2(new_n758), .C1(new_n756), .C2(new_n1121), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(G132), .A2(new_n739), .B1(new_n787), .B2(G137), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n1201), .B1(new_n1167), .B2(new_n762), .C1(new_n789), .C2(new_n772), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n1195), .A2(new_n1197), .B1(new_n1200), .B2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(new_n725), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1204), .B(new_n706), .C1(G68), .C2(new_n801), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(new_n857), .B2(new_n711), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(new_n1076), .B2(new_n705), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1192), .A2(new_n1207), .ZN(G381));
  NAND2_X1  g1008(.A1(new_n1107), .A2(new_n1129), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(G375), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  AND3_X1   g1011(.A1(new_n988), .A2(new_n780), .A3(new_n1020), .ZN(new_n1212));
  INV_X1    g1012(.A(G384), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(G390), .B1(KEYINPUT123), .B2(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(KEYINPUT123), .B2(new_n1214), .ZN(new_n1216));
  OR4_X1    g1016(.A1(G387), .A2(G381), .A3(new_n1211), .A4(new_n1216), .ZN(G407));
  NAND2_X1  g1017(.A1(new_n627), .A2(G213), .ZN(new_n1218));
  XOR2_X1   g1018(.A(new_n1218), .B(KEYINPUT124), .Z(new_n1219));
  OAI211_X1 g1019(.A(G407), .B(G213), .C1(new_n1211), .C2(new_n1219), .ZN(G409));
  NAND2_X1  g1020(.A1(new_n962), .A2(new_n963), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(new_n704), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n981), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n1222), .A2(new_n1223), .B1(new_n931), .B2(new_n923), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(G393), .A2(G396), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n988), .A2(new_n780), .A3(new_n1020), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n983), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1227), .A2(G390), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1050), .B1(new_n986), .B2(new_n960), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n958), .A2(KEYINPUT108), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n652), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1047), .B1(new_n1231), .B2(new_n1053), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n780), .B1(new_n988), .B2(new_n1020), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1212), .A2(new_n1233), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1232), .A2(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1224), .B1(new_n1228), .B2(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1232), .B1(new_n1234), .B2(new_n983), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1237), .B(new_n982), .C1(new_n1232), .C2(new_n1234), .ZN(new_n1238));
  AND2_X1   g1038(.A1(new_n1236), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(G2897), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1218), .A2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT60), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1191), .A2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1246), .A2(KEYINPUT60), .A3(new_n1094), .A4(new_n1062), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1245), .A2(new_n653), .A3(new_n1190), .A4(new_n1247), .ZN(new_n1248));
  AND3_X1   g1048(.A1(new_n1248), .A2(G384), .A3(new_n1207), .ZN(new_n1249));
  AOI21_X1  g1049(.A(G384), .B1(new_n1248), .B2(new_n1207), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT125), .ZN(new_n1251));
  NOR3_X1   g1051(.A1(new_n1249), .A2(new_n1250), .A3(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1248), .A2(new_n1207), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n1213), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1248), .A2(G384), .A3(new_n1207), .ZN(new_n1255));
  AOI21_X1  g1055(.A(KEYINPUT125), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1243), .B1(new_n1252), .B2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT127), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1219), .A2(new_n1241), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1257), .A2(new_n1258), .A3(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1251), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1254), .A2(KEYINPUT125), .A3(new_n1255), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1242), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  AOI211_X1 g1066(.A(new_n1241), .B(new_n1219), .C1(new_n1254), .C2(new_n1255), .ZN(new_n1267));
  OAI21_X1  g1067(.A(KEYINPUT127), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1153), .A2(new_n963), .A3(new_n1182), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1181), .A2(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1270), .A2(new_n1107), .A3(new_n1129), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1271), .B1(new_n1132), .B2(G375), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n1219), .ZN(new_n1273));
  AND3_X1   g1073(.A1(new_n1263), .A2(new_n1268), .A3(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1272), .A2(new_n1275), .A3(new_n1219), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(KEYINPUT62), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT61), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT62), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1272), .A2(new_n1275), .A3(new_n1279), .A4(new_n1218), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1277), .A2(new_n1278), .A3(new_n1280), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1240), .B1(new_n1274), .B2(new_n1281), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1272), .A2(new_n1275), .A3(KEYINPUT63), .A4(new_n1219), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1239), .A2(new_n1283), .A3(new_n1278), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1218), .ZN(new_n1285));
  OAI221_X1 g1085(.A(new_n1181), .B1(new_n1184), .B2(new_n1185), .C1(new_n1130), .C2(new_n1131), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1285), .B1(new_n1286), .B2(new_n1271), .ZN(new_n1287));
  AOI21_X1  g1087(.A(KEYINPUT63), .B1(new_n1287), .B2(new_n1275), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1284), .A2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT126), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1287), .A2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1272), .A2(new_n1218), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(KEYINPUT126), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1291), .A2(new_n1293), .A3(new_n1263), .A4(new_n1268), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1289), .A2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1282), .A2(new_n1295), .ZN(G405));
  AND3_X1   g1096(.A1(G375), .A2(new_n1107), .A3(new_n1129), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1132), .A2(G375), .ZN(new_n1298));
  NOR3_X1   g1098(.A1(new_n1297), .A2(new_n1298), .A3(new_n1259), .ZN(new_n1299));
  OR2_X1    g1099(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1299), .B1(new_n1275), .B2(new_n1300), .ZN(new_n1301));
  XNOR2_X1  g1101(.A(new_n1301), .B(new_n1239), .ZN(G402));
endmodule


