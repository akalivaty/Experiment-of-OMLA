//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 1 0 0 0 0 0 0 1 0 0 0 1 0 1 0 0 1 0 1 0 0 0 1 1 0 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 0 0 1 0 1 1 0 0 1 1 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:17 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n210, new_n211, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1277, new_n1278, new_n1279,
    new_n1280, new_n1281, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  NOR2_X1   g0009(.A1(G97), .A2(G107), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n211), .A2(G87), .ZN(G355));
  INV_X1    g0012(.A(G1), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(G13), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n217), .B(G250), .C1(G257), .C2(G264), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT0), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n206), .A2(new_n207), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n221), .A2(new_n214), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(KEYINPUT65), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n229));
  NAND3_X1  g0029(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n226), .A2(KEYINPUT65), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n216), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n219), .B(new_n223), .C1(KEYINPUT1), .C2(new_n232), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XOR2_X1   g0034(.A(G238), .B(G244), .Z(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G226), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT67), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G358));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n207), .A2(G68), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n202), .A2(G50), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G58), .B(G77), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n247), .B(new_n252), .Z(G351));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n221), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT70), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT70), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n254), .A2(new_n257), .A3(new_n221), .ZN(new_n258));
  AND2_X1   g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G13), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(G1), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G20), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  XOR2_X1   g0063(.A(KEYINPUT8), .B(G58), .Z(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(KEYINPUT71), .ZN(new_n265));
  XNOR2_X1  g0065(.A(KEYINPUT8), .B(G58), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT71), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n213), .A2(G20), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n265), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  XNOR2_X1  g0070(.A(new_n266), .B(KEYINPUT71), .ZN(new_n271));
  OAI22_X1  g0071(.A1(new_n263), .A2(new_n270), .B1(new_n262), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n255), .ZN(new_n273));
  AND2_X1   g0073(.A1(KEYINPUT3), .A2(G33), .ZN(new_n274));
  NOR2_X1   g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(KEYINPUT7), .B1(new_n276), .B2(new_n214), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT7), .ZN(new_n278));
  NOR4_X1   g0078(.A1(new_n274), .A2(new_n275), .A3(new_n278), .A4(G20), .ZN(new_n279));
  OAI21_X1  g0079(.A(G68), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G58), .A2(G68), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n203), .A2(new_n205), .A3(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(G20), .A2(G33), .ZN(new_n283));
  AOI22_X1  g0083(.A1(new_n282), .A2(G20), .B1(G159), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n280), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT16), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n273), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  OR2_X1    g0087(.A1(KEYINPUT3), .A2(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(KEYINPUT3), .A2(G33), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n288), .A2(KEYINPUT7), .A3(new_n214), .A4(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(KEYINPUT76), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT76), .ZN(new_n292));
  NAND4_X1  g0092(.A1(new_n276), .A2(new_n292), .A3(KEYINPUT7), .A4(new_n214), .ZN(new_n293));
  XNOR2_X1  g0093(.A(KEYINPUT3), .B(G33), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n278), .B1(new_n294), .B2(G20), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n291), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G68), .ZN(new_n297));
  AND2_X1   g0097(.A1(new_n284), .A2(KEYINPUT16), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n272), .B1(new_n287), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(G33), .A2(G41), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n301), .A2(G1), .A3(G13), .ZN(new_n302));
  INV_X1    g0102(.A(G223), .ZN(new_n303));
  INV_X1    g0103(.A(G1698), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G226), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G1698), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n305), .B(new_n307), .C1(new_n274), .C2(new_n275), .ZN(new_n308));
  NAND2_X1  g0108(.A1(G33), .A2(G87), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n302), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G41), .ZN(new_n311));
  INV_X1    g0111(.A(G45), .ZN(new_n312));
  AOI21_X1  g0112(.A(G1), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n313), .A2(new_n302), .A3(G274), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n213), .B1(G41), .B2(G45), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n302), .A2(G232), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G179), .ZN(new_n318));
  NOR3_X1   g0118(.A1(new_n310), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n308), .A2(new_n309), .ZN(new_n320));
  INV_X1    g0120(.A(new_n302), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n311), .A2(new_n312), .ZN(new_n323));
  AND2_X1   g0123(.A1(G1), .A2(G13), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n213), .A2(new_n323), .B1(new_n324), .B2(new_n301), .ZN(new_n325));
  INV_X1    g0125(.A(G274), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n326), .B1(new_n324), .B2(new_n301), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n325), .A2(G232), .B1(new_n327), .B2(new_n313), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n322), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n319), .B1(new_n329), .B2(G169), .ZN(new_n330));
  OAI21_X1  g0130(.A(KEYINPUT18), .B1(new_n300), .B2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n322), .A2(G190), .A3(new_n328), .ZN(new_n332));
  OAI21_X1  g0132(.A(G200), .B1(new_n310), .B2(new_n317), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI211_X1 g0134(.A(new_n272), .B(new_n334), .C1(new_n287), .C2(new_n299), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(KEYINPUT17), .ZN(new_n336));
  INV_X1    g0136(.A(new_n272), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n202), .B1(new_n295), .B2(new_n290), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n282), .A2(G20), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n283), .A2(G159), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n286), .B1(new_n338), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n255), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n284), .A2(KEYINPUT16), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n344), .B1(G68), .B2(new_n296), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n337), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT18), .ZN(new_n347));
  INV_X1    g0147(.A(new_n330), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n334), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n350), .B(new_n337), .C1(new_n343), .C2(new_n345), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT17), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AND4_X1   g0153(.A1(new_n331), .A2(new_n336), .A3(new_n349), .A4(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n208), .A2(G20), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n283), .A2(G150), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n265), .A2(new_n268), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT72), .ZN(new_n358));
  INV_X1    g0158(.A(G33), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n358), .B1(new_n359), .B2(G20), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n214), .A2(KEYINPUT72), .A3(G33), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n355), .B(new_n356), .C1(new_n357), .C2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n256), .A2(new_n258), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NOR3_X1   g0165(.A1(new_n260), .A2(new_n214), .A3(G1), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n269), .A2(G50), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n367), .A2(new_n369), .B1(new_n207), .B2(new_n366), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n365), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT9), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n365), .A2(new_n370), .A3(KEYINPUT9), .ZN(new_n374));
  INV_X1    g0174(.A(new_n314), .ZN(new_n375));
  XNOR2_X1  g0175(.A(KEYINPUT68), .B(G226), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n375), .B1(new_n325), .B2(new_n376), .ZN(new_n377));
  OAI211_X1 g0177(.A(G223), .B(G1698), .C1(new_n274), .C2(new_n275), .ZN(new_n378));
  INV_X1    g0178(.A(G77), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n378), .B1(new_n379), .B2(new_n294), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n294), .A2(new_n304), .ZN(new_n381));
  INV_X1    g0181(.A(G222), .ZN(new_n382));
  OAI21_X1  g0182(.A(KEYINPUT69), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(G1698), .B1(new_n288), .B2(new_n289), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT69), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n384), .A2(new_n385), .A3(G222), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n380), .B1(new_n383), .B2(new_n386), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n377), .B1(new_n387), .B2(new_n302), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(G200), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n373), .A2(new_n374), .A3(new_n389), .ZN(new_n390));
  OAI211_X1 g0190(.A(G190), .B(new_n377), .C1(new_n387), .C2(new_n302), .ZN(new_n391));
  XNOR2_X1  g0191(.A(new_n391), .B(KEYINPUT73), .ZN(new_n392));
  OAI21_X1  g0192(.A(KEYINPUT10), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT73), .ZN(new_n394));
  XNOR2_X1  g0194(.A(new_n391), .B(new_n394), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n371), .A2(new_n372), .B1(G200), .B2(new_n388), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT10), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n395), .A2(new_n396), .A3(new_n397), .A4(new_n374), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n393), .A2(new_n398), .ZN(new_n399));
  OR2_X1    g0199(.A1(new_n388), .A2(G179), .ZN(new_n400));
  INV_X1    g0200(.A(G169), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n388), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n400), .A2(new_n371), .A3(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n366), .A2(new_n255), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n405), .A2(G77), .A3(new_n269), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(G77), .B2(new_n262), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n264), .A2(new_n283), .B1(G20), .B2(G77), .ZN(new_n408));
  XNOR2_X1  g0208(.A(KEYINPUT15), .B(G87), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n410), .A2(new_n360), .A3(new_n361), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n273), .B1(new_n408), .B2(new_n411), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n407), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n294), .A2(G238), .A3(G1698), .ZN(new_n414));
  INV_X1    g0214(.A(G107), .ZN(new_n415));
  INV_X1    g0215(.A(G232), .ZN(new_n416));
  OAI221_X1 g0216(.A(new_n414), .B1(new_n415), .B2(new_n294), .C1(new_n381), .C2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n321), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n375), .B1(G244), .B2(new_n325), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(G190), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n413), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(G200), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n423), .B1(new_n418), .B2(new_n419), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n420), .A2(G179), .ZN(new_n426));
  AOI21_X1  g0226(.A(G169), .B1(new_n418), .B2(new_n419), .ZN(new_n427));
  NOR3_X1   g0227(.A1(new_n426), .A2(new_n413), .A3(new_n427), .ZN(new_n428));
  NOR3_X1   g0228(.A1(new_n404), .A2(new_n425), .A3(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT13), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n416), .A2(G1698), .ZN(new_n431));
  OAI221_X1 g0231(.A(new_n431), .B1(G226), .B2(G1698), .C1(new_n274), .C2(new_n275), .ZN(new_n432));
  NAND2_X1  g0232(.A1(G33), .A2(G97), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n321), .ZN(new_n435));
  INV_X1    g0235(.A(G238), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n302), .A2(new_n315), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n314), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n430), .B1(new_n435), .B2(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n302), .B1(new_n432), .B2(new_n433), .ZN(new_n441));
  NOR3_X1   g0241(.A1(new_n441), .A2(new_n438), .A3(KEYINPUT13), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n443), .A2(new_n423), .ZN(new_n444));
  AOI22_X1  g0244(.A1(new_n283), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n445), .B1(new_n362), .B2(new_n379), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n446), .A2(new_n364), .ZN(new_n447));
  OR2_X1    g0247(.A1(new_n447), .A2(KEYINPUT11), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(KEYINPUT11), .ZN(new_n449));
  OR3_X1    g0249(.A1(new_n262), .A2(KEYINPUT12), .A3(G68), .ZN(new_n450));
  OAI21_X1  g0250(.A(KEYINPUT12), .B1(new_n262), .B2(G68), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n202), .B1(new_n213), .B2(G20), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n450), .A2(new_n451), .B1(new_n405), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n448), .A2(new_n449), .A3(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT74), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(KEYINPUT13), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n435), .A2(new_n439), .A3(new_n456), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n455), .B(KEYINPUT13), .C1(new_n441), .C2(new_n438), .ZN(new_n458));
  AND3_X1   g0258(.A1(new_n457), .A2(new_n458), .A3(G190), .ZN(new_n459));
  NOR3_X1   g0259(.A1(new_n444), .A2(new_n454), .A3(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(KEYINPUT14), .B1(new_n443), .B2(new_n401), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT14), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n462), .B(G169), .C1(new_n440), .C2(new_n442), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n457), .A2(new_n458), .A3(G179), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT75), .ZN(new_n465));
  AND2_X1   g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n464), .A2(new_n465), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n461), .B(new_n463), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n460), .B1(new_n468), .B2(new_n454), .ZN(new_n469));
  AND4_X1   g0269(.A1(new_n354), .A2(new_n399), .A3(new_n429), .A4(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(G33), .A2(G283), .ZN(new_n471));
  OAI211_X1 g0271(.A(G250), .B(G1698), .C1(new_n274), .C2(new_n275), .ZN(new_n472));
  OAI211_X1 g0272(.A(G244), .B(new_n304), .C1(new_n274), .C2(new_n275), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT4), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n471), .B(new_n472), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(KEYINPUT4), .B1(new_n384), .B2(G244), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n321), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n213), .A2(G45), .ZN(new_n478));
  OR2_X1    g0278(.A1(KEYINPUT5), .A2(G41), .ZN(new_n479));
  NAND2_X1  g0279(.A1(KEYINPUT5), .A2(G41), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n327), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n312), .A2(G1), .ZN(new_n483));
  INV_X1    g0283(.A(new_n480), .ZN(new_n484));
  NOR2_X1   g0284(.A1(KEYINPUT5), .A2(G41), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AND3_X1   g0286(.A1(new_n486), .A2(G257), .A3(new_n302), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n477), .A2(new_n482), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n401), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT6), .ZN(new_n491));
  AND2_X1   g0291(.A1(G97), .A2(G107), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n491), .B1(new_n492), .B2(new_n210), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n415), .A2(KEYINPUT6), .A3(G97), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(G20), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n283), .A2(G77), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n415), .B1(new_n295), .B2(new_n290), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n255), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(G97), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n213), .A2(new_n501), .A3(G13), .A4(G20), .ZN(new_n502));
  XNOR2_X1  g0302(.A(new_n502), .B(KEYINPUT77), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n213), .A2(G33), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n256), .A2(new_n262), .A3(new_n258), .A4(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n503), .B1(new_n505), .B2(new_n501), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n500), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n473), .A2(new_n474), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n294), .A2(KEYINPUT4), .A3(G244), .A4(new_n304), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n509), .A2(new_n510), .A3(new_n471), .A4(new_n472), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n487), .B1(new_n511), .B2(new_n321), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n512), .A2(new_n318), .A3(new_n482), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n490), .A2(new_n508), .A3(new_n513), .ZN(new_n514));
  OAI21_X1  g0314(.A(G107), .B1(new_n277), .B2(new_n279), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n495), .A2(G20), .B1(G77), .B2(new_n283), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n506), .B1(new_n517), .B2(new_n255), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n477), .A2(G190), .A3(new_n482), .A4(new_n488), .ZN(new_n519));
  INV_X1    g0319(.A(new_n482), .ZN(new_n520));
  AOI211_X1 g0320(.A(new_n487), .B(new_n520), .C1(new_n511), .C2(new_n321), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n518), .B(new_n519), .C1(new_n521), .C2(new_n423), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n514), .A2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT79), .ZN(new_n525));
  XNOR2_X1  g0325(.A(KEYINPUT5), .B(G41), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n526), .A2(new_n483), .B1(new_n324), .B2(new_n301), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n527), .A2(G270), .B1(new_n327), .B2(new_n481), .ZN(new_n528));
  OAI211_X1 g0328(.A(G264), .B(G1698), .C1(new_n274), .C2(new_n275), .ZN(new_n529));
  OAI211_X1 g0329(.A(G257), .B(new_n304), .C1(new_n274), .C2(new_n275), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n288), .A2(G303), .A3(new_n289), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n321), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n423), .B1(new_n528), .B2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(G116), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT78), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT78), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(G116), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n536), .A2(new_n538), .A3(G20), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n471), .B(new_n214), .C1(G33), .C2(new_n501), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n539), .A2(new_n255), .A3(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT20), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n539), .A2(KEYINPUT20), .A3(new_n255), .A4(new_n540), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n504), .A2(G116), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(new_n539), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n405), .A2(new_n547), .B1(new_n548), .B2(new_n261), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n545), .A2(new_n549), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n525), .B1(new_n534), .B2(new_n550), .ZN(new_n551));
  XNOR2_X1  g0351(.A(KEYINPUT78), .B(G116), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n552), .A2(G20), .A3(new_n261), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n273), .A2(new_n262), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n553), .B1(new_n554), .B2(new_n546), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n555), .B1(new_n543), .B2(new_n544), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n486), .A2(G270), .A3(new_n302), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n482), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n558), .B1(new_n321), .B2(new_n532), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n556), .B(KEYINPUT79), .C1(new_n559), .C2(new_n423), .ZN(new_n560));
  INV_X1    g0360(.A(new_n559), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n551), .B(new_n560), .C1(new_n421), .C2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n360), .A2(G97), .A3(new_n361), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT19), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n294), .A2(new_n214), .A3(G68), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n214), .B1(new_n433), .B2(new_n564), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n567), .B1(G87), .B2(new_n211), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n565), .A2(new_n566), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n255), .ZN(new_n570));
  INV_X1    g0370(.A(new_n505), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n410), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n409), .A2(new_n366), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n570), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n537), .A2(G116), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n535), .A2(KEYINPUT78), .ZN(new_n576));
  OAI21_X1  g0376(.A(G33), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  OAI211_X1 g0377(.A(G238), .B(new_n304), .C1(new_n274), .C2(new_n275), .ZN(new_n578));
  OAI211_X1 g0378(.A(G244), .B(G1698), .C1(new_n274), .C2(new_n275), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n321), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n302), .A2(G274), .A3(new_n483), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n302), .A2(G250), .A3(new_n478), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n401), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n584), .B1(new_n580), .B2(new_n321), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n318), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n574), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n586), .A2(G200), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n569), .A2(new_n255), .B1(new_n366), .B2(new_n409), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n571), .A2(G87), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n588), .A2(G190), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n591), .A2(new_n592), .A3(new_n593), .A4(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n486), .A2(G264), .A3(new_n302), .ZN(new_n596));
  AND2_X1   g0396(.A1(new_n596), .A2(new_n482), .ZN(new_n597));
  OAI211_X1 g0397(.A(G257), .B(G1698), .C1(new_n274), .C2(new_n275), .ZN(new_n598));
  OAI211_X1 g0398(.A(G250), .B(new_n304), .C1(new_n274), .C2(new_n275), .ZN(new_n599));
  INV_X1    g0399(.A(G294), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n598), .B(new_n599), .C1(new_n359), .C2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n321), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n597), .A2(new_n602), .A3(new_n421), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n596), .A2(new_n482), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n604), .B1(new_n321), .B2(new_n601), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n603), .B1(new_n605), .B2(G200), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n214), .B(G87), .C1(new_n274), .C2(new_n275), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(KEYINPUT22), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT22), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n294), .A2(new_n609), .A3(new_n214), .A4(G87), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT24), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n359), .B1(new_n536), .B2(new_n538), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT23), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n614), .B1(new_n214), .B2(G107), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n415), .A2(KEYINPUT23), .A3(G20), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n613), .A2(new_n214), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  AND3_X1   g0417(.A1(new_n611), .A2(new_n612), .A3(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n612), .B1(new_n611), .B2(new_n617), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n255), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n366), .A2(new_n415), .ZN(new_n621));
  XNOR2_X1  g0421(.A(new_n621), .B(KEYINPUT25), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n505), .A2(new_n415), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n606), .A2(new_n620), .A3(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n562), .A2(new_n590), .A3(new_n595), .A4(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n597), .A2(new_n602), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n401), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n597), .A2(new_n602), .A3(new_n318), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n611), .A2(new_n617), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(KEYINPUT24), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n611), .A2(new_n612), .A3(new_n617), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n273), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n624), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n628), .B(new_n629), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n528), .A2(G179), .A3(new_n533), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n550), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n401), .B1(new_n528), .B2(new_n533), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n638), .A2(new_n550), .A3(KEYINPUT21), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n638), .A2(new_n550), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT21), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n635), .A2(new_n640), .A3(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n626), .A2(new_n644), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n470), .A2(new_n524), .A3(new_n645), .ZN(G372));
  INV_X1    g0446(.A(new_n590), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n490), .A2(new_n513), .A3(new_n508), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n648), .A2(KEYINPUT26), .A3(new_n590), .A4(new_n595), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT26), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n595), .A2(new_n590), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n650), .B1(new_n651), .B2(new_n514), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n647), .B1(new_n649), .B2(new_n652), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n625), .A2(new_n590), .A3(new_n595), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n524), .A2(new_n654), .A3(new_n644), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n470), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g0457(.A(new_n657), .B(KEYINPUT80), .Z(new_n658));
  INV_X1    g0458(.A(KEYINPUT82), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n399), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n393), .A2(KEYINPUT82), .A3(new_n398), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT81), .ZN(new_n663));
  NOR3_X1   g0463(.A1(new_n300), .A2(KEYINPUT18), .A3(new_n330), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n347), .B1(new_n346), .B2(new_n348), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n663), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n331), .A2(new_n349), .A3(KEYINPUT81), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n336), .A2(new_n353), .ZN(new_n669));
  INV_X1    g0469(.A(new_n460), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n428), .B1(new_n468), .B2(new_n454), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n668), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n404), .B1(new_n662), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n658), .A2(new_n674), .ZN(G369));
  NAND2_X1  g0475(.A1(new_n261), .A2(new_n214), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n676), .A2(KEYINPUT27), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(KEYINPUT27), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(G213), .A3(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(G343), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n682), .B1(new_n633), .B2(new_n634), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n635), .A2(new_n625), .A3(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT83), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n629), .B1(new_n605), .B2(G169), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n687), .B1(new_n620), .B2(new_n624), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n682), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n684), .A2(new_n685), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n686), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT84), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n686), .A2(KEYINPUT84), .A3(new_n689), .A4(new_n690), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n643), .A2(new_n637), .A3(new_n639), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(new_n681), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  AOI22_X1  g0498(.A1(new_n695), .A2(new_n698), .B1(new_n688), .B2(new_n681), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n696), .A2(new_n550), .A3(new_n682), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n562), .B1(new_n556), .B2(new_n681), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n700), .B1(new_n701), .B2(new_n696), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(G330), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n695), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n699), .A2(new_n705), .ZN(G399));
  INV_X1    g0506(.A(new_n217), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(G41), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR3_X1   g0509(.A1(new_n211), .A2(G87), .A3(G116), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(G1), .A3(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n220), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n711), .B1(new_n712), .B2(new_n709), .ZN(new_n713));
  XNOR2_X1  g0513(.A(new_n713), .B(KEYINPUT28), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT29), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n523), .A2(KEYINPUT86), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT86), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n514), .A2(new_n522), .A3(new_n717), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n716), .A2(new_n654), .A3(new_n644), .A4(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n653), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n715), .B1(new_n720), .B2(new_n681), .ZN(new_n721));
  AOI211_X1 g0521(.A(KEYINPUT29), .B(new_n682), .C1(new_n653), .C2(new_n655), .ZN(new_n722));
  OR2_X1    g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n696), .A2(new_n688), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n724), .A2(new_n654), .A3(new_n524), .A4(new_n562), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT85), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n636), .A2(new_n512), .A3(new_n605), .A4(new_n588), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT30), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n627), .A2(new_n586), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n730), .A2(KEYINPUT30), .A3(new_n512), .A4(new_n636), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n588), .A2(G179), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n561), .A2(new_n489), .A3(new_n627), .A4(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n729), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(KEYINPUT31), .B1(new_n734), .B2(new_n682), .ZN(new_n735));
  OAI22_X1  g0535(.A1(new_n725), .A2(new_n682), .B1(new_n726), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n734), .A2(new_n682), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT31), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n734), .A2(KEYINPUT31), .A3(new_n682), .ZN(new_n740));
  AOI21_X1  g0540(.A(KEYINPUT85), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OR2_X1    g0541(.A1(new_n736), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n723), .B1(G330), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n714), .B1(new_n743), .B2(G1), .ZN(new_n744));
  XOR2_X1   g0544(.A(new_n744), .B(KEYINPUT87), .Z(G364));
  NOR2_X1   g0545(.A1(new_n260), .A2(G20), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n213), .B1(new_n746), .B2(G45), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n708), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n707), .A2(new_n276), .ZN(new_n751));
  AOI22_X1  g0551(.A1(new_n751), .A2(G355), .B1(new_n535), .B2(new_n707), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n707), .A2(new_n294), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n753), .B1(new_n712), .B2(G45), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n252), .A2(new_n312), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n752), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(G13), .A2(G33), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(G20), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n221), .B1(G20), .B2(new_n401), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n750), .B1(new_n756), .B2(new_n761), .ZN(new_n762));
  XNOR2_X1  g0562(.A(new_n762), .B(KEYINPUT88), .ZN(new_n763));
  INV_X1    g0563(.A(new_n759), .ZN(new_n764));
  NOR4_X1   g0564(.A1(new_n214), .A2(new_n421), .A3(new_n423), .A4(G179), .ZN(new_n765));
  XOR2_X1   g0565(.A(new_n765), .B(KEYINPUT91), .Z(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G303), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G179), .A2(G200), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n214), .B1(new_n768), .B2(G190), .ZN(new_n769));
  OAI211_X1 g0569(.A(new_n767), .B(new_n276), .C1(new_n600), .C2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(G20), .A2(G179), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(KEYINPUT89), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G190), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n423), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n770), .B1(G326), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n421), .A2(G20), .ZN(new_n776));
  INV_X1    g0576(.A(KEYINPUT90), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NOR3_X1   g0578(.A1(new_n778), .A2(G179), .A3(new_n423), .ZN(new_n779));
  INV_X1    g0579(.A(new_n768), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  AOI22_X1  g0581(.A1(new_n779), .A2(G283), .B1(new_n781), .B2(G329), .ZN(new_n782));
  XNOR2_X1  g0582(.A(new_n782), .B(KEYINPUT92), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n773), .A2(G200), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G322), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n772), .A2(new_n421), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(G200), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(new_n423), .ZN(new_n788));
  XNOR2_X1  g0588(.A(KEYINPUT33), .B(G317), .ZN(new_n789));
  AOI22_X1  g0589(.A1(G311), .A2(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n775), .A2(new_n783), .A3(new_n785), .A4(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n765), .ZN(new_n792));
  INV_X1    g0592(.A(G87), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n294), .B1(new_n501), .B2(new_n769), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n779), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(new_n415), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n794), .B(new_n796), .C1(new_n788), .C2(G68), .ZN(new_n797));
  INV_X1    g0597(.A(new_n784), .ZN(new_n798));
  INV_X1    g0598(.A(new_n787), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n201), .A2(new_n798), .B1(new_n799), .B2(new_n379), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n800), .B1(G50), .B2(new_n774), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n781), .A2(G159), .ZN(new_n802));
  XOR2_X1   g0602(.A(new_n802), .B(KEYINPUT32), .Z(new_n803));
  NAND3_X1  g0603(.A1(new_n797), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n791), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n760), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n763), .B1(new_n702), .B2(new_n764), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n702), .A2(G330), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n703), .A2(new_n750), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  XNOR2_X1  g0610(.A(KEYINPUT93), .B(KEYINPUT94), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n810), .B(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(G396));
  NAND2_X1  g0613(.A1(new_n742), .A2(G330), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n656), .A2(new_n681), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n422), .A2(new_n424), .B1(new_n413), .B2(new_n681), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n427), .A2(new_n413), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(G179), .B2(new_n420), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n428), .A2(new_n681), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n815), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n821), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n656), .A2(new_n681), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n749), .B1(new_n814), .B2(new_n825), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(new_n814), .B2(new_n825), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n760), .A2(new_n757), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n749), .B1(G77), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n795), .A2(new_n202), .ZN(new_n831));
  INV_X1    g0631(.A(new_n781), .ZN(new_n832));
  INV_X1    g0632(.A(G132), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n294), .B1(new_n201), .B2(new_n769), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n831), .B(new_n834), .C1(G50), .C2(new_n766), .ZN(new_n835));
  AOI22_X1  g0635(.A1(G137), .A2(new_n774), .B1(new_n788), .B2(G150), .ZN(new_n836));
  AOI22_X1  g0636(.A1(G143), .A2(new_n784), .B1(new_n787), .B2(G159), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g0638(.A(KEYINPUT96), .B(KEYINPUT34), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n835), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n838), .A2(new_n839), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n795), .A2(new_n793), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(G311), .B2(new_n781), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n766), .A2(G107), .ZN(new_n844));
  INV_X1    g0644(.A(new_n769), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n294), .B1(new_n845), .B2(G97), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n843), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  XOR2_X1   g0647(.A(KEYINPUT95), .B(G283), .Z(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  AOI22_X1  g0649(.A1(G303), .A2(new_n774), .B1(new_n788), .B2(new_n849), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n850), .B1(new_n600), .B2(new_n798), .C1(new_n552), .C2(new_n799), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n840), .A2(new_n841), .B1(new_n847), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n830), .B1(new_n852), .B2(new_n760), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n758), .B2(new_n823), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n827), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(G384));
  NOR2_X1   g0656(.A1(new_n746), .A2(new_n213), .ZN(new_n857));
  INV_X1    g0657(.A(G330), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT101), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n341), .B1(new_n296), .B2(G68), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n299), .B(new_n364), .C1(KEYINPUT16), .C2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n330), .B1(new_n861), .B2(new_n337), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n859), .B1(new_n862), .B2(new_n335), .ZN(new_n863));
  OR2_X1    g0663(.A1(new_n860), .A2(KEYINPUT16), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n259), .B1(new_n297), .B2(new_n298), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n272), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n351), .B(KEYINPUT101), .C1(new_n866), .C2(new_n330), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n861), .A2(new_n337), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT100), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n868), .A2(new_n869), .A3(new_n680), .ZN(new_n870));
  OAI21_X1  g0670(.A(KEYINPUT100), .B1(new_n866), .B2(new_n679), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n863), .A2(new_n867), .A3(new_n870), .A4(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(KEYINPUT37), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n300), .A2(new_n679), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT37), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n346), .A2(new_n348), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n875), .A2(new_n876), .A3(new_n877), .A4(new_n351), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n873), .A2(new_n878), .ZN(new_n879));
  AND2_X1   g0679(.A1(new_n871), .A2(new_n870), .ZN(new_n880));
  OR2_X1    g0680(.A1(new_n354), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n879), .A2(KEYINPUT38), .A3(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT38), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n877), .A2(new_n351), .ZN(new_n884));
  NOR3_X1   g0684(.A1(new_n884), .A2(new_n874), .A3(KEYINPUT37), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n885), .B1(new_n872), .B2(KEYINPUT37), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n354), .A2(new_n880), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n883), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n882), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n740), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n890), .A2(new_n735), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n645), .A2(new_n524), .A3(new_n681), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n468), .A2(new_n454), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n454), .A2(new_n682), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n894), .A2(new_n670), .A3(new_n895), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n454), .B(new_n682), .C1(new_n468), .C2(new_n460), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n821), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n893), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(KEYINPUT40), .B1(new_n889), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n875), .B1(new_n668), .B2(new_n669), .ZN(new_n901));
  OAI21_X1  g0701(.A(KEYINPUT37), .B1(new_n884), .B2(new_n874), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n878), .A2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n883), .B1(new_n901), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n882), .A2(new_n905), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n893), .A2(new_n898), .A3(KEYINPUT40), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n900), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n470), .A2(new_n893), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n858), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n910), .B1(new_n908), .B2(new_n909), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n668), .A2(new_n680), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n824), .A2(new_n820), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n896), .A2(new_n897), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n912), .B1(new_n916), .B2(new_n889), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT39), .ZN(new_n918));
  NOR3_X1   g0718(.A1(new_n886), .A2(new_n887), .A3(new_n883), .ZN(new_n919));
  AND3_X1   g0719(.A1(new_n331), .A2(new_n349), .A3(KEYINPUT81), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT81), .B1(new_n331), .B2(new_n349), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n669), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n874), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT38), .B1(new_n923), .B2(new_n903), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n918), .B1(new_n919), .B2(new_n924), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n894), .A2(new_n682), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n882), .A2(KEYINPUT39), .A3(new_n888), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n917), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n470), .B1(new_n721), .B2(new_n722), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n674), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n929), .B(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n857), .B1(new_n911), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n932), .B2(new_n911), .ZN(new_n934));
  OR2_X1    g0734(.A1(new_n495), .A2(KEYINPUT35), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n495), .A2(KEYINPUT35), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n935), .A2(G116), .A3(new_n222), .A4(new_n936), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT36), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n220), .A2(G77), .A3(new_n281), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT97), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  XOR2_X1   g0741(.A(new_n248), .B(KEYINPUT98), .Z(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n939), .B2(new_n940), .ZN(new_n943));
  OAI211_X1 g0743(.A(G1), .B(new_n260), .C1(new_n941), .C2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n938), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(KEYINPUT99), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n934), .A2(new_n946), .ZN(G367));
  OAI21_X1  g0747(.A(new_n761), .B1(new_n217), .B2(new_n409), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n948), .B1(new_n753), .B2(new_n243), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n294), .B1(new_n845), .B2(G107), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n792), .A2(new_n552), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n950), .B1(new_n951), .B2(KEYINPUT46), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n766), .A2(KEYINPUT46), .A3(G116), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n779), .A2(G97), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n781), .A2(G317), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  AOI211_X1 g0756(.A(new_n952), .B(new_n956), .C1(G311), .C2(new_n774), .ZN(new_n957));
  AOI22_X1  g0757(.A1(G303), .A2(new_n784), .B1(new_n787), .B2(new_n849), .ZN(new_n958));
  INV_X1    g0758(.A(new_n788), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n957), .B(new_n958), .C1(new_n600), .C2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n779), .A2(G77), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n781), .A2(G137), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n845), .A2(G68), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n276), .B1(new_n765), .B2(G58), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n961), .A2(new_n962), .A3(new_n963), .A4(new_n964), .ZN(new_n965));
  AOI22_X1  g0765(.A1(G50), .A2(new_n787), .B1(new_n774), .B2(G143), .ZN(new_n966));
  INV_X1    g0766(.A(G150), .ZN(new_n967));
  INV_X1    g0767(.A(G159), .ZN(new_n968));
  OAI221_X1 g0768(.A(new_n966), .B1(new_n967), .B2(new_n798), .C1(new_n968), .C2(new_n959), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n960), .B1(new_n965), .B2(new_n969), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT47), .ZN(new_n971));
  AOI211_X1 g0771(.A(new_n750), .B(new_n949), .C1(new_n971), .C2(new_n760), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n592), .A2(new_n593), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n973), .A2(new_n681), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n651), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n647), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n759), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n972), .A2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT45), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n695), .A2(new_n698), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n688), .A2(new_n681), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n716), .B(new_n718), .C1(new_n518), .C2(new_n681), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n648), .A2(new_n682), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n981), .B1(new_n984), .B2(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n699), .A2(KEYINPUT45), .A3(new_n987), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n984), .A2(KEYINPUT44), .A3(new_n988), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT44), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n699), .B2(new_n987), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n991), .A2(new_n705), .A3(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n695), .A2(new_n698), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n697), .B1(new_n693), .B2(new_n694), .ZN(new_n998));
  OR3_X1    g0798(.A1(new_n997), .A2(new_n703), .A3(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n703), .B1(new_n997), .B2(new_n998), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n743), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT103), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n705), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n996), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n990), .A2(new_n989), .B1(new_n992), .B2(new_n994), .ZN(new_n1007));
  NOR3_X1   g0807(.A1(new_n1007), .A2(new_n1004), .A3(new_n705), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n743), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n708), .B(KEYINPUT41), .Z(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n748), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n985), .A2(new_n635), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n682), .B1(new_n1013), .B2(new_n514), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT42), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n982), .B2(new_n988), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n998), .A2(KEYINPUT42), .A3(new_n987), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1014), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  AND2_X1   g0818(.A1(new_n978), .A2(KEYINPUT102), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n978), .A2(KEYINPUT102), .ZN(new_n1020));
  NOR3_X1   g0820(.A1(new_n1019), .A2(new_n1020), .A3(KEYINPUT43), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1021), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT43), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1023), .B1(new_n1024), .B2(new_n978), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1022), .B1(new_n1018), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n695), .A2(new_n704), .A3(new_n987), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n980), .B1(new_n1012), .B2(new_n1030), .ZN(G387));
  NOR2_X1   g0831(.A1(new_n1003), .A2(new_n709), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1001), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1032), .B1(new_n743), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n710), .ZN(new_n1035));
  AOI211_X1 g0835(.A(G45), .B(new_n1035), .C1(G68), .C2(G77), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n264), .A2(new_n207), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT50), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n753), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n1040), .A2(KEYINPUT104), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(KEYINPUT104), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n1041), .B(new_n1042), .C1(new_n312), .C2(new_n239), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n751), .A2(new_n1035), .B1(new_n415), .B2(new_n707), .ZN(new_n1044));
  AOI21_X1  g0844(.A(KEYINPUT105), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NOR3_X1   g0845(.A1(new_n1045), .A2(new_n759), .A3(new_n760), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1043), .A2(KEYINPUT105), .A3(new_n1044), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n750), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(G68), .A2(new_n787), .B1(new_n788), .B2(new_n271), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT106), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n845), .A2(new_n410), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n276), .B1(new_n765), .B2(G77), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n954), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(G150), .B2(new_n781), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(G50), .A2(new_n784), .B1(new_n774), .B2(G159), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1050), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n294), .B1(new_n781), .B2(G326), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n792), .A2(new_n600), .B1(new_n769), .B2(new_n848), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(G303), .A2(new_n787), .B1(new_n784), .B2(G317), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(G311), .A2(new_n788), .B1(new_n774), .B2(G322), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT48), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1058), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(new_n1062), .B2(new_n1061), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT49), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1057), .B1(new_n552), .B2(new_n795), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  AND2_X1   g0866(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1056), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1068), .A2(new_n760), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1048), .B(new_n1069), .C1(new_n695), .C2(new_n764), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1034), .B(new_n1070), .C1(new_n747), .C2(new_n1001), .ZN(G393));
  AND3_X1   g0871(.A1(new_n991), .A2(new_n705), .A3(new_n995), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n705), .B1(new_n991), .B2(new_n995), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n1072), .A2(new_n1073), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1074), .B(new_n708), .C1(new_n1008), .C2(new_n1006), .ZN(new_n1075));
  AND2_X1   g0875(.A1(new_n753), .A2(new_n247), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n761), .B1(new_n501), .B2(new_n217), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n276), .B(new_n842), .C1(G77), .C2(new_n845), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n1078), .B1(new_n207), .B2(new_n959), .C1(new_n266), .C2(new_n799), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(G150), .A2(new_n774), .B1(new_n784), .B2(G159), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT107), .ZN(new_n1081));
  AND2_X1   g0881(.A1(new_n1081), .A2(KEYINPUT51), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n781), .A2(G143), .B1(G68), .B2(new_n765), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT108), .ZN(new_n1084));
  NOR3_X1   g0884(.A1(new_n1079), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(KEYINPUT51), .B2(new_n1081), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n294), .B(new_n796), .C1(new_n765), .C2(new_n849), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n781), .A2(G322), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1087), .B(new_n1088), .C1(new_n600), .C2(new_n799), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n788), .A2(G303), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n552), .B2(new_n769), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1089), .B1(KEYINPUT109), .B2(new_n1091), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(G311), .A2(new_n784), .B1(new_n774), .B2(G317), .ZN(new_n1093));
  XOR2_X1   g0893(.A(new_n1093), .B(KEYINPUT52), .Z(new_n1094));
  OAI211_X1 g0894(.A(new_n1092), .B(new_n1094), .C1(KEYINPUT109), .C2(new_n1091), .ZN(new_n1095));
  AND2_X1   g0895(.A1(new_n1086), .A2(new_n1095), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n749), .B1(new_n1076), .B2(new_n1077), .C1(new_n1096), .C2(new_n806), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(new_n759), .B2(new_n988), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1098), .B1(new_n1099), .B2(new_n748), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1075), .A2(KEYINPUT110), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(KEYINPUT110), .B1(new_n1075), .B2(new_n1100), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(G390));
  AOI21_X1  g0905(.A(new_n858), .B1(new_n891), .B2(new_n892), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n898), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n824), .A2(new_n820), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n926), .B1(new_n1109), .B2(new_n914), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(new_n925), .B2(new_n927), .ZN(new_n1111));
  AND3_X1   g0911(.A1(new_n720), .A2(new_n681), .A3(new_n819), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n820), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n914), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n926), .ZN(new_n1115));
  AND3_X1   g0915(.A1(new_n906), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1108), .B1(new_n1111), .B2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1115), .B1(new_n913), .B2(new_n915), .ZN(new_n1118));
  AND3_X1   g0918(.A1(new_n882), .A2(KEYINPUT39), .A3(new_n888), .ZN(new_n1119));
  AOI21_X1  g0919(.A(KEYINPUT39), .B1(new_n882), .B2(new_n905), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1118), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n906), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n898), .B(G330), .C1(new_n736), .C2(new_n741), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1121), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1117), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n739), .A2(new_n740), .ZN(new_n1126));
  NOR4_X1   g0926(.A1(new_n626), .A2(new_n644), .A3(new_n523), .A4(new_n682), .ZN(new_n1127));
  OAI211_X1 g0927(.A(G330), .B(new_n823), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n915), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n682), .B1(new_n653), .B2(new_n719), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1113), .B1(new_n1130), .B2(new_n819), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1129), .A2(new_n1123), .A3(new_n1131), .ZN(new_n1132));
  OAI211_X1 g0932(.A(G330), .B(new_n823), .C1(new_n736), .C2(new_n741), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n1133), .A2(new_n915), .B1(new_n898), .B2(new_n1106), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1132), .B1(new_n1134), .B2(new_n913), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1106), .A2(new_n470), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n930), .A2(new_n674), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT111), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n930), .A2(new_n674), .A3(new_n1136), .A4(KEYINPUT111), .ZN(new_n1140));
  AND3_X1   g0940(.A1(new_n1135), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1125), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1141), .A2(new_n1117), .A3(new_n1124), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1143), .A2(new_n708), .A3(new_n1144), .ZN(new_n1145));
  AND2_X1   g0945(.A1(new_n1117), .A2(new_n1124), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n757), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n749), .B1(new_n271), .B2(new_n829), .ZN(new_n1148));
  AOI211_X1 g0948(.A(new_n294), .B(new_n831), .C1(G77), .C2(new_n845), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n766), .A2(G87), .B1(G294), .B2(new_n781), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(G97), .A2(new_n787), .B1(new_n774), .B2(G283), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(G107), .A2(new_n788), .B1(new_n784), .B2(G116), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .A4(new_n1152), .ZN(new_n1153));
  OR3_X1    g0953(.A1(new_n792), .A2(KEYINPUT53), .A3(new_n967), .ZN(new_n1154));
  OAI21_X1  g0954(.A(KEYINPUT53), .B1(new_n792), .B2(new_n967), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1154), .B(new_n1155), .C1(new_n968), .C2(new_n769), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(G128), .B2(new_n774), .ZN(new_n1157));
  XOR2_X1   g0957(.A(KEYINPUT54), .B(G143), .Z(new_n1158));
  AOI22_X1  g0958(.A1(G137), .A2(new_n788), .B1(new_n787), .B2(new_n1158), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1157), .B(new_n1159), .C1(new_n833), .C2(new_n798), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n276), .B1(new_n781), .B2(G125), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n795), .B2(new_n207), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1162), .B(KEYINPUT112), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1153), .B1(new_n1160), .B2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1148), .B1(new_n1164), .B2(new_n760), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n1146), .A2(new_n748), .B1(new_n1147), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1145), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(KEYINPUT113), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT113), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1145), .A2(new_n1166), .A3(new_n1169), .ZN(new_n1170));
  AND2_X1   g0970(.A1(new_n1168), .A2(new_n1170), .ZN(G378));
  NAND2_X1  g0971(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1144), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n661), .ZN(new_n1175));
  AOI21_X1  g0975(.A(KEYINPUT82), .B1(new_n393), .B2(new_n398), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n403), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n371), .A2(new_n680), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n662), .A2(new_n403), .A3(new_n1178), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1182), .A2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1180), .A2(new_n1181), .A3(new_n1183), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n906), .A2(new_n907), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(G330), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1187), .B1(new_n1189), .B2(new_n900), .ZN(new_n1190));
  AND3_X1   g0990(.A1(new_n1180), .A2(new_n1181), .A3(new_n1183), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1183), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n889), .A2(new_n899), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT40), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n858), .B1(new_n906), .B2(new_n907), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1193), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1190), .A2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(new_n929), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1190), .A2(new_n1198), .A3(new_n928), .A4(new_n917), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1174), .A2(KEYINPUT57), .A3(new_n1200), .A4(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n929), .A2(KEYINPUT118), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1199), .A2(new_n1203), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1190), .A2(new_n1198), .A3(new_n929), .A4(KEYINPUT118), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n1204), .A2(new_n1205), .B1(new_n1144), .B2(new_n1173), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1202), .B(new_n708), .C1(KEYINPUT57), .C2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n747), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1193), .A2(new_n757), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n749), .B1(G50), .B2(new_n829), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(G132), .A2(new_n788), .B1(new_n787), .B2(G137), .ZN(new_n1211));
  XOR2_X1   g1011(.A(new_n1211), .B(KEYINPUT116), .Z(new_n1212));
  NAND2_X1  g1012(.A1(new_n774), .A2(G125), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n784), .A2(G128), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n765), .A2(new_n1158), .B1(new_n845), .B2(G150), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .A4(new_n1215), .ZN(new_n1216));
  XOR2_X1   g1016(.A(new_n1216), .B(KEYINPUT59), .Z(new_n1217));
  NAND2_X1  g1017(.A1(new_n779), .A2(G159), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(G33), .A2(G41), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1219), .B(KEYINPUT114), .ZN(new_n1220));
  XOR2_X1   g1020(.A(KEYINPUT117), .B(G124), .Z(new_n1221));
  NAND2_X1  g1021(.A1(new_n781), .A2(new_n1221), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1217), .A2(new_n1218), .A3(new_n1220), .A4(new_n1222), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(G116), .A2(new_n774), .B1(new_n787), .B2(new_n410), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1224), .B1(new_n501), .B2(new_n959), .C1(new_n415), .C2(new_n798), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n795), .A2(new_n201), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n781), .A2(G283), .ZN(new_n1227));
  AOI211_X1 g1027(.A(G41), .B(new_n294), .C1(new_n765), .C2(G77), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1227), .A2(new_n1228), .A3(new_n963), .ZN(new_n1229));
  NOR3_X1   g1029(.A1(new_n1225), .A2(new_n1226), .A3(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1230), .A2(KEYINPUT58), .ZN(new_n1231));
  OR2_X1    g1031(.A1(new_n1230), .A2(KEYINPUT58), .ZN(new_n1232));
  AOI211_X1 g1032(.A(G50), .B(new_n1220), .C1(new_n311), .C2(new_n276), .ZN(new_n1233));
  XOR2_X1   g1033(.A(new_n1233), .B(KEYINPUT115), .Z(new_n1234));
  NAND4_X1  g1034(.A1(new_n1223), .A2(new_n1231), .A3(new_n1232), .A4(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1210), .B1(new_n1235), .B2(new_n760), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1208), .B1(new_n1209), .B2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1207), .A2(new_n1237), .ZN(G375));
  XOR2_X1   g1038(.A(new_n1010), .B(KEYINPUT119), .Z(new_n1239));
  NAND2_X1  g1039(.A1(new_n1142), .A2(new_n1239), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1173), .A2(new_n1135), .ZN(new_n1241));
  OR2_X1    g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT120), .ZN(new_n1243));
  OR2_X1    g1043(.A1(new_n1134), .A2(new_n913), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n1243), .B(new_n747), .C1(new_n1244), .C2(new_n1132), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n749), .B1(G68), .B2(new_n829), .ZN(new_n1246));
  XOR2_X1   g1046(.A(new_n1246), .B(KEYINPUT121), .Z(new_n1247));
  NOR2_X1   g1047(.A1(new_n914), .A2(new_n758), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n276), .B(new_n1226), .C1(G50), .C2(new_n845), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n766), .A2(G159), .B1(G128), .B2(new_n781), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(G132), .A2(new_n774), .B1(new_n784), .B2(G137), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(G150), .A2(new_n787), .B1(new_n788), .B2(new_n1158), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1249), .A2(new_n1250), .A3(new_n1251), .A4(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n774), .A2(G294), .ZN(new_n1254));
  OAI221_X1 g1054(.A(new_n1254), .B1(new_n799), .B2(new_n415), .C1(new_n552), .C2(new_n959), .ZN(new_n1255));
  XNOR2_X1  g1055(.A(new_n1255), .B(KEYINPUT122), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n784), .A2(G283), .B1(new_n410), .B2(new_n845), .ZN(new_n1257));
  XNOR2_X1  g1057(.A(new_n1257), .B(KEYINPUT123), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n766), .A2(G97), .B1(G303), .B2(new_n781), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1258), .A2(new_n276), .A3(new_n961), .A4(new_n1259), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1253), .B1(new_n1256), .B2(new_n1260), .ZN(new_n1261));
  AOI211_X1 g1061(.A(new_n1247), .B(new_n1248), .C1(new_n760), .C2(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(KEYINPUT120), .B1(new_n1135), .B2(new_n748), .ZN(new_n1263));
  NOR3_X1   g1063(.A1(new_n1245), .A2(new_n1262), .A3(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1242), .A2(new_n1264), .ZN(G381));
  OR2_X1    g1065(.A1(G393), .A2(G396), .ZN(new_n1266));
  NOR4_X1   g1066(.A1(new_n1266), .A2(G384), .A3(new_n1167), .A4(G381), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1073), .A2(KEYINPUT103), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n999), .A2(new_n743), .A3(new_n1000), .A4(new_n1005), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1269), .B1(new_n1007), .B2(new_n705), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1002), .B1(new_n1268), .B2(new_n1270), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n747), .B1(new_n1271), .B2(new_n1010), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1030), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(new_n1272), .A2(new_n1273), .B1(new_n979), .B2(new_n972), .ZN(new_n1274));
  INV_X1    g1074(.A(G375), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1267), .A2(new_n1274), .A3(new_n1104), .A4(new_n1275), .ZN(G407));
  INV_X1    g1076(.A(new_n1167), .ZN(new_n1277));
  INV_X1    g1077(.A(G213), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1278), .A2(G343), .ZN(new_n1279));
  XOR2_X1   g1079(.A(new_n1279), .B(KEYINPUT124), .Z(new_n1280));
  NAND3_X1  g1080(.A1(new_n1275), .A2(new_n1277), .A3(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(G407), .A2(G213), .A3(new_n1281), .ZN(G409));
  OAI21_X1  g1082(.A(G387), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1075), .A2(new_n1100), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT110), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1274), .A2(new_n1286), .A3(new_n1101), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT125), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1283), .A2(new_n1287), .A3(new_n1288), .ZN(new_n1289));
  XNOR2_X1  g1089(.A(G393), .B(new_n812), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1290), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1292), .A2(new_n1283), .A3(new_n1287), .A4(new_n1288), .ZN(new_n1293));
  AND2_X1   g1093(.A1(new_n1291), .A2(new_n1293), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1207), .A2(new_n1168), .A3(new_n1170), .A4(new_n1237), .ZN(new_n1295));
  AND2_X1   g1095(.A1(new_n1206), .A2(new_n1239), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1200), .A2(new_n748), .A3(new_n1201), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1209), .A2(new_n1236), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1277), .B1(new_n1296), .B2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1295), .A2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1279), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1241), .B1(KEYINPUT60), .B2(new_n1142), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1172), .A2(KEYINPUT60), .A3(new_n1244), .A4(new_n1132), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n708), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1264), .B1(new_n1304), .B2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(new_n855), .ZN(new_n1308));
  OAI211_X1 g1108(.A(G384), .B(new_n1264), .C1(new_n1304), .C2(new_n1306), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1280), .A2(G2897), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1279), .A2(G2897), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1312), .B1(new_n1310), .B2(new_n1313), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1280), .B1(new_n1295), .B2(new_n1300), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT63), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1310), .A2(new_n1316), .ZN(new_n1317));
  AOI22_X1  g1117(.A1(new_n1303), .A2(new_n1314), .B1(new_n1315), .B2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT61), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1310), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1301), .A2(new_n1302), .A3(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1321), .A2(new_n1316), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1294), .A2(new_n1318), .A3(new_n1319), .A4(new_n1322), .ZN(new_n1323));
  XOR2_X1   g1123(.A(KEYINPUT126), .B(KEYINPUT61), .Z(new_n1324));
  INV_X1    g1124(.A(new_n1314), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1324), .B1(new_n1325), .B2(new_n1315), .ZN(new_n1326));
  AOI211_X1 g1126(.A(new_n1279), .B(new_n1310), .C1(new_n1295), .C2(new_n1300), .ZN(new_n1327));
  OAI21_X1  g1127(.A(KEYINPUT127), .B1(new_n1327), .B2(KEYINPUT62), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT127), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT62), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1321), .A2(new_n1329), .A3(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1328), .A2(new_n1331), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1315), .A2(KEYINPUT62), .A3(new_n1320), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1326), .B1(new_n1332), .B2(new_n1333), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1323), .B1(new_n1334), .B2(new_n1294), .ZN(G405));
  NAND2_X1  g1135(.A1(G375), .A2(new_n1277), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1336), .A2(new_n1295), .ZN(new_n1337));
  AND3_X1   g1137(.A1(new_n1291), .A2(new_n1293), .A3(new_n1337), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1337), .B1(new_n1291), .B2(new_n1293), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1310), .B1(new_n1338), .B2(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1291), .A2(new_n1293), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1337), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1341), .A2(new_n1342), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1291), .A2(new_n1293), .A3(new_n1337), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1343), .A2(new_n1320), .A3(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1340), .A2(new_n1345), .ZN(G402));
endmodule


