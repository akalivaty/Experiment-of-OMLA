

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587;

  XOR2_X2 U322 ( .A(n577), .B(KEYINPUT41), .Z(n502) );
  XNOR2_X1 U323 ( .A(n410), .B(KEYINPUT37), .ZN(n411) );
  XOR2_X1 U324 ( .A(n309), .B(n308), .Z(n558) );
  XOR2_X1 U325 ( .A(G134GAT), .B(G106GAT), .Z(n290) );
  XOR2_X1 U326 ( .A(n327), .B(n422), .Z(n291) );
  XOR2_X1 U327 ( .A(n470), .B(n469), .Z(n292) );
  XNOR2_X1 U328 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U329 ( .A(KEYINPUT54), .B(KEYINPUT122), .ZN(n469) );
  XNOR2_X1 U330 ( .A(n334), .B(n333), .ZN(n336) );
  XNOR2_X1 U331 ( .A(n297), .B(n290), .ZN(n302) );
  XNOR2_X1 U332 ( .A(n353), .B(n341), .ZN(n342) );
  XNOR2_X1 U333 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U334 ( .A(n343), .B(n342), .ZN(n358) );
  XOR2_X1 U335 ( .A(KEYINPUT36), .B(n558), .Z(n585) );
  XNOR2_X1 U336 ( .A(n412), .B(n411), .ZN(n516) );
  XOR2_X1 U337 ( .A(n475), .B(KEYINPUT124), .Z(n567) );
  XNOR2_X1 U338 ( .A(n476), .B(G190GAT), .ZN(n477) );
  XNOR2_X1 U339 ( .A(n454), .B(G50GAT), .ZN(n455) );
  XNOR2_X1 U340 ( .A(n478), .B(n477), .ZN(G1351GAT) );
  XNOR2_X1 U341 ( .A(n456), .B(n455), .ZN(G1331GAT) );
  XOR2_X1 U342 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n294) );
  XNOR2_X1 U343 ( .A(G92GAT), .B(KEYINPUT73), .ZN(n293) );
  XNOR2_X1 U344 ( .A(n294), .B(n293), .ZN(n304) );
  XOR2_X1 U345 ( .A(G99GAT), .B(G85GAT), .Z(n414) );
  XOR2_X1 U346 ( .A(KEYINPUT72), .B(n414), .Z(n296) );
  XOR2_X1 U347 ( .A(G50GAT), .B(G162GAT), .Z(n327) );
  XNOR2_X1 U348 ( .A(G218GAT), .B(n327), .ZN(n295) );
  XNOR2_X1 U349 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U350 ( .A(G36GAT), .B(G190GAT), .ZN(n298) );
  XNOR2_X1 U351 ( .A(n298), .B(KEYINPUT74), .ZN(n347) );
  XOR2_X1 U352 ( .A(n347), .B(KEYINPUT11), .Z(n300) );
  NAND2_X1 U353 ( .A1(G232GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U354 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U355 ( .A(n304), .B(n303), .ZN(n309) );
  XOR2_X1 U356 ( .A(KEYINPUT68), .B(KEYINPUT8), .Z(n306) );
  XNOR2_X1 U357 ( .A(G43GAT), .B(G29GAT), .ZN(n305) );
  XNOR2_X1 U358 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U359 ( .A(KEYINPUT7), .B(n307), .ZN(n445) );
  INV_X1 U360 ( .A(n445), .ZN(n308) );
  XOR2_X1 U361 ( .A(G127GAT), .B(KEYINPUT0), .Z(n311) );
  XNOR2_X1 U362 ( .A(G113GAT), .B(G134GAT), .ZN(n310) );
  XNOR2_X1 U363 ( .A(n311), .B(n310), .ZN(n366) );
  XOR2_X1 U364 ( .A(G120GAT), .B(G71GAT), .Z(n430) );
  XOR2_X1 U365 ( .A(n366), .B(n430), .Z(n313) );
  NAND2_X1 U366 ( .A1(G227GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U367 ( .A(n313), .B(n312), .ZN(n317) );
  XOR2_X1 U368 ( .A(G176GAT), .B(G183GAT), .Z(n315) );
  XNOR2_X1 U369 ( .A(KEYINPUT20), .B(KEYINPUT79), .ZN(n314) );
  XNOR2_X1 U370 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U371 ( .A(n317), .B(n316), .Z(n325) );
  XOR2_X1 U372 ( .A(KEYINPUT17), .B(KEYINPUT80), .Z(n319) );
  XNOR2_X1 U373 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n318) );
  XNOR2_X1 U374 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U375 ( .A(G169GAT), .B(n320), .Z(n357) );
  XOR2_X1 U376 ( .A(G190GAT), .B(G99GAT), .Z(n322) );
  XNOR2_X1 U377 ( .A(G43GAT), .B(G15GAT), .ZN(n321) );
  XNOR2_X1 U378 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U379 ( .A(n357), .B(n323), .ZN(n324) );
  XOR2_X1 U380 ( .A(n325), .B(n324), .Z(n531) );
  INV_X1 U381 ( .A(n531), .ZN(n521) );
  XNOR2_X1 U382 ( .A(G106GAT), .B(G78GAT), .ZN(n326) );
  XNOR2_X1 U383 ( .A(n326), .B(G148GAT), .ZN(n422) );
  NAND2_X1 U384 ( .A1(G228GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U385 ( .A(n291), .B(n328), .ZN(n334) );
  XOR2_X1 U386 ( .A(KEYINPUT82), .B(KEYINPUT3), .Z(n330) );
  XNOR2_X1 U387 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n329) );
  XNOR2_X1 U388 ( .A(n330), .B(n329), .ZN(n377) );
  XNOR2_X1 U389 ( .A(n377), .B(KEYINPUT23), .ZN(n332) );
  INV_X1 U390 ( .A(KEYINPUT24), .ZN(n331) );
  INV_X1 U391 ( .A(KEYINPUT83), .ZN(n335) );
  XNOR2_X1 U392 ( .A(n336), .B(n335), .ZN(n343) );
  XNOR2_X1 U393 ( .A(G211GAT), .B(G218GAT), .ZN(n337) );
  XNOR2_X1 U394 ( .A(n337), .B(KEYINPUT21), .ZN(n338) );
  XOR2_X1 U395 ( .A(n338), .B(KEYINPUT81), .Z(n340) );
  XNOR2_X1 U396 ( .A(G197GAT), .B(G204GAT), .ZN(n339) );
  XNOR2_X1 U397 ( .A(n340), .B(n339), .ZN(n353) );
  XOR2_X1 U398 ( .A(G22GAT), .B(G155GAT), .Z(n399) );
  XNOR2_X1 U399 ( .A(n399), .B(KEYINPUT22), .ZN(n341) );
  NOR2_X1 U400 ( .A1(n521), .A2(n358), .ZN(n345) );
  INV_X1 U401 ( .A(KEYINPUT26), .ZN(n344) );
  XNOR2_X1 U402 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U403 ( .A(KEYINPUT91), .B(n346), .Z(n549) );
  INV_X1 U404 ( .A(n549), .ZN(n572) );
  XOR2_X1 U405 ( .A(KEYINPUT89), .B(n347), .Z(n349) );
  NAND2_X1 U406 ( .A1(G226GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U407 ( .A(n349), .B(n348), .ZN(n351) );
  XNOR2_X1 U408 ( .A(G176GAT), .B(G92GAT), .ZN(n350) );
  XNOR2_X1 U409 ( .A(n350), .B(G64GAT), .ZN(n413) );
  XOR2_X1 U410 ( .A(n351), .B(n413), .Z(n355) );
  XNOR2_X1 U411 ( .A(G8GAT), .B(G183GAT), .ZN(n352) );
  XNOR2_X1 U412 ( .A(n352), .B(KEYINPUT75), .ZN(n396) );
  XNOR2_X1 U413 ( .A(n353), .B(n396), .ZN(n354) );
  XNOR2_X1 U414 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U415 ( .A(n357), .B(n356), .ZN(n519) );
  XNOR2_X1 U416 ( .A(KEYINPUT27), .B(n519), .ZN(n387) );
  NAND2_X1 U417 ( .A1(n572), .A2(n387), .ZN(n362) );
  NAND2_X1 U418 ( .A1(n521), .A2(n519), .ZN(n359) );
  NAND2_X1 U419 ( .A1(n358), .A2(n359), .ZN(n360) );
  XOR2_X1 U420 ( .A(KEYINPUT25), .B(n360), .Z(n361) );
  NAND2_X1 U421 ( .A1(n362), .A2(n361), .ZN(n363) );
  XNOR2_X1 U422 ( .A(n363), .B(KEYINPUT92), .ZN(n385) );
  XOR2_X1 U423 ( .A(KEYINPUT5), .B(KEYINPUT88), .Z(n365) );
  XNOR2_X1 U424 ( .A(KEYINPUT87), .B(KEYINPUT85), .ZN(n364) );
  XNOR2_X1 U425 ( .A(n365), .B(n364), .ZN(n370) );
  XOR2_X1 U426 ( .A(n366), .B(KEYINPUT4), .Z(n368) );
  NAND2_X1 U427 ( .A1(G225GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U428 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U429 ( .A(n370), .B(n369), .ZN(n384) );
  XOR2_X1 U430 ( .A(KEYINPUT84), .B(KEYINPUT1), .Z(n372) );
  XNOR2_X1 U431 ( .A(G155GAT), .B(G148GAT), .ZN(n371) );
  XNOR2_X1 U432 ( .A(n372), .B(n371), .ZN(n376) );
  XOR2_X1 U433 ( .A(KEYINPUT86), .B(G57GAT), .Z(n374) );
  XNOR2_X1 U434 ( .A(G1GAT), .B(KEYINPUT6), .ZN(n373) );
  XNOR2_X1 U435 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U436 ( .A(n376), .B(n375), .Z(n382) );
  XOR2_X1 U437 ( .A(G85GAT), .B(G162GAT), .Z(n379) );
  XNOR2_X1 U438 ( .A(G29GAT), .B(n377), .ZN(n378) );
  XNOR2_X1 U439 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U440 ( .A(G120GAT), .B(n380), .ZN(n381) );
  XNOR2_X1 U441 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U442 ( .A(n384), .B(n383), .ZN(n517) );
  INV_X1 U443 ( .A(n517), .ZN(n571) );
  NAND2_X1 U444 ( .A1(n385), .A2(n571), .ZN(n391) );
  XNOR2_X1 U445 ( .A(KEYINPUT64), .B(KEYINPUT28), .ZN(n386) );
  XOR2_X1 U446 ( .A(n386), .B(n358), .Z(n525) );
  INV_X1 U447 ( .A(n525), .ZN(n533) );
  NAND2_X1 U448 ( .A1(n387), .A2(n517), .ZN(n388) );
  XOR2_X1 U449 ( .A(KEYINPUT90), .B(n388), .Z(n529) );
  NAND2_X1 U450 ( .A1(n533), .A2(n529), .ZN(n389) );
  OR2_X1 U451 ( .A1(n521), .A2(n389), .ZN(n390) );
  AND2_X1 U452 ( .A1(n391), .A2(n390), .ZN(n392) );
  XOR2_X1 U453 ( .A(n392), .B(KEYINPUT93), .Z(n483) );
  NOR2_X1 U454 ( .A1(n585), .A2(n483), .ZN(n409) );
  XOR2_X1 U455 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n398) );
  XOR2_X1 U456 ( .A(KEYINPUT14), .B(KEYINPUT76), .Z(n394) );
  XNOR2_X1 U457 ( .A(G64GAT), .B(KEYINPUT77), .ZN(n393) );
  XNOR2_X1 U458 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U459 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U460 ( .A(n398), .B(n397), .ZN(n403) );
  XOR2_X1 U461 ( .A(G57GAT), .B(KEYINPUT13), .Z(n429) );
  XOR2_X1 U462 ( .A(n429), .B(n399), .Z(n401) );
  NAND2_X1 U463 ( .A1(G231GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U464 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U465 ( .A(n403), .B(n402), .Z(n408) );
  XOR2_X1 U466 ( .A(G15GAT), .B(G1GAT), .Z(n438) );
  XOR2_X1 U467 ( .A(G78GAT), .B(G211GAT), .Z(n405) );
  XNOR2_X1 U468 ( .A(G127GAT), .B(G71GAT), .ZN(n404) );
  XNOR2_X1 U469 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U470 ( .A(n438), .B(n406), .ZN(n407) );
  XOR2_X1 U471 ( .A(n408), .B(n407), .Z(n582) );
  INV_X1 U472 ( .A(n582), .ZN(n479) );
  NAND2_X1 U473 ( .A1(n409), .A2(n479), .ZN(n412) );
  XNOR2_X1 U474 ( .A(KEYINPUT97), .B(KEYINPUT98), .ZN(n410) );
  XNOR2_X1 U475 ( .A(n414), .B(n413), .ZN(n415) );
  AND2_X1 U476 ( .A1(G230GAT), .A2(G233GAT), .ZN(n416) );
  NAND2_X1 U477 ( .A1(n415), .A2(n416), .ZN(n420) );
  INV_X1 U478 ( .A(n415), .ZN(n418) );
  INV_X1 U479 ( .A(n416), .ZN(n417) );
  NAND2_X1 U480 ( .A1(n418), .A2(n417), .ZN(n419) );
  NAND2_X1 U481 ( .A1(n420), .A2(n419), .ZN(n421) );
  XOR2_X1 U482 ( .A(n421), .B(KEYINPUT31), .Z(n424) );
  XNOR2_X1 U483 ( .A(n422), .B(KEYINPUT33), .ZN(n423) );
  XNOR2_X1 U484 ( .A(n424), .B(n423), .ZN(n428) );
  XOR2_X1 U485 ( .A(KEYINPUT70), .B(KEYINPUT32), .Z(n426) );
  XNOR2_X1 U486 ( .A(G204GAT), .B(KEYINPUT69), .ZN(n425) );
  XOR2_X1 U487 ( .A(n426), .B(n425), .Z(n427) );
  XNOR2_X1 U488 ( .A(n428), .B(n427), .ZN(n432) );
  XNOR2_X1 U489 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U490 ( .A(n432), .B(n431), .ZN(n577) );
  XOR2_X1 U491 ( .A(KEYINPUT67), .B(KEYINPUT65), .Z(n434) );
  XNOR2_X1 U492 ( .A(G141GAT), .B(G8GAT), .ZN(n433) );
  XNOR2_X1 U493 ( .A(n434), .B(n433), .ZN(n449) );
  XOR2_X1 U494 ( .A(G22GAT), .B(G197GAT), .Z(n436) );
  XNOR2_X1 U495 ( .A(G50GAT), .B(G36GAT), .ZN(n435) );
  XNOR2_X1 U496 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U497 ( .A(n437), .B(G113GAT), .Z(n440) );
  XNOR2_X1 U498 ( .A(G169GAT), .B(n438), .ZN(n439) );
  XNOR2_X1 U499 ( .A(n440), .B(n439), .ZN(n444) );
  XOR2_X1 U500 ( .A(KEYINPUT29), .B(KEYINPUT66), .Z(n442) );
  NAND2_X1 U501 ( .A1(G229GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U502 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U503 ( .A(n444), .B(n443), .Z(n447) );
  XOR2_X1 U504 ( .A(n445), .B(KEYINPUT30), .Z(n446) );
  XNOR2_X1 U505 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U506 ( .A(n449), .B(n448), .ZN(n574) );
  NOR2_X1 U507 ( .A1(n577), .A2(n574), .ZN(n450) );
  XNOR2_X1 U508 ( .A(KEYINPUT71), .B(n450), .ZN(n485) );
  NOR2_X1 U509 ( .A1(n516), .A2(n485), .ZN(n453) );
  XNOR2_X1 U510 ( .A(KEYINPUT99), .B(KEYINPUT100), .ZN(n451) );
  XOR2_X1 U511 ( .A(n451), .B(KEYINPUT38), .Z(n452) );
  XNOR2_X1 U512 ( .A(n453), .B(n452), .ZN(n498) );
  NAND2_X1 U513 ( .A1(n498), .A2(n525), .ZN(n456) );
  XOR2_X1 U514 ( .A(KEYINPUT103), .B(KEYINPUT102), .Z(n454) );
  XOR2_X1 U515 ( .A(KEYINPUT123), .B(KEYINPUT55), .Z(n473) );
  AND2_X1 U516 ( .A1(n571), .A2(n358), .ZN(n471) );
  NOR2_X1 U517 ( .A1(n479), .A2(n585), .ZN(n458) );
  XNOR2_X1 U518 ( .A(KEYINPUT45), .B(KEYINPUT110), .ZN(n457) );
  XNOR2_X1 U519 ( .A(n458), .B(n457), .ZN(n460) );
  INV_X1 U520 ( .A(n574), .ZN(n562) );
  NOR2_X1 U521 ( .A1(n562), .A2(n577), .ZN(n459) );
  NAND2_X1 U522 ( .A1(n460), .A2(n459), .ZN(n466) );
  NAND2_X1 U523 ( .A1(n562), .A2(n502), .ZN(n461) );
  XNOR2_X1 U524 ( .A(n461), .B(KEYINPUT46), .ZN(n463) );
  NOR2_X1 U525 ( .A1(n558), .A2(n582), .ZN(n462) );
  AND2_X1 U526 ( .A1(n463), .A2(n462), .ZN(n464) );
  XNOR2_X1 U527 ( .A(KEYINPUT47), .B(n464), .ZN(n465) );
  NAND2_X1 U528 ( .A1(n466), .A2(n465), .ZN(n468) );
  XOR2_X1 U529 ( .A(KEYINPUT48), .B(KEYINPUT111), .Z(n467) );
  XNOR2_X1 U530 ( .A(n468), .B(n467), .ZN(n530) );
  NAND2_X1 U531 ( .A1(n519), .A2(n530), .ZN(n470) );
  NAND2_X1 U532 ( .A1(n471), .A2(n292), .ZN(n472) );
  XNOR2_X1 U533 ( .A(n473), .B(n472), .ZN(n474) );
  NAND2_X1 U534 ( .A1(n474), .A2(n521), .ZN(n475) );
  NAND2_X1 U535 ( .A1(n567), .A2(n558), .ZN(n478) );
  XOR2_X1 U536 ( .A(KEYINPUT58), .B(KEYINPUT125), .Z(n476) );
  XNOR2_X1 U537 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n487) );
  OR2_X1 U538 ( .A1(n479), .A2(n558), .ZN(n480) );
  XNOR2_X1 U539 ( .A(n480), .B(KEYINPUT78), .ZN(n481) );
  XNOR2_X1 U540 ( .A(n481), .B(KEYINPUT16), .ZN(n482) );
  NOR2_X1 U541 ( .A1(n483), .A2(n482), .ZN(n484) );
  XOR2_X1 U542 ( .A(KEYINPUT94), .B(n484), .Z(n503) );
  NOR2_X1 U543 ( .A1(n503), .A2(n485), .ZN(n493) );
  NAND2_X1 U544 ( .A1(n517), .A2(n493), .ZN(n486) );
  XNOR2_X1 U545 ( .A(n487), .B(n486), .ZN(G1324GAT) );
  NAND2_X1 U546 ( .A1(n519), .A2(n493), .ZN(n488) );
  XNOR2_X1 U547 ( .A(n488), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U548 ( .A(KEYINPUT96), .B(KEYINPUT35), .Z(n490) );
  NAND2_X1 U549 ( .A1(n493), .A2(n521), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n490), .B(n489), .ZN(n492) );
  XOR2_X1 U551 ( .A(G15GAT), .B(KEYINPUT95), .Z(n491) );
  XNOR2_X1 U552 ( .A(n492), .B(n491), .ZN(G1326GAT) );
  NAND2_X1 U553 ( .A1(n493), .A2(n525), .ZN(n494) );
  XNOR2_X1 U554 ( .A(n494), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U555 ( .A(G29GAT), .B(KEYINPUT39), .Z(n496) );
  NAND2_X1 U556 ( .A1(n498), .A2(n517), .ZN(n495) );
  XNOR2_X1 U557 ( .A(n496), .B(n495), .ZN(G1328GAT) );
  NAND2_X1 U558 ( .A1(n519), .A2(n498), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n497), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U560 ( .A1(n498), .A2(n521), .ZN(n500) );
  XOR2_X1 U561 ( .A(KEYINPUT101), .B(KEYINPUT40), .Z(n499) );
  XNOR2_X1 U562 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U563 ( .A(n501), .B(G43GAT), .ZN(G1330GAT) );
  XNOR2_X1 U564 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n505) );
  NAND2_X1 U565 ( .A1(n502), .A2(n574), .ZN(n515) );
  NOR2_X1 U566 ( .A1(n503), .A2(n515), .ZN(n510) );
  NAND2_X1 U567 ( .A1(n517), .A2(n510), .ZN(n504) );
  XNOR2_X1 U568 ( .A(n505), .B(n504), .ZN(G1332GAT) );
  NAND2_X1 U569 ( .A1(n519), .A2(n510), .ZN(n506) );
  XNOR2_X1 U570 ( .A(n506), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U571 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n508) );
  NAND2_X1 U572 ( .A1(n510), .A2(n521), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U574 ( .A(G71GAT), .B(n509), .ZN(G1334GAT) );
  XOR2_X1 U575 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n512) );
  NAND2_X1 U576 ( .A1(n510), .A2(n525), .ZN(n511) );
  XNOR2_X1 U577 ( .A(n512), .B(n511), .ZN(n514) );
  XOR2_X1 U578 ( .A(G78GAT), .B(KEYINPUT106), .Z(n513) );
  XNOR2_X1 U579 ( .A(n514), .B(n513), .ZN(G1335GAT) );
  NOR2_X1 U580 ( .A1(n516), .A2(n515), .ZN(n526) );
  NAND2_X1 U581 ( .A1(n517), .A2(n526), .ZN(n518) );
  XNOR2_X1 U582 ( .A(G85GAT), .B(n518), .ZN(G1336GAT) );
  NAND2_X1 U583 ( .A1(n519), .A2(n526), .ZN(n520) );
  XNOR2_X1 U584 ( .A(n520), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U585 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n523) );
  NAND2_X1 U586 ( .A1(n526), .A2(n521), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U588 ( .A(G99GAT), .B(n524), .ZN(G1338GAT) );
  NAND2_X1 U589 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U590 ( .A(n527), .B(KEYINPUT44), .ZN(n528) );
  XNOR2_X1 U591 ( .A(G106GAT), .B(n528), .ZN(G1339GAT) );
  NAND2_X1 U592 ( .A1(n530), .A2(n529), .ZN(n548) );
  NOR2_X1 U593 ( .A1(n531), .A2(n548), .ZN(n532) );
  XNOR2_X1 U594 ( .A(KEYINPUT112), .B(n532), .ZN(n534) );
  NAND2_X1 U595 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U596 ( .A(n535), .B(KEYINPUT113), .ZN(n544) );
  NAND2_X1 U597 ( .A1(n544), .A2(n562), .ZN(n536) );
  XNOR2_X1 U598 ( .A(n536), .B(KEYINPUT114), .ZN(n537) );
  XNOR2_X1 U599 ( .A(G113GAT), .B(n537), .ZN(G1340GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n539) );
  NAND2_X1 U601 ( .A1(n544), .A2(n502), .ZN(n538) );
  XNOR2_X1 U602 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U603 ( .A(G120GAT), .B(n540), .Z(G1341GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n542) );
  NAND2_X1 U605 ( .A1(n544), .A2(n582), .ZN(n541) );
  XNOR2_X1 U606 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U607 ( .A(G127GAT), .B(n543), .Z(G1342GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n546) );
  NAND2_X1 U609 ( .A1(n544), .A2(n558), .ZN(n545) );
  XNOR2_X1 U610 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U611 ( .A(G134GAT), .B(n547), .Z(G1343GAT) );
  XNOR2_X1 U612 ( .A(G141GAT), .B(KEYINPUT118), .ZN(n551) );
  NOR2_X1 U613 ( .A1(n549), .A2(n548), .ZN(n559) );
  NAND2_X1 U614 ( .A1(n562), .A2(n559), .ZN(n550) );
  XNOR2_X1 U615 ( .A(n551), .B(n550), .ZN(G1344GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT52), .B(KEYINPUT119), .Z(n553) );
  NAND2_X1 U617 ( .A1(n559), .A2(n502), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n553), .B(n552), .ZN(n555) );
  XOR2_X1 U619 ( .A(G148GAT), .B(KEYINPUT53), .Z(n554) );
  XNOR2_X1 U620 ( .A(n555), .B(n554), .ZN(G1345GAT) );
  NAND2_X1 U621 ( .A1(n582), .A2(n559), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n556), .B(KEYINPUT120), .ZN(n557) );
  XNOR2_X1 U623 ( .A(G155GAT), .B(n557), .ZN(G1346GAT) );
  XOR2_X1 U624 ( .A(G162GAT), .B(KEYINPUT121), .Z(n561) );
  NAND2_X1 U625 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n561), .B(n560), .ZN(G1347GAT) );
  NAND2_X1 U627 ( .A1(n562), .A2(n567), .ZN(n563) );
  XNOR2_X1 U628 ( .A(G169GAT), .B(n563), .ZN(G1348GAT) );
  NAND2_X1 U629 ( .A1(n567), .A2(n502), .ZN(n565) );
  XOR2_X1 U630 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U632 ( .A(G176GAT), .B(n566), .ZN(G1349GAT) );
  NAND2_X1 U633 ( .A1(n567), .A2(n582), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n568), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n570) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n570), .B(n569), .ZN(n576) );
  AND2_X1 U638 ( .A1(n571), .A2(n292), .ZN(n573) );
  NAND2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n584) );
  NOR2_X1 U640 ( .A1(n574), .A2(n584), .ZN(n575) );
  XOR2_X1 U641 ( .A(n576), .B(n575), .Z(G1352GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT61), .B(KEYINPUT127), .Z(n579) );
  INV_X1 U643 ( .A(n584), .ZN(n581) );
  NAND2_X1 U644 ( .A1(n581), .A2(n577), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(n580) );
  XOR2_X1 U646 ( .A(G204GAT), .B(n580), .Z(G1353GAT) );
  NAND2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n583), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U650 ( .A(KEYINPUT62), .B(n586), .Z(n587) );
  XNOR2_X1 U651 ( .A(G218GAT), .B(n587), .ZN(G1355GAT) );
endmodule

