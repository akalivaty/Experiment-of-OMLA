

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U550 ( .A1(n675), .A2(n748), .ZN(n714) );
  NOR2_X2 U551 ( .A1(G2105), .A2(n523), .ZN(n882) );
  XNOR2_X1 U552 ( .A(n707), .B(KEYINPUT90), .ZN(n782) );
  XOR2_X1 U553 ( .A(G543), .B(KEYINPUT0), .Z(n515) );
  XOR2_X1 U554 ( .A(KEYINPUT31), .B(n721), .Z(n516) );
  OR2_X1 U555 ( .A1(n938), .A2(n686), .ZN(n687) );
  NOR2_X1 U556 ( .A1(n720), .A2(n719), .ZN(n721) );
  INV_X1 U557 ( .A(KEYINPUT95), .ZN(n731) );
  XNOR2_X1 U558 ( .A(n732), .B(n731), .ZN(n735) );
  XNOR2_X1 U559 ( .A(KEYINPUT97), .B(KEYINPUT32), .ZN(n728) );
  XNOR2_X1 U560 ( .A(n729), .B(n728), .ZN(n739) );
  NOR2_X1 U561 ( .A1(n739), .A2(n738), .ZN(n792) );
  INV_X1 U562 ( .A(n782), .ZN(n794) );
  INV_X1 U563 ( .A(KEYINPUT17), .ZN(n517) );
  NAND2_X1 U564 ( .A1(n885), .A2(G137), .ZN(n519) );
  NOR2_X1 U565 ( .A1(n538), .A2(n634), .ZN(n643) );
  NOR2_X1 U566 ( .A1(G651), .A2(n634), .ZN(n641) );
  NAND2_X1 U567 ( .A1(n582), .A2(n581), .ZN(n954) );
  NOR2_X1 U568 ( .A1(n528), .A2(n527), .ZN(G160) );
  NOR2_X1 U569 ( .A1(G2104), .A2(G2105), .ZN(n518) );
  XNOR2_X2 U570 ( .A(n518), .B(n517), .ZN(n885) );
  XOR2_X1 U571 ( .A(KEYINPUT65), .B(n519), .Z(n522) );
  INV_X1 U572 ( .A(G2104), .ZN(n523) );
  NAND2_X1 U573 ( .A1(G101), .A2(n882), .ZN(n520) );
  XOR2_X1 U574 ( .A(KEYINPUT23), .B(n520), .Z(n521) );
  NAND2_X1 U575 ( .A1(n522), .A2(n521), .ZN(n528) );
  AND2_X1 U576 ( .A1(n523), .A2(G2105), .ZN(n877) );
  NAND2_X1 U577 ( .A1(G125), .A2(n877), .ZN(n526) );
  NAND2_X1 U578 ( .A1(G2105), .A2(G2104), .ZN(n524) );
  XOR2_X1 U579 ( .A(KEYINPUT64), .B(n524), .Z(n878) );
  NAND2_X1 U580 ( .A1(G113), .A2(n878), .ZN(n525) );
  NAND2_X1 U581 ( .A1(n526), .A2(n525), .ZN(n527) );
  NAND2_X1 U582 ( .A1(G138), .A2(n885), .ZN(n530) );
  NAND2_X1 U583 ( .A1(G102), .A2(n882), .ZN(n529) );
  NAND2_X1 U584 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U585 ( .A(KEYINPUT84), .B(n531), .ZN(n535) );
  NAND2_X1 U586 ( .A1(G126), .A2(n877), .ZN(n533) );
  NAND2_X1 U587 ( .A1(G114), .A2(n878), .ZN(n532) );
  NAND2_X1 U588 ( .A1(n533), .A2(n532), .ZN(n534) );
  NOR2_X1 U589 ( .A1(n535), .A2(n534), .ZN(G164) );
  NOR2_X1 U590 ( .A1(G651), .A2(G543), .ZN(n637) );
  NAND2_X1 U591 ( .A1(G91), .A2(n637), .ZN(n537) );
  INV_X1 U592 ( .A(G651), .ZN(n538) );
  XNOR2_X1 U593 ( .A(KEYINPUT66), .B(n515), .ZN(n634) );
  NAND2_X1 U594 ( .A1(G78), .A2(n643), .ZN(n536) );
  NAND2_X1 U595 ( .A1(n537), .A2(n536), .ZN(n543) );
  NOR2_X1 U596 ( .A1(G543), .A2(n538), .ZN(n539) );
  XOR2_X1 U597 ( .A(KEYINPUT1), .B(n539), .Z(n638) );
  NAND2_X1 U598 ( .A1(G65), .A2(n638), .ZN(n541) );
  NAND2_X1 U599 ( .A1(G53), .A2(n641), .ZN(n540) );
  NAND2_X1 U600 ( .A1(n541), .A2(n540), .ZN(n542) );
  OR2_X1 U601 ( .A1(n543), .A2(n542), .ZN(G299) );
  NAND2_X1 U602 ( .A1(G64), .A2(n638), .ZN(n545) );
  NAND2_X1 U603 ( .A1(G52), .A2(n641), .ZN(n544) );
  NAND2_X1 U604 ( .A1(n545), .A2(n544), .ZN(n550) );
  NAND2_X1 U605 ( .A1(G90), .A2(n637), .ZN(n547) );
  NAND2_X1 U606 ( .A1(G77), .A2(n643), .ZN(n546) );
  NAND2_X1 U607 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U608 ( .A(KEYINPUT9), .B(n548), .Z(n549) );
  NOR2_X1 U609 ( .A1(n550), .A2(n549), .ZN(G171) );
  AND2_X1 U610 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U611 ( .A1(G123), .A2(n877), .ZN(n551) );
  XNOR2_X1 U612 ( .A(n551), .B(KEYINPUT18), .ZN(n558) );
  NAND2_X1 U613 ( .A1(G99), .A2(n882), .ZN(n553) );
  NAND2_X1 U614 ( .A1(G111), .A2(n878), .ZN(n552) );
  NAND2_X1 U615 ( .A1(n553), .A2(n552), .ZN(n556) );
  NAND2_X1 U616 ( .A1(G135), .A2(n885), .ZN(n554) );
  XNOR2_X1 U617 ( .A(KEYINPUT73), .B(n554), .ZN(n555) );
  NOR2_X1 U618 ( .A1(n556), .A2(n555), .ZN(n557) );
  NAND2_X1 U619 ( .A1(n558), .A2(n557), .ZN(n990) );
  XNOR2_X1 U620 ( .A(G2096), .B(n990), .ZN(n559) );
  OR2_X1 U621 ( .A1(G2100), .A2(n559), .ZN(G156) );
  INV_X1 U622 ( .A(G132), .ZN(G219) );
  INV_X1 U623 ( .A(G82), .ZN(G220) );
  INV_X1 U624 ( .A(G57), .ZN(G237) );
  INV_X1 U625 ( .A(G120), .ZN(G236) );
  NAND2_X1 U626 ( .A1(G63), .A2(n638), .ZN(n561) );
  NAND2_X1 U627 ( .A1(G51), .A2(n641), .ZN(n560) );
  NAND2_X1 U628 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U629 ( .A(KEYINPUT6), .B(n562), .ZN(n568) );
  NAND2_X1 U630 ( .A1(n637), .A2(G89), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n563), .B(KEYINPUT4), .ZN(n565) );
  NAND2_X1 U632 ( .A1(G76), .A2(n643), .ZN(n564) );
  NAND2_X1 U633 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U634 ( .A(n566), .B(KEYINPUT5), .Z(n567) );
  NOR2_X1 U635 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U636 ( .A(KEYINPUT7), .B(n569), .Z(n570) );
  XNOR2_X1 U637 ( .A(KEYINPUT70), .B(n570), .ZN(G168) );
  XOR2_X1 U638 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U639 ( .A1(G7), .A2(G661), .ZN(n571) );
  XNOR2_X1 U640 ( .A(n571), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U641 ( .A(G223), .ZN(n819) );
  NAND2_X1 U642 ( .A1(n819), .A2(G567), .ZN(n572) );
  XOR2_X1 U643 ( .A(KEYINPUT11), .B(n572), .Z(G234) );
  NAND2_X1 U644 ( .A1(G68), .A2(n643), .ZN(n575) );
  NAND2_X1 U645 ( .A1(n637), .A2(G81), .ZN(n573) );
  XNOR2_X1 U646 ( .A(n573), .B(KEYINPUT12), .ZN(n574) );
  NAND2_X1 U647 ( .A1(n575), .A2(n574), .ZN(n577) );
  XNOR2_X1 U648 ( .A(KEYINPUT67), .B(KEYINPUT13), .ZN(n576) );
  XNOR2_X1 U649 ( .A(n577), .B(n576), .ZN(n580) );
  NAND2_X1 U650 ( .A1(n638), .A2(G56), .ZN(n578) );
  XOR2_X1 U651 ( .A(KEYINPUT14), .B(n578), .Z(n579) );
  NOR2_X1 U652 ( .A1(n580), .A2(n579), .ZN(n582) );
  NAND2_X1 U653 ( .A1(n641), .A2(G43), .ZN(n581) );
  INV_X1 U654 ( .A(G860), .ZN(n596) );
  OR2_X1 U655 ( .A1(n954), .A2(n596), .ZN(G153) );
  INV_X1 U656 ( .A(G868), .ZN(n648) );
  NOR2_X1 U657 ( .A1(G171), .A2(n648), .ZN(n583) );
  XNOR2_X1 U658 ( .A(n583), .B(KEYINPUT68), .ZN(n592) );
  NAND2_X1 U659 ( .A1(G92), .A2(n637), .ZN(n585) );
  NAND2_X1 U660 ( .A1(G79), .A2(n643), .ZN(n584) );
  NAND2_X1 U661 ( .A1(n585), .A2(n584), .ZN(n589) );
  NAND2_X1 U662 ( .A1(G66), .A2(n638), .ZN(n587) );
  NAND2_X1 U663 ( .A1(G54), .A2(n641), .ZN(n586) );
  NAND2_X1 U664 ( .A1(n587), .A2(n586), .ZN(n588) );
  NOR2_X1 U665 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U666 ( .A(KEYINPUT15), .B(n590), .Z(n938) );
  NOR2_X1 U667 ( .A1(n938), .A2(G868), .ZN(n591) );
  NOR2_X1 U668 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U669 ( .A(KEYINPUT69), .B(n593), .ZN(G284) );
  INV_X1 U670 ( .A(G171), .ZN(G301) );
  NAND2_X1 U671 ( .A1(G868), .A2(G286), .ZN(n595) );
  NAND2_X1 U672 ( .A1(G299), .A2(n648), .ZN(n594) );
  NAND2_X1 U673 ( .A1(n595), .A2(n594), .ZN(G297) );
  NAND2_X1 U674 ( .A1(n596), .A2(G559), .ZN(n597) );
  NAND2_X1 U675 ( .A1(n597), .A2(n938), .ZN(n598) );
  XNOR2_X1 U676 ( .A(n598), .B(KEYINPUT71), .ZN(n599) );
  XOR2_X1 U677 ( .A(KEYINPUT16), .B(n599), .Z(G148) );
  NAND2_X1 U678 ( .A1(n938), .A2(G868), .ZN(n600) );
  NOR2_X1 U679 ( .A1(G559), .A2(n600), .ZN(n601) );
  XNOR2_X1 U680 ( .A(n601), .B(KEYINPUT72), .ZN(n603) );
  NOR2_X1 U681 ( .A1(n954), .A2(G868), .ZN(n602) );
  NOR2_X1 U682 ( .A1(n603), .A2(n602), .ZN(G282) );
  NAND2_X1 U683 ( .A1(G559), .A2(n938), .ZN(n604) );
  XOR2_X1 U684 ( .A(n954), .B(n604), .Z(n657) );
  XOR2_X1 U685 ( .A(n657), .B(KEYINPUT74), .Z(n605) );
  NOR2_X1 U686 ( .A1(G860), .A2(n605), .ZN(n606) );
  XOR2_X1 U687 ( .A(KEYINPUT78), .B(n606), .Z(n616) );
  NAND2_X1 U688 ( .A1(n641), .A2(G55), .ZN(n607) );
  XNOR2_X1 U689 ( .A(n607), .B(KEYINPUT76), .ZN(n609) );
  NAND2_X1 U690 ( .A1(G67), .A2(n638), .ZN(n608) );
  NAND2_X1 U691 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U692 ( .A(KEYINPUT77), .B(n610), .ZN(n615) );
  NAND2_X1 U693 ( .A1(G93), .A2(n637), .ZN(n612) );
  NAND2_X1 U694 ( .A1(G80), .A2(n643), .ZN(n611) );
  NAND2_X1 U695 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U696 ( .A(KEYINPUT75), .B(n613), .ZN(n614) );
  NAND2_X1 U697 ( .A1(n615), .A2(n614), .ZN(n654) );
  XNOR2_X1 U698 ( .A(n616), .B(n654), .ZN(G145) );
  AND2_X1 U699 ( .A1(n638), .A2(G60), .ZN(n620) );
  NAND2_X1 U700 ( .A1(G85), .A2(n637), .ZN(n618) );
  NAND2_X1 U701 ( .A1(G72), .A2(n643), .ZN(n617) );
  NAND2_X1 U702 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U703 ( .A1(n620), .A2(n619), .ZN(n622) );
  NAND2_X1 U704 ( .A1(n641), .A2(G47), .ZN(n621) );
  NAND2_X1 U705 ( .A1(n622), .A2(n621), .ZN(G290) );
  NAND2_X1 U706 ( .A1(G73), .A2(n643), .ZN(n623) );
  XOR2_X1 U707 ( .A(KEYINPUT2), .B(n623), .Z(n628) );
  NAND2_X1 U708 ( .A1(G86), .A2(n637), .ZN(n625) );
  NAND2_X1 U709 ( .A1(G61), .A2(n638), .ZN(n624) );
  NAND2_X1 U710 ( .A1(n625), .A2(n624), .ZN(n626) );
  XOR2_X1 U711 ( .A(KEYINPUT79), .B(n626), .Z(n627) );
  NOR2_X1 U712 ( .A1(n628), .A2(n627), .ZN(n630) );
  NAND2_X1 U713 ( .A1(n641), .A2(G48), .ZN(n629) );
  NAND2_X1 U714 ( .A1(n630), .A2(n629), .ZN(G305) );
  NAND2_X1 U715 ( .A1(G49), .A2(n641), .ZN(n632) );
  NAND2_X1 U716 ( .A1(G74), .A2(G651), .ZN(n631) );
  NAND2_X1 U717 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U718 ( .A1(n638), .A2(n633), .ZN(n636) );
  NAND2_X1 U719 ( .A1(G87), .A2(n634), .ZN(n635) );
  NAND2_X1 U720 ( .A1(n636), .A2(n635), .ZN(G288) );
  NAND2_X1 U721 ( .A1(G88), .A2(n637), .ZN(n640) );
  NAND2_X1 U722 ( .A1(G62), .A2(n638), .ZN(n639) );
  NAND2_X1 U723 ( .A1(n640), .A2(n639), .ZN(n647) );
  NAND2_X1 U724 ( .A1(G50), .A2(n641), .ZN(n642) );
  XNOR2_X1 U725 ( .A(n642), .B(KEYINPUT80), .ZN(n645) );
  NAND2_X1 U726 ( .A1(n643), .A2(G75), .ZN(n644) );
  NAND2_X1 U727 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U728 ( .A1(n647), .A2(n646), .ZN(G166) );
  NAND2_X1 U729 ( .A1(n648), .A2(n654), .ZN(n649) );
  XNOR2_X1 U730 ( .A(n649), .B(KEYINPUT82), .ZN(n660) );
  XOR2_X1 U731 ( .A(G290), .B(G305), .Z(n650) );
  XNOR2_X1 U732 ( .A(G299), .B(n650), .ZN(n653) );
  XOR2_X1 U733 ( .A(KEYINPUT19), .B(KEYINPUT81), .Z(n651) );
  XNOR2_X1 U734 ( .A(G288), .B(n651), .ZN(n652) );
  XOR2_X1 U735 ( .A(n653), .B(n652), .Z(n656) );
  XOR2_X1 U736 ( .A(G166), .B(n654), .Z(n655) );
  XNOR2_X1 U737 ( .A(n656), .B(n655), .ZN(n892) );
  XNOR2_X1 U738 ( .A(n892), .B(n657), .ZN(n658) );
  NAND2_X1 U739 ( .A1(G868), .A2(n658), .ZN(n659) );
  NAND2_X1 U740 ( .A1(n660), .A2(n659), .ZN(G295) );
  NAND2_X1 U741 ( .A1(G2084), .A2(G2078), .ZN(n661) );
  XOR2_X1 U742 ( .A(KEYINPUT20), .B(n661), .Z(n662) );
  NAND2_X1 U743 ( .A1(G2090), .A2(n662), .ZN(n663) );
  XNOR2_X1 U744 ( .A(KEYINPUT21), .B(n663), .ZN(n664) );
  NAND2_X1 U745 ( .A1(n664), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U746 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U747 ( .A1(G236), .A2(G237), .ZN(n665) );
  NAND2_X1 U748 ( .A1(G69), .A2(n665), .ZN(n666) );
  XNOR2_X1 U749 ( .A(KEYINPUT83), .B(n666), .ZN(n667) );
  NAND2_X1 U750 ( .A1(n667), .A2(G108), .ZN(n826) );
  NAND2_X1 U751 ( .A1(G567), .A2(n826), .ZN(n672) );
  NOR2_X1 U752 ( .A1(G220), .A2(G219), .ZN(n668) );
  XOR2_X1 U753 ( .A(KEYINPUT22), .B(n668), .Z(n669) );
  NOR2_X1 U754 ( .A1(G218), .A2(n669), .ZN(n670) );
  NAND2_X1 U755 ( .A1(G96), .A2(n670), .ZN(n827) );
  NAND2_X1 U756 ( .A1(G2106), .A2(n827), .ZN(n671) );
  NAND2_X1 U757 ( .A1(n672), .A2(n671), .ZN(n849) );
  NAND2_X1 U758 ( .A1(G483), .A2(G661), .ZN(n673) );
  NOR2_X1 U759 ( .A1(n849), .A2(n673), .ZN(n825) );
  NAND2_X1 U760 ( .A1(n825), .A2(G36), .ZN(G176) );
  XNOR2_X1 U761 ( .A(KEYINPUT85), .B(G166), .ZN(G303) );
  NAND2_X1 U762 ( .A1(G160), .A2(G40), .ZN(n747) );
  INV_X1 U763 ( .A(n747), .ZN(n675) );
  NOR2_X1 U764 ( .A1(G164), .A2(G1384), .ZN(n748) );
  INV_X1 U765 ( .A(G1996), .ZN(n970) );
  NOR2_X1 U766 ( .A1(n714), .A2(n970), .ZN(n677) );
  INV_X1 U767 ( .A(KEYINPUT26), .ZN(n676) );
  XNOR2_X1 U768 ( .A(n677), .B(n676), .ZN(n680) );
  AND2_X1 U769 ( .A1(n714), .A2(G1341), .ZN(n678) );
  NOR2_X1 U770 ( .A1(n678), .A2(n954), .ZN(n679) );
  AND2_X1 U771 ( .A1(n680), .A2(n679), .ZN(n686) );
  NAND2_X1 U772 ( .A1(n938), .A2(n686), .ZN(n685) );
  NAND2_X1 U773 ( .A1(n714), .A2(G1348), .ZN(n681) );
  XNOR2_X1 U774 ( .A(n681), .B(KEYINPUT92), .ZN(n683) );
  INV_X1 U775 ( .A(n714), .ZN(n702) );
  NAND2_X1 U776 ( .A1(n702), .A2(G2067), .ZN(n682) );
  NAND2_X1 U777 ( .A1(n683), .A2(n682), .ZN(n684) );
  NAND2_X1 U778 ( .A1(n685), .A2(n684), .ZN(n688) );
  NAND2_X1 U779 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U780 ( .A(KEYINPUT93), .B(n689), .ZN(n696) );
  AND2_X1 U781 ( .A1(n702), .A2(G2072), .ZN(n691) );
  XOR2_X1 U782 ( .A(KEYINPUT27), .B(KEYINPUT91), .Z(n690) );
  XNOR2_X1 U783 ( .A(n691), .B(n690), .ZN(n693) );
  NAND2_X1 U784 ( .A1(n714), .A2(G1956), .ZN(n692) );
  NAND2_X1 U785 ( .A1(n693), .A2(n692), .ZN(n697) );
  NOR2_X1 U786 ( .A1(G299), .A2(n697), .ZN(n694) );
  XNOR2_X1 U787 ( .A(n694), .B(KEYINPUT94), .ZN(n695) );
  NOR2_X1 U788 ( .A1(n696), .A2(n695), .ZN(n700) );
  NAND2_X1 U789 ( .A1(G299), .A2(n697), .ZN(n698) );
  XOR2_X1 U790 ( .A(KEYINPUT28), .B(n698), .Z(n699) );
  NOR2_X1 U791 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U792 ( .A(n701), .B(KEYINPUT29), .ZN(n706) );
  OR2_X1 U793 ( .A1(n702), .A2(G1961), .ZN(n704) );
  XNOR2_X1 U794 ( .A(G2078), .B(KEYINPUT25), .ZN(n969) );
  NAND2_X1 U795 ( .A1(n702), .A2(n969), .ZN(n703) );
  NAND2_X1 U796 ( .A1(n704), .A2(n703), .ZN(n718) );
  NAND2_X1 U797 ( .A1(G171), .A2(n718), .ZN(n705) );
  NAND2_X1 U798 ( .A1(n706), .A2(n705), .ZN(n730) );
  INV_X1 U799 ( .A(G8), .ZN(n713) );
  NAND2_X1 U800 ( .A1(n714), .A2(G8), .ZN(n707) );
  NOR2_X1 U801 ( .A1(n782), .A2(G1971), .ZN(n709) );
  NOR2_X1 U802 ( .A1(G2090), .A2(n714), .ZN(n708) );
  NOR2_X1 U803 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U804 ( .A1(n710), .A2(G303), .ZN(n711) );
  XNOR2_X1 U805 ( .A(n711), .B(KEYINPUT96), .ZN(n712) );
  OR2_X1 U806 ( .A1(n713), .A2(n712), .ZN(n723) );
  AND2_X1 U807 ( .A1(n730), .A2(n723), .ZN(n722) );
  NOR2_X1 U808 ( .A1(n782), .A2(G1966), .ZN(n736) );
  NOR2_X1 U809 ( .A1(G2084), .A2(n714), .ZN(n733) );
  NOR2_X1 U810 ( .A1(n736), .A2(n733), .ZN(n715) );
  NAND2_X1 U811 ( .A1(G8), .A2(n715), .ZN(n716) );
  XNOR2_X1 U812 ( .A(n716), .B(KEYINPUT30), .ZN(n717) );
  NOR2_X1 U813 ( .A1(n717), .A2(G168), .ZN(n720) );
  NOR2_X1 U814 ( .A1(G171), .A2(n718), .ZN(n719) );
  NAND2_X1 U815 ( .A1(n722), .A2(n516), .ZN(n727) );
  INV_X1 U816 ( .A(n723), .ZN(n725) );
  AND2_X1 U817 ( .A1(G286), .A2(G8), .ZN(n724) );
  OR2_X1 U818 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U819 ( .A1(n727), .A2(n726), .ZN(n729) );
  NAND2_X1 U820 ( .A1(n516), .A2(n730), .ZN(n732) );
  NAND2_X1 U821 ( .A1(n733), .A2(G8), .ZN(n734) );
  NAND2_X1 U822 ( .A1(n735), .A2(n734), .ZN(n737) );
  NOR2_X1 U823 ( .A1(n737), .A2(n736), .ZN(n738) );
  INV_X1 U824 ( .A(n792), .ZN(n741) );
  NOR2_X1 U825 ( .A1(G1976), .A2(G288), .ZN(n744) );
  NOR2_X1 U826 ( .A1(G1971), .A2(G303), .ZN(n740) );
  NOR2_X1 U827 ( .A1(n744), .A2(n740), .ZN(n943) );
  NAND2_X1 U828 ( .A1(n741), .A2(n943), .ZN(n742) );
  NAND2_X1 U829 ( .A1(G1976), .A2(G288), .ZN(n946) );
  NAND2_X1 U830 ( .A1(n742), .A2(n946), .ZN(n743) );
  XNOR2_X1 U831 ( .A(KEYINPUT98), .B(n743), .ZN(n784) );
  AND2_X1 U832 ( .A1(n744), .A2(KEYINPUT33), .ZN(n745) );
  AND2_X1 U833 ( .A1(n745), .A2(n794), .ZN(n746) );
  XNOR2_X1 U834 ( .A(G1981), .B(G305), .ZN(n958) );
  NOR2_X1 U835 ( .A1(n746), .A2(n958), .ZN(n780) );
  NOR2_X1 U836 ( .A1(n748), .A2(n747), .ZN(n814) );
  NAND2_X1 U837 ( .A1(G140), .A2(n885), .ZN(n750) );
  NAND2_X1 U838 ( .A1(G104), .A2(n882), .ZN(n749) );
  NAND2_X1 U839 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U840 ( .A(KEYINPUT34), .B(n751), .ZN(n756) );
  NAND2_X1 U841 ( .A1(G128), .A2(n877), .ZN(n753) );
  NAND2_X1 U842 ( .A1(G116), .A2(n878), .ZN(n752) );
  NAND2_X1 U843 ( .A1(n753), .A2(n752), .ZN(n754) );
  XOR2_X1 U844 ( .A(KEYINPUT35), .B(n754), .Z(n755) );
  NOR2_X1 U845 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U846 ( .A(KEYINPUT36), .B(n757), .ZN(n858) );
  XNOR2_X1 U847 ( .A(KEYINPUT37), .B(G2067), .ZN(n811) );
  NOR2_X1 U848 ( .A1(n858), .A2(n811), .ZN(n997) );
  NAND2_X1 U849 ( .A1(n814), .A2(n997), .ZN(n809) );
  NAND2_X1 U850 ( .A1(G129), .A2(n877), .ZN(n759) );
  NAND2_X1 U851 ( .A1(G117), .A2(n878), .ZN(n758) );
  NAND2_X1 U852 ( .A1(n759), .A2(n758), .ZN(n763) );
  NAND2_X1 U853 ( .A1(G105), .A2(n882), .ZN(n760) );
  XNOR2_X1 U854 ( .A(n760), .B(KEYINPUT38), .ZN(n761) );
  XNOR2_X1 U855 ( .A(n761), .B(KEYINPUT87), .ZN(n762) );
  NOR2_X1 U856 ( .A1(n763), .A2(n762), .ZN(n765) );
  NAND2_X1 U857 ( .A1(n885), .A2(G141), .ZN(n764) );
  NAND2_X1 U858 ( .A1(n765), .A2(n764), .ZN(n859) );
  NAND2_X1 U859 ( .A1(G1996), .A2(n859), .ZN(n766) );
  XNOR2_X1 U860 ( .A(n766), .B(KEYINPUT88), .ZN(n775) );
  NAND2_X1 U861 ( .A1(G119), .A2(n877), .ZN(n768) );
  NAND2_X1 U862 ( .A1(G107), .A2(n878), .ZN(n767) );
  NAND2_X1 U863 ( .A1(n768), .A2(n767), .ZN(n769) );
  XOR2_X1 U864 ( .A(KEYINPUT86), .B(n769), .Z(n773) );
  NAND2_X1 U865 ( .A1(n885), .A2(G131), .ZN(n771) );
  NAND2_X1 U866 ( .A1(G95), .A2(n882), .ZN(n770) );
  AND2_X1 U867 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U868 ( .A1(n773), .A2(n772), .ZN(n862) );
  NAND2_X1 U869 ( .A1(G1991), .A2(n862), .ZN(n774) );
  NAND2_X1 U870 ( .A1(n775), .A2(n774), .ZN(n998) );
  NAND2_X1 U871 ( .A1(n814), .A2(n998), .ZN(n802) );
  NAND2_X1 U872 ( .A1(n809), .A2(n802), .ZN(n776) );
  XNOR2_X1 U873 ( .A(n776), .B(KEYINPUT89), .ZN(n778) );
  XNOR2_X1 U874 ( .A(G1986), .B(G290), .ZN(n950) );
  NAND2_X1 U875 ( .A1(n814), .A2(n950), .ZN(n777) );
  NAND2_X1 U876 ( .A1(n778), .A2(n777), .ZN(n798) );
  INV_X1 U877 ( .A(n798), .ZN(n779) );
  AND2_X1 U878 ( .A1(n780), .A2(n779), .ZN(n785) );
  INV_X1 U879 ( .A(n785), .ZN(n781) );
  OR2_X1 U880 ( .A1(n782), .A2(n781), .ZN(n783) );
  NOR2_X1 U881 ( .A1(n784), .A2(n783), .ZN(n787) );
  AND2_X1 U882 ( .A1(n785), .A2(KEYINPUT33), .ZN(n786) );
  NOR2_X1 U883 ( .A1(n787), .A2(n786), .ZN(n800) );
  NOR2_X1 U884 ( .A1(G1981), .A2(G305), .ZN(n788) );
  XNOR2_X1 U885 ( .A(n788), .B(KEYINPUT24), .ZN(n789) );
  AND2_X1 U886 ( .A1(n789), .A2(n794), .ZN(n796) );
  INV_X1 U887 ( .A(G2090), .ZN(n992) );
  NAND2_X1 U888 ( .A1(G8), .A2(n992), .ZN(n790) );
  NOR2_X1 U889 ( .A1(n790), .A2(G303), .ZN(n791) );
  NOR2_X1 U890 ( .A1(n792), .A2(n791), .ZN(n793) );
  NOR2_X1 U891 ( .A1(n794), .A2(n793), .ZN(n795) );
  NOR2_X1 U892 ( .A1(n796), .A2(n795), .ZN(n797) );
  OR2_X1 U893 ( .A1(n798), .A2(n797), .ZN(n799) );
  NAND2_X1 U894 ( .A1(n800), .A2(n799), .ZN(n801) );
  XNOR2_X1 U895 ( .A(n801), .B(KEYINPUT99), .ZN(n816) );
  NOR2_X1 U896 ( .A1(G1996), .A2(n859), .ZN(n994) );
  INV_X1 U897 ( .A(n802), .ZN(n806) );
  NOR2_X1 U898 ( .A1(G1986), .A2(G290), .ZN(n803) );
  XNOR2_X1 U899 ( .A(n803), .B(KEYINPUT100), .ZN(n804) );
  NOR2_X1 U900 ( .A1(G1991), .A2(n862), .ZN(n989) );
  NOR2_X1 U901 ( .A1(n804), .A2(n989), .ZN(n805) );
  NOR2_X1 U902 ( .A1(n806), .A2(n805), .ZN(n807) );
  NOR2_X1 U903 ( .A1(n994), .A2(n807), .ZN(n808) );
  XNOR2_X1 U904 ( .A(n808), .B(KEYINPUT39), .ZN(n810) );
  NAND2_X1 U905 ( .A1(n810), .A2(n809), .ZN(n812) );
  NAND2_X1 U906 ( .A1(n858), .A2(n811), .ZN(n999) );
  NAND2_X1 U907 ( .A1(n812), .A2(n999), .ZN(n813) );
  NAND2_X1 U908 ( .A1(n814), .A2(n813), .ZN(n815) );
  NAND2_X1 U909 ( .A1(n816), .A2(n815), .ZN(n818) );
  XOR2_X1 U910 ( .A(KEYINPUT101), .B(KEYINPUT40), .Z(n817) );
  XNOR2_X1 U911 ( .A(n818), .B(n817), .ZN(G329) );
  NAND2_X1 U912 ( .A1(n819), .A2(G2106), .ZN(n820) );
  XOR2_X1 U913 ( .A(KEYINPUT103), .B(n820), .Z(G217) );
  NAND2_X1 U914 ( .A1(G15), .A2(G2), .ZN(n821) );
  XOR2_X1 U915 ( .A(KEYINPUT104), .B(n821), .Z(n822) );
  NAND2_X1 U916 ( .A1(G661), .A2(n822), .ZN(G259) );
  NAND2_X1 U917 ( .A1(G3), .A2(G1), .ZN(n823) );
  XOR2_X1 U918 ( .A(KEYINPUT105), .B(n823), .Z(n824) );
  NAND2_X1 U919 ( .A1(n825), .A2(n824), .ZN(G188) );
  INV_X1 U921 ( .A(G108), .ZN(G238) );
  INV_X1 U922 ( .A(G96), .ZN(G221) );
  NOR2_X1 U923 ( .A1(n827), .A2(n826), .ZN(G325) );
  INV_X1 U924 ( .A(G325), .ZN(G261) );
  XOR2_X1 U925 ( .A(KEYINPUT107), .B(G2090), .Z(n829) );
  XNOR2_X1 U926 ( .A(G2084), .B(G2078), .ZN(n828) );
  XNOR2_X1 U927 ( .A(n829), .B(n828), .ZN(n830) );
  XOR2_X1 U928 ( .A(n830), .B(G2100), .Z(n832) );
  XNOR2_X1 U929 ( .A(G2067), .B(G2072), .ZN(n831) );
  XNOR2_X1 U930 ( .A(n832), .B(n831), .ZN(n836) );
  XOR2_X1 U931 ( .A(G2096), .B(KEYINPUT43), .Z(n834) );
  XNOR2_X1 U932 ( .A(KEYINPUT42), .B(G2678), .ZN(n833) );
  XNOR2_X1 U933 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U934 ( .A(n836), .B(n835), .Z(G227) );
  XOR2_X1 U935 ( .A(G1976), .B(G1971), .Z(n838) );
  XNOR2_X1 U936 ( .A(G1986), .B(G1961), .ZN(n837) );
  XNOR2_X1 U937 ( .A(n838), .B(n837), .ZN(n848) );
  XOR2_X1 U938 ( .A(KEYINPUT110), .B(KEYINPUT41), .Z(n840) );
  XNOR2_X1 U939 ( .A(G1996), .B(G2474), .ZN(n839) );
  XNOR2_X1 U940 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U941 ( .A(G1956), .B(G1966), .Z(n842) );
  XNOR2_X1 U942 ( .A(G1991), .B(G1981), .ZN(n841) );
  XNOR2_X1 U943 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U944 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U945 ( .A(KEYINPUT109), .B(KEYINPUT108), .ZN(n845) );
  XNOR2_X1 U946 ( .A(n846), .B(n845), .ZN(n847) );
  XNOR2_X1 U947 ( .A(n848), .B(n847), .ZN(G229) );
  XOR2_X1 U948 ( .A(KEYINPUT106), .B(n849), .Z(G319) );
  NAND2_X1 U949 ( .A1(G124), .A2(n877), .ZN(n850) );
  XOR2_X1 U950 ( .A(KEYINPUT111), .B(n850), .Z(n851) );
  XNOR2_X1 U951 ( .A(n851), .B(KEYINPUT44), .ZN(n853) );
  NAND2_X1 U952 ( .A1(G100), .A2(n882), .ZN(n852) );
  NAND2_X1 U953 ( .A1(n853), .A2(n852), .ZN(n857) );
  NAND2_X1 U954 ( .A1(G136), .A2(n885), .ZN(n855) );
  NAND2_X1 U955 ( .A1(G112), .A2(n878), .ZN(n854) );
  NAND2_X1 U956 ( .A1(n855), .A2(n854), .ZN(n856) );
  NOR2_X1 U957 ( .A1(n857), .A2(n856), .ZN(G162) );
  XNOR2_X1 U958 ( .A(G160), .B(n858), .ZN(n860) );
  XNOR2_X1 U959 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U960 ( .A(n861), .B(KEYINPUT48), .Z(n866) );
  XNOR2_X1 U961 ( .A(G162), .B(n862), .ZN(n863) );
  XNOR2_X1 U962 ( .A(n863), .B(n990), .ZN(n864) );
  XNOR2_X1 U963 ( .A(n864), .B(KEYINPUT46), .ZN(n865) );
  XNOR2_X1 U964 ( .A(n866), .B(n865), .ZN(n876) );
  NAND2_X1 U965 ( .A1(G130), .A2(n877), .ZN(n868) );
  NAND2_X1 U966 ( .A1(G118), .A2(n878), .ZN(n867) );
  NAND2_X1 U967 ( .A1(n868), .A2(n867), .ZN(n874) );
  NAND2_X1 U968 ( .A1(n885), .A2(G142), .ZN(n869) );
  XNOR2_X1 U969 ( .A(n869), .B(KEYINPUT112), .ZN(n871) );
  NAND2_X1 U970 ( .A1(G106), .A2(n882), .ZN(n870) );
  NAND2_X1 U971 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U972 ( .A(n872), .B(KEYINPUT45), .Z(n873) );
  NOR2_X1 U973 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U974 ( .A(n876), .B(n875), .Z(n890) );
  NAND2_X1 U975 ( .A1(G127), .A2(n877), .ZN(n880) );
  NAND2_X1 U976 ( .A1(G115), .A2(n878), .ZN(n879) );
  NAND2_X1 U977 ( .A1(n880), .A2(n879), .ZN(n881) );
  XNOR2_X1 U978 ( .A(n881), .B(KEYINPUT47), .ZN(n884) );
  NAND2_X1 U979 ( .A1(G103), .A2(n882), .ZN(n883) );
  NAND2_X1 U980 ( .A1(n884), .A2(n883), .ZN(n888) );
  NAND2_X1 U981 ( .A1(G139), .A2(n885), .ZN(n886) );
  XNOR2_X1 U982 ( .A(KEYINPUT113), .B(n886), .ZN(n887) );
  NOR2_X1 U983 ( .A1(n888), .A2(n887), .ZN(n1001) );
  XOR2_X1 U984 ( .A(n1001), .B(G164), .Z(n889) );
  XNOR2_X1 U985 ( .A(n890), .B(n889), .ZN(n891) );
  NOR2_X1 U986 ( .A1(G37), .A2(n891), .ZN(G395) );
  XNOR2_X1 U987 ( .A(n954), .B(n892), .ZN(n894) );
  XNOR2_X1 U988 ( .A(G171), .B(n938), .ZN(n893) );
  XNOR2_X1 U989 ( .A(n894), .B(n893), .ZN(n895) );
  XNOR2_X1 U990 ( .A(n895), .B(G286), .ZN(n896) );
  NOR2_X1 U991 ( .A1(G37), .A2(n896), .ZN(G397) );
  NOR2_X1 U992 ( .A1(G227), .A2(G229), .ZN(n898) );
  XNOR2_X1 U993 ( .A(KEYINPUT49), .B(KEYINPUT114), .ZN(n897) );
  XNOR2_X1 U994 ( .A(n898), .B(n897), .ZN(n910) );
  XOR2_X1 U995 ( .A(KEYINPUT102), .B(G2446), .Z(n900) );
  XNOR2_X1 U996 ( .A(G2443), .B(G2454), .ZN(n899) );
  XNOR2_X1 U997 ( .A(n900), .B(n899), .ZN(n901) );
  XOR2_X1 U998 ( .A(n901), .B(G2451), .Z(n903) );
  XNOR2_X1 U999 ( .A(G1341), .B(G1348), .ZN(n902) );
  XNOR2_X1 U1000 ( .A(n903), .B(n902), .ZN(n907) );
  XOR2_X1 U1001 ( .A(G2435), .B(G2427), .Z(n905) );
  XNOR2_X1 U1002 ( .A(G2430), .B(G2438), .ZN(n904) );
  XNOR2_X1 U1003 ( .A(n905), .B(n904), .ZN(n906) );
  XOR2_X1 U1004 ( .A(n907), .B(n906), .Z(n908) );
  NAND2_X1 U1005 ( .A1(G14), .A2(n908), .ZN(n913) );
  NAND2_X1 U1006 ( .A1(n913), .A2(G319), .ZN(n909) );
  NOR2_X1 U1007 ( .A1(n910), .A2(n909), .ZN(n912) );
  NOR2_X1 U1008 ( .A1(G395), .A2(G397), .ZN(n911) );
  NAND2_X1 U1009 ( .A1(n912), .A2(n911), .ZN(G225) );
  INV_X1 U1010 ( .A(G225), .ZN(G308) );
  INV_X1 U1011 ( .A(G69), .ZN(G235) );
  INV_X1 U1012 ( .A(n913), .ZN(G401) );
  XNOR2_X1 U1013 ( .A(KEYINPUT123), .B(G1961), .ZN(n914) );
  XNOR2_X1 U1014 ( .A(n914), .B(G5), .ZN(n924) );
  XNOR2_X1 U1015 ( .A(G1971), .B(G22), .ZN(n916) );
  XNOR2_X1 U1016 ( .A(G23), .B(G1976), .ZN(n915) );
  NOR2_X1 U1017 ( .A1(n916), .A2(n915), .ZN(n917) );
  XOR2_X1 U1018 ( .A(KEYINPUT124), .B(n917), .Z(n919) );
  XNOR2_X1 U1019 ( .A(G1986), .B(G24), .ZN(n918) );
  NOR2_X1 U1020 ( .A1(n919), .A2(n918), .ZN(n920) );
  XOR2_X1 U1021 ( .A(KEYINPUT58), .B(n920), .Z(n922) );
  XNOR2_X1 U1022 ( .A(G1966), .B(G21), .ZN(n921) );
  NOR2_X1 U1023 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1024 ( .A1(n924), .A2(n923), .ZN(n934) );
  XOR2_X1 U1025 ( .A(G1348), .B(KEYINPUT59), .Z(n925) );
  XNOR2_X1 U1026 ( .A(G4), .B(n925), .ZN(n927) );
  XNOR2_X1 U1027 ( .A(G20), .B(G1956), .ZN(n926) );
  NOR2_X1 U1028 ( .A1(n927), .A2(n926), .ZN(n931) );
  XNOR2_X1 U1029 ( .A(G1981), .B(G6), .ZN(n929) );
  XNOR2_X1 U1030 ( .A(G1341), .B(G19), .ZN(n928) );
  NOR2_X1 U1031 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1032 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1033 ( .A(KEYINPUT60), .B(n932), .ZN(n933) );
  NOR2_X1 U1034 ( .A1(n934), .A2(n933), .ZN(n935) );
  XOR2_X1 U1035 ( .A(KEYINPUT61), .B(n935), .Z(n936) );
  NOR2_X1 U1036 ( .A1(G16), .A2(n936), .ZN(n937) );
  XNOR2_X1 U1037 ( .A(KEYINPUT125), .B(n937), .ZN(n965) );
  XNOR2_X1 U1038 ( .A(KEYINPUT56), .B(G16), .ZN(n963) );
  XNOR2_X1 U1039 ( .A(G301), .B(G1961), .ZN(n940) );
  XOR2_X1 U1040 ( .A(n938), .B(G1348), .Z(n939) );
  NOR2_X1 U1041 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1042 ( .A(KEYINPUT120), .B(n941), .ZN(n952) );
  NAND2_X1 U1043 ( .A1(G1971), .A2(G303), .ZN(n942) );
  NAND2_X1 U1044 ( .A1(n943), .A2(n942), .ZN(n945) );
  XNOR2_X1 U1045 ( .A(G1956), .B(G299), .ZN(n944) );
  NOR2_X1 U1046 ( .A1(n945), .A2(n944), .ZN(n947) );
  NAND2_X1 U1047 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1048 ( .A(KEYINPUT121), .B(n948), .Z(n949) );
  NOR2_X1 U1049 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1050 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1051 ( .A(KEYINPUT122), .B(n953), .ZN(n956) );
  XNOR2_X1 U1052 ( .A(G1341), .B(n954), .ZN(n955) );
  NOR2_X1 U1053 ( .A1(n956), .A2(n955), .ZN(n961) );
  XOR2_X1 U1054 ( .A(G168), .B(G1966), .Z(n957) );
  NOR2_X1 U1055 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1056 ( .A(KEYINPUT57), .B(n959), .Z(n960) );
  NAND2_X1 U1057 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1060 ( .A(n966), .B(KEYINPUT126), .ZN(n1021) );
  XOR2_X1 U1061 ( .A(G2084), .B(G34), .Z(n967) );
  XNOR2_X1 U1062 ( .A(KEYINPUT54), .B(n967), .ZN(n984) );
  XNOR2_X1 U1063 ( .A(G2090), .B(G35), .ZN(n982) );
  XOR2_X1 U1064 ( .A(G1991), .B(G25), .Z(n968) );
  NAND2_X1 U1065 ( .A1(n968), .A2(G28), .ZN(n979) );
  XOR2_X1 U1066 ( .A(n969), .B(G27), .Z(n972) );
  XOR2_X1 U1067 ( .A(n970), .B(G32), .Z(n971) );
  NOR2_X1 U1068 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1069 ( .A(KEYINPUT118), .B(n973), .ZN(n977) );
  XNOR2_X1 U1070 ( .A(G2067), .B(G26), .ZN(n975) );
  XNOR2_X1 U1071 ( .A(G33), .B(G2072), .ZN(n974) );
  NOR2_X1 U1072 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1073 ( .A1(n977), .A2(n976), .ZN(n978) );
  NOR2_X1 U1074 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1075 ( .A(KEYINPUT53), .B(n980), .ZN(n981) );
  NOR2_X1 U1076 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1078 ( .A(n985), .B(KEYINPUT119), .ZN(n986) );
  XOR2_X1 U1079 ( .A(KEYINPUT55), .B(KEYINPUT116), .Z(n1013) );
  XNOR2_X1 U1080 ( .A(n986), .B(n1013), .ZN(n987) );
  NOR2_X1 U1081 ( .A1(G29), .A2(n987), .ZN(n1018) );
  XOR2_X1 U1082 ( .A(G160), .B(G2084), .Z(n988) );
  NOR2_X1 U1083 ( .A1(n989), .A2(n988), .ZN(n991) );
  NAND2_X1 U1084 ( .A1(n991), .A2(n990), .ZN(n1011) );
  XNOR2_X1 U1085 ( .A(G162), .B(n992), .ZN(n993) );
  NOR2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1087 ( .A(n995), .B(KEYINPUT51), .ZN(n996) );
  NOR2_X1 U1088 ( .A1(n997), .A2(n996), .ZN(n1009) );
  INV_X1 U1089 ( .A(n998), .ZN(n1000) );
  NAND2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1007) );
  XNOR2_X1 U1091 ( .A(G2072), .B(n1001), .ZN(n1003) );
  XNOR2_X1 U1092 ( .A(G164), .B(G2078), .ZN(n1002) );
  NAND2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XOR2_X1 U1094 ( .A(KEYINPUT50), .B(n1004), .Z(n1005) );
  XNOR2_X1 U1095 ( .A(KEYINPUT115), .B(n1005), .ZN(n1006) );
  NOR2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NOR2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1099 ( .A(KEYINPUT52), .B(n1012), .ZN(n1014) );
  NAND2_X1 U1100 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1101 ( .A1(n1015), .A2(G29), .ZN(n1016) );
  XNOR2_X1 U1102 ( .A(KEYINPUT117), .B(n1016), .ZN(n1017) );
  NOR2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1104 ( .A1(G11), .A2(n1019), .ZN(n1020) );
  NOR2_X1 U1105 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XOR2_X1 U1106 ( .A(KEYINPUT62), .B(n1022), .Z(n1023) );
  XNOR2_X1 U1107 ( .A(KEYINPUT127), .B(n1023), .ZN(G311) );
  INV_X1 U1108 ( .A(G311), .ZN(G150) );
endmodule

