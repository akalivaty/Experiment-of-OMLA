//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 1 0 1 0 1 1 1 0 1 1 1 0 1 1 1 1 0 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 0 0 0 0 0 0 1 1 1 0 0 0 1 1 0 1 0 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:46 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1298, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G68), .A3(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(G13), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  XOR2_X1   g0015(.A(KEYINPUT64), .B(KEYINPUT0), .Z(new_n216));
  XNOR2_X1  g0016(.A(new_n215), .B(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(G50), .B1(G58), .B2(G68), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n220), .A2(new_n210), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(KEYINPUT1), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT65), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n228));
  AND3_X1   g0028(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n211), .B1(new_n225), .B2(new_n229), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n217), .B(new_n222), .C1(new_n223), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(new_n223), .B2(new_n230), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  INV_X1    g0033(.A(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(KEYINPUT2), .B(G226), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G358));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G107), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(KEYINPUT81), .ZN(new_n249));
  INV_X1    g0049(.A(G1698), .ZN(new_n250));
  AND2_X1   g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  NOR2_X1   g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  OAI211_X1 g0052(.A(G257), .B(new_n250), .C1(new_n251), .C2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT80), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT3), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND4_X1  g0060(.A1(new_n260), .A2(KEYINPUT80), .A3(G257), .A4(new_n250), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n251), .A2(new_n252), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G303), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n260), .A2(G264), .A3(G1698), .ZN(new_n264));
  NAND4_X1  g0064(.A1(new_n255), .A2(new_n261), .A3(new_n263), .A4(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n220), .ZN(new_n266));
  NAND2_X1  g0066(.A1(G33), .A2(G41), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n265), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n209), .A2(G45), .ZN(new_n271));
  OR2_X1    g0071(.A1(KEYINPUT5), .A2(G41), .ZN(new_n272));
  NAND2_X1  g0072(.A1(KEYINPUT5), .A2(G41), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT66), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n267), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(KEYINPUT66), .A2(G33), .A3(G41), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n276), .A2(new_n266), .A3(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n274), .A2(new_n278), .A3(G274), .ZN(new_n279));
  INV_X1    g0079(.A(G45), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n280), .A2(G1), .ZN(new_n281));
  INV_X1    g0081(.A(new_n273), .ZN(new_n282));
  NOR2_X1   g0082(.A1(KEYINPUT5), .A2(G41), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n281), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n278), .A2(new_n284), .A3(G270), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n279), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n270), .A2(G179), .A3(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G116), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n209), .A2(G33), .ZN(new_n293));
  NAND3_X1  g0093(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n294));
  NAND4_X1  g0094(.A1(new_n289), .A2(new_n293), .A3(new_n220), .A4(new_n294), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n292), .B1(new_n295), .B2(new_n291), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT20), .ZN(new_n297));
  NAND2_X1  g0097(.A1(G33), .A2(G283), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(new_n210), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n205), .A2(KEYINPUT77), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT77), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G97), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n299), .B1(new_n303), .B2(new_n257), .ZN(new_n304));
  AOI22_X1  g0104(.A1(new_n294), .A2(new_n220), .B1(G20), .B2(new_n291), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n297), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(G33), .B1(new_n300), .B2(new_n302), .ZN(new_n308));
  OAI211_X1 g0108(.A(KEYINPUT20), .B(new_n305), .C1(new_n308), .C2(new_n299), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n296), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n249), .B1(new_n288), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n310), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n286), .B1(new_n265), .B2(new_n269), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n312), .A2(new_n313), .A3(KEYINPUT81), .A4(G179), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT21), .ZN(new_n316));
  INV_X1    g0116(.A(G169), .ZN(new_n317));
  NOR4_X1   g0117(.A1(new_n313), .A2(new_n310), .A3(new_n316), .A4(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n307), .A2(new_n309), .ZN(new_n320));
  INV_X1    g0120(.A(new_n296), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n317), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n270), .A2(new_n287), .ZN(new_n323));
  AOI21_X1  g0123(.A(KEYINPUT21), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  AND3_X1   g0125(.A1(new_n315), .A2(new_n319), .A3(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT70), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT9), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n290), .A2(new_n201), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n289), .A2(new_n220), .A3(new_n294), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n209), .A2(G20), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G50), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n329), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT68), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n329), .B(KEYINPUT68), .C1(new_n330), .C2(new_n332), .ZN(new_n336));
  AND2_X1   g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(G20), .B1(new_n203), .B2(G68), .ZN(new_n338));
  INV_X1    g0138(.A(G150), .ZN(new_n339));
  NOR2_X1   g0139(.A1(G20), .A2(G33), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n210), .A2(G33), .ZN(new_n342));
  XNOR2_X1  g0142(.A(KEYINPUT8), .B(G58), .ZN(new_n343));
  OAI221_X1 g0143(.A(new_n338), .B1(new_n339), .B2(new_n341), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n294), .A2(new_n220), .ZN(new_n345));
  AND2_X1   g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n327), .B(new_n328), .C1(new_n337), .C2(new_n346), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n335), .A2(new_n336), .B1(new_n344), .B2(new_n345), .ZN(new_n348));
  OAI21_X1  g0148(.A(KEYINPUT70), .B1(new_n348), .B2(KEYINPUT9), .ZN(new_n349));
  AND2_X1   g0149(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n260), .A2(new_n250), .ZN(new_n351));
  INV_X1    g0151(.A(G222), .ZN(new_n352));
  INV_X1    g0152(.A(G77), .ZN(new_n353));
  OAI22_X1  g0153(.A1(new_n351), .A2(new_n352), .B1(new_n353), .B2(new_n260), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(G1698), .B1(new_n251), .B2(new_n252), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(KEYINPUT67), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT67), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n358), .B(G1698), .C1(new_n251), .C2(new_n252), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(G223), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n268), .B1(new_n355), .B2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(G41), .ZN(new_n363));
  AOI21_X1  g0163(.A(G1), .B1(new_n363), .B2(new_n280), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n220), .B1(new_n275), .B2(new_n267), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n364), .B1(new_n365), .B2(new_n277), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(G226), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n278), .A2(G274), .A3(new_n364), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(G200), .B1(new_n362), .B2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n369), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n354), .B1(new_n360), .B2(G223), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n371), .B(G190), .C1(new_n372), .C2(new_n268), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT71), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n348), .A2(KEYINPUT9), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n370), .A2(new_n373), .A3(new_n374), .A4(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(KEYINPUT10), .B1(new_n350), .B2(new_n376), .ZN(new_n377));
  AND2_X1   g0177(.A1(new_n370), .A2(new_n375), .ZN(new_n378));
  AND2_X1   g0178(.A1(new_n373), .A2(new_n374), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT10), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n347), .A2(new_n349), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n378), .A2(new_n379), .A3(new_n380), .A4(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n377), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n371), .B1(new_n372), .B2(new_n268), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n348), .B1(new_n384), .B2(new_n317), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n385), .B1(G179), .B2(new_n384), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n260), .A2(KEYINPUT69), .A3(G232), .A4(new_n250), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT69), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n388), .B1(new_n262), .B2(G107), .ZN(new_n389));
  OAI211_X1 g0189(.A(G232), .B(new_n250), .C1(new_n251), .C2(new_n252), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n387), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(G238), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n393), .B1(new_n357), .B2(new_n359), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n269), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n366), .A2(G244), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n368), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n395), .A2(G190), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n331), .A2(G77), .ZN(new_n400));
  OAI22_X1  g0200(.A1(new_n330), .A2(new_n400), .B1(G77), .B2(new_n289), .ZN(new_n401));
  NAND2_X1  g0201(.A1(G20), .A2(G77), .ZN(new_n402));
  XNOR2_X1  g0202(.A(KEYINPUT15), .B(G87), .ZN(new_n403));
  OAI221_X1 g0203(.A(new_n402), .B1(new_n403), .B2(new_n342), .C1(new_n341), .C2(new_n343), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n401), .B1(new_n404), .B2(new_n345), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n358), .B1(new_n260), .B2(G1698), .ZN(new_n406));
  INV_X1    g0206(.A(new_n359), .ZN(new_n407));
  OAI21_X1  g0207(.A(G238), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(KEYINPUT69), .B1(new_n260), .B2(new_n206), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(new_n390), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n408), .A2(new_n387), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n397), .B1(new_n411), .B2(new_n269), .ZN(new_n412));
  INV_X1    g0212(.A(G200), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n399), .B(new_n405), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n395), .A2(new_n398), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n405), .B1(new_n415), .B2(new_n317), .ZN(new_n416));
  INV_X1    g0216(.A(G179), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n412), .A2(new_n417), .ZN(new_n418));
  AND2_X1   g0218(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n383), .A2(new_n386), .A3(new_n414), .A4(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n234), .A2(G1698), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(G226), .B2(G1698), .ZN(new_n423));
  OAI22_X1  g0223(.A1(new_n423), .A2(new_n262), .B1(new_n257), .B2(new_n205), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n269), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT13), .ZN(new_n426));
  INV_X1    g0226(.A(new_n364), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n278), .A2(new_n427), .A3(G238), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n425), .A2(new_n426), .A3(new_n368), .A4(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT72), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(G226), .A2(G1698), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n432), .B1(new_n234), .B2(G1698), .ZN(new_n433));
  AOI22_X1  g0233(.A1(new_n433), .A2(new_n260), .B1(G33), .B2(G97), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n368), .B(new_n428), .C1(new_n434), .C2(new_n268), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n417), .B1(new_n435), .B2(KEYINPUT13), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n424), .A2(new_n269), .B1(new_n366), .B2(G238), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n437), .A2(KEYINPUT72), .A3(new_n426), .A4(new_n368), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n431), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT74), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT74), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n431), .A2(new_n436), .A3(new_n438), .A4(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT14), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n435), .A2(KEYINPUT13), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(new_n429), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n444), .B1(new_n446), .B2(G169), .ZN(new_n447));
  AOI211_X1 g0247(.A(KEYINPUT14), .B(new_n317), .C1(new_n445), .C2(new_n429), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n443), .A2(new_n449), .ZN(new_n450));
  OAI22_X1  g0250(.A1(new_n341), .A2(new_n201), .B1(new_n210), .B2(G68), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n342), .A2(new_n353), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n345), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  XNOR2_X1  g0253(.A(new_n453), .B(KEYINPUT11), .ZN(new_n454));
  INV_X1    g0254(.A(G68), .ZN(new_n455));
  AOI21_X1  g0255(.A(KEYINPUT73), .B1(new_n290), .B2(new_n455), .ZN(new_n456));
  XNOR2_X1  g0256(.A(new_n456), .B(KEYINPUT12), .ZN(new_n457));
  INV_X1    g0257(.A(new_n330), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n458), .A2(G68), .A3(new_n331), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n454), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n450), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n460), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n431), .A2(G190), .A3(new_n438), .A4(new_n445), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n446), .A2(G200), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n278), .A2(new_n427), .A3(G232), .ZN(new_n467));
  NAND2_X1  g0267(.A1(G33), .A2(G87), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT76), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(KEYINPUT76), .A2(G33), .A3(G87), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(G223), .A2(G1698), .ZN(new_n473));
  INV_X1    g0273(.A(G226), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n473), .B1(new_n474), .B2(G1698), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n472), .B1(new_n260), .B2(new_n475), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n368), .B(new_n467), .C1(new_n476), .C2(new_n268), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(new_n317), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n478), .B1(G179), .B2(new_n477), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n258), .A2(new_n210), .A3(new_n259), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT7), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n258), .A2(KEYINPUT7), .A3(new_n210), .A4(new_n259), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n455), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n202), .A2(new_n455), .ZN(new_n485));
  NOR2_X1   g0285(.A1(G58), .A2(G68), .ZN(new_n486));
  OAI21_X1  g0286(.A(G20), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(G159), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n487), .B1(new_n488), .B2(new_n341), .ZN(new_n489));
  OAI21_X1  g0289(.A(KEYINPUT75), .B1(new_n484), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(KEYINPUT16), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT16), .ZN(new_n492));
  OAI211_X1 g0292(.A(KEYINPUT75), .B(new_n492), .C1(new_n484), .C2(new_n489), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n491), .A2(new_n345), .A3(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(new_n343), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n331), .ZN(new_n496));
  OAI22_X1  g0296(.A1(new_n496), .A2(new_n330), .B1(new_n289), .B2(new_n495), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n479), .B1(new_n494), .B2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT18), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n490), .A2(KEYINPUT16), .B1(new_n220), .B2(new_n294), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n497), .B1(new_n502), .B2(new_n493), .ZN(new_n503));
  OAI21_X1  g0303(.A(KEYINPUT18), .B1(new_n503), .B2(new_n479), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n477), .A2(new_n413), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n505), .B1(G190), .B2(new_n477), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n494), .A2(new_n498), .A3(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT17), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n503), .A2(KEYINPUT17), .A3(new_n506), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n501), .A2(new_n504), .A3(new_n509), .A4(new_n510), .ZN(new_n511));
  NOR3_X1   g0311(.A1(new_n421), .A2(new_n466), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n413), .B1(new_n270), .B2(new_n287), .ZN(new_n513));
  OAI21_X1  g0313(.A(KEYINPUT82), .B1(new_n513), .B2(new_n312), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT82), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n515), .B(new_n310), .C1(new_n313), .C2(new_n413), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n313), .A2(G190), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n514), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT83), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT83), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n514), .A2(new_n517), .A3(new_n520), .A4(new_n516), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT23), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n523), .B1(new_n210), .B2(G107), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n210), .A2(G33), .A3(G116), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n210), .B(G87), .C1(new_n251), .C2(new_n252), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(KEYINPUT22), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT22), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n260), .A2(new_n531), .A3(new_n210), .A4(G87), .ZN(new_n532));
  AOI211_X1 g0332(.A(KEYINPUT24), .B(new_n528), .C1(new_n530), .C2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT24), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n530), .A2(new_n532), .ZN(new_n535));
  INV_X1    g0335(.A(new_n528), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n345), .B1(new_n533), .B2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n295), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n290), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT25), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(new_n289), .B2(G107), .ZN(new_n542));
  AOI22_X1  g0342(.A1(G107), .A2(new_n539), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n538), .A2(new_n543), .ZN(new_n544));
  OAI211_X1 g0344(.A(G257), .B(G1698), .C1(new_n251), .C2(new_n252), .ZN(new_n545));
  OAI211_X1 g0345(.A(G250), .B(new_n250), .C1(new_n251), .C2(new_n252), .ZN(new_n546));
  NAND2_X1  g0346(.A1(G33), .A2(G294), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT84), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n268), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n545), .A2(new_n546), .A3(KEYINPUT84), .A4(new_n547), .ZN(new_n551));
  AND2_X1   g0351(.A1(new_n278), .A2(new_n284), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n550), .A2(new_n551), .B1(G264), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n553), .A2(new_n417), .A3(new_n279), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n548), .A2(new_n549), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n555), .A2(new_n269), .A3(new_n551), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n552), .A2(G264), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n556), .A2(new_n279), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n317), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n544), .A2(new_n554), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n558), .A2(G200), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n553), .A2(G190), .A3(new_n279), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n561), .A2(new_n562), .A3(new_n538), .A4(new_n543), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n289), .A2(G97), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n565), .B1(new_n539), .B2(G97), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(KEYINPUT7), .B1(new_n262), .B2(new_n210), .ZN(new_n568));
  INV_X1    g0368(.A(new_n483), .ZN(new_n569));
  OAI21_X1  g0369(.A(G107), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n340), .A2(G77), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n206), .A2(KEYINPUT6), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n572), .B1(new_n300), .B2(new_n302), .ZN(new_n573));
  NAND2_X1  g0373(.A1(G97), .A2(G107), .ZN(new_n574));
  AOI21_X1  g0374(.A(KEYINPUT6), .B1(new_n207), .B2(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(G20), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n570), .A2(new_n571), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n567), .B1(new_n577), .B2(new_n345), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n278), .A2(new_n284), .A3(G257), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n279), .A2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  AND2_X1   g0381(.A1(KEYINPUT4), .A2(G244), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n250), .B(new_n582), .C1(new_n251), .C2(new_n252), .ZN(new_n583));
  INV_X1    g0383(.A(G244), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n584), .B1(new_n258), .B2(new_n259), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n583), .B(new_n298), .C1(new_n585), .C2(KEYINPUT4), .ZN(new_n586));
  OAI21_X1  g0386(.A(G250), .B1(new_n251), .B2(new_n252), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n250), .B1(new_n587), .B2(KEYINPUT4), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n269), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n581), .A2(new_n589), .A3(G190), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT78), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n580), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n279), .A2(new_n579), .A3(KEYINPUT78), .ZN(new_n593));
  INV_X1    g0393(.A(G250), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n594), .B1(new_n258), .B2(new_n259), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT4), .ZN(new_n596));
  OAI21_X1  g0396(.A(G1698), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n596), .B1(new_n262), .B2(new_n584), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n597), .A2(new_n298), .A3(new_n583), .A4(new_n598), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n592), .A2(new_n593), .B1(new_n599), .B2(new_n269), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n578), .B(new_n590), .C1(new_n600), .C2(new_n413), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n581), .A2(new_n589), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n317), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n576), .A2(new_n571), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n206), .B1(new_n482), .B2(new_n483), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n345), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n566), .ZN(new_n607));
  AND3_X1   g0407(.A1(new_n279), .A2(new_n579), .A3(KEYINPUT78), .ZN(new_n608));
  AOI21_X1  g0408(.A(KEYINPUT78), .B1(new_n279), .B2(new_n579), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n417), .B(new_n589), .C1(new_n608), .C2(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n603), .A2(new_n607), .A3(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n403), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n612), .A2(new_n289), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT19), .ZN(new_n614));
  XNOR2_X1  g0414(.A(KEYINPUT77), .B(G97), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n614), .B1(new_n615), .B2(new_n342), .ZN(new_n616));
  NOR2_X1   g0416(.A1(G87), .A2(G107), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n300), .A2(new_n302), .A3(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n210), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n260), .A2(new_n210), .A3(G68), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n616), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n613), .B1(new_n623), .B2(new_n345), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n539), .A2(new_n612), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(G33), .A2(G116), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n393), .A2(new_n250), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n584), .A2(G1698), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n627), .B1(new_n630), .B2(new_n262), .ZN(new_n631));
  AOI21_X1  g0431(.A(G250), .B1(new_n209), .B2(G45), .ZN(new_n632));
  INV_X1    g0432(.A(G274), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n632), .B1(new_n633), .B2(new_n281), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n631), .A2(new_n269), .B1(new_n634), .B2(new_n278), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n317), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n635), .A2(new_n417), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n626), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(G87), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n295), .A2(new_n640), .ZN(new_n641));
  AOI211_X1 g0441(.A(new_n613), .B(new_n641), .C1(new_n623), .C2(new_n345), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n636), .A2(G200), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n634), .A2(new_n278), .ZN(new_n644));
  NOR2_X1   g0444(.A1(G238), .A2(G1698), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n645), .B1(new_n584), .B2(G1698), .ZN(new_n646));
  AOI22_X1  g0446(.A1(new_n646), .A2(new_n260), .B1(G33), .B2(G116), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n644), .B(G190), .C1(new_n647), .C2(new_n268), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n648), .A2(KEYINPUT79), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT79), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n650), .B1(new_n635), .B2(G190), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n642), .B(new_n643), .C1(new_n649), .C2(new_n651), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n601), .A2(new_n611), .A3(new_n639), .A4(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n564), .A2(new_n653), .ZN(new_n654));
  AND4_X1   g0454(.A1(new_n326), .A2(new_n512), .A3(new_n522), .A4(new_n654), .ZN(G372));
  INV_X1    g0455(.A(new_n386), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n501), .A2(new_n504), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n461), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n659), .B1(new_n465), .B2(new_n419), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n509), .A2(new_n510), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n658), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT86), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n383), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n377), .A2(new_n382), .A3(KEYINPUT86), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n656), .B1(new_n662), .B2(new_n666), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n603), .A2(new_n607), .A3(new_n610), .ZN(new_n668));
  OAI21_X1  g0468(.A(KEYINPUT85), .B1(new_n647), .B2(new_n268), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT85), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n631), .A2(new_n670), .A3(new_n269), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n644), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n317), .ZN(new_n674));
  AOI22_X1  g0474(.A1(new_n624), .A2(new_n625), .B1(new_n417), .B2(new_n635), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT26), .ZN(new_n677));
  AOI22_X1  g0477(.A1(new_n669), .A2(new_n671), .B1(new_n278), .B2(new_n634), .ZN(new_n678));
  OAI211_X1 g0478(.A(new_n642), .B(new_n648), .C1(new_n678), .C2(new_n413), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n668), .A2(new_n676), .A3(new_n677), .A4(new_n679), .ZN(new_n680));
  AOI22_X1  g0480(.A1(new_n317), .A2(new_n602), .B1(new_n606), .B2(new_n566), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n652), .A2(new_n681), .A3(new_n639), .A4(new_n610), .ZN(new_n682));
  AOI22_X1  g0482(.A1(new_n682), .A2(KEYINPUT26), .B1(new_n675), .B2(new_n674), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n318), .A2(new_n324), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n684), .A2(new_n315), .A3(new_n560), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n413), .B1(new_n672), .B2(new_n644), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  OAI211_X1 g0487(.A(new_n624), .B(new_n648), .C1(new_n640), .C2(new_n295), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  AOI22_X1  g0489(.A1(new_n687), .A2(new_n689), .B1(new_n674), .B2(new_n675), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n690), .A2(new_n563), .A3(new_n611), .A4(new_n601), .ZN(new_n691));
  OAI211_X1 g0491(.A(new_n680), .B(new_n683), .C1(new_n685), .C2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n512), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n667), .A2(new_n693), .ZN(G369));
  NAND3_X1  g0494(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(KEYINPUT27), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT27), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n697), .A2(new_n209), .A3(new_n210), .A4(G13), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n696), .A2(G213), .A3(new_n698), .ZN(new_n699));
  XOR2_X1   g0499(.A(new_n699), .B(KEYINPUT87), .Z(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(G343), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n544), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n560), .A2(new_n563), .A3(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT89), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n560), .A2(new_n563), .A3(KEYINPUT89), .A4(new_n703), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OR2_X1    g0508(.A1(new_n560), .A2(new_n701), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n702), .A2(new_n312), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n522), .A2(new_n326), .A3(new_n711), .ZN(new_n712));
  OR2_X1    g0512(.A1(new_n326), .A2(new_n711), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT88), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n714), .A2(new_n715), .A3(G330), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n715), .B1(new_n714), .B2(G330), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n710), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  OR2_X1    g0519(.A1(new_n560), .A2(new_n702), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n326), .A2(new_n702), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n721), .A2(new_n707), .A3(new_n706), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n719), .A2(new_n720), .A3(new_n722), .ZN(G399));
  NAND3_X1  g0523(.A1(new_n615), .A2(new_n291), .A3(new_n617), .ZN(new_n724));
  XNOR2_X1  g0524(.A(new_n724), .B(KEYINPUT90), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n213), .A2(G41), .ZN(new_n726));
  NOR3_X1   g0526(.A1(new_n725), .A2(new_n209), .A3(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n727), .B1(new_n219), .B2(new_n726), .ZN(new_n728));
  XOR2_X1   g0528(.A(new_n728), .B(KEYINPUT91), .Z(new_n729));
  XNOR2_X1  g0529(.A(new_n729), .B(KEYINPUT28), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n522), .A2(new_n654), .A3(new_n326), .A4(new_n701), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT30), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n553), .A2(new_n635), .A3(new_n589), .A4(new_n581), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n732), .B1(new_n733), .B2(new_n288), .ZN(new_n734));
  INV_X1    g0534(.A(new_n288), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n602), .A2(new_n636), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n735), .A2(new_n736), .A3(KEYINPUT30), .A4(new_n553), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n589), .B1(new_n608), .B2(new_n609), .ZN(new_n739));
  AND3_X1   g0539(.A1(new_n558), .A2(new_n739), .A3(KEYINPUT92), .ZN(new_n740));
  AOI21_X1  g0540(.A(KEYINPUT92), .B1(new_n558), .B2(new_n739), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n673), .A2(new_n417), .A3(new_n323), .ZN(new_n742));
  NOR3_X1   g0542(.A1(new_n740), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n702), .B1(new_n738), .B2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT31), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  OAI211_X1 g0546(.A(KEYINPUT31), .B(new_n702), .C1(new_n738), .C2(new_n743), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n731), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G330), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n692), .A2(new_n701), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT93), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT29), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n652), .A2(new_n639), .ZN(new_n755));
  OAI21_X1  g0555(.A(KEYINPUT26), .B1(new_n755), .B2(new_n611), .ZN(new_n756));
  AND3_X1   g0556(.A1(new_n756), .A2(new_n680), .A3(new_n676), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n684), .A2(new_n315), .A3(new_n560), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n601), .A2(new_n611), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n626), .A2(new_n638), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n678), .A2(G169), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n679), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n758), .A2(new_n763), .A3(new_n563), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n702), .B1(new_n757), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(KEYINPUT93), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n753), .A2(new_n754), .A3(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(KEYINPUT26), .B1(new_n762), .B2(new_n611), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n668), .A2(new_n677), .A3(new_n639), .A4(new_n652), .ZN(new_n769));
  AND3_X1   g0569(.A1(new_n768), .A2(new_n676), .A3(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n702), .B1(new_n770), .B2(new_n764), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(KEYINPUT29), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n750), .B1(new_n767), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n730), .B1(new_n773), .B2(G1), .ZN(G364));
  NOR2_X1   g0574(.A1(G13), .A2(G33), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(G20), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n220), .B1(G20), .B2(new_n317), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n213), .A2(new_n260), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n782), .B1(new_n280), .B2(new_n219), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n783), .B1(new_n244), .B2(new_n280), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n213), .A2(new_n262), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n785), .A2(G355), .B1(new_n291), .B2(new_n213), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n780), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n210), .A2(new_n417), .ZN(new_n788));
  INV_X1    g0588(.A(G190), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n788), .A2(new_n789), .A3(G200), .ZN(new_n790));
  XOR2_X1   g0590(.A(KEYINPUT33), .B(G317), .Z(new_n791));
  NOR2_X1   g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n210), .A2(G190), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n417), .A2(G200), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(G311), .ZN(new_n796));
  INV_X1    g0596(.A(G322), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n210), .A2(new_n789), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(new_n794), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n262), .B1(new_n795), .B2(new_n796), .C1(new_n797), .C2(new_n799), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n788), .A2(G190), .A3(G200), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n792), .B(new_n800), .C1(G326), .C2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n417), .A2(new_n413), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n804), .B(KEYINPUT95), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(new_n793), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(G329), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n413), .A2(G179), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(KEYINPUT96), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(new_n793), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n811), .A2(new_n798), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  AOI22_X1  g0615(.A1(G283), .A2(new_n813), .B1(new_n815), .B2(G303), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n210), .B1(new_n806), .B2(G190), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(G294), .ZN(new_n819));
  NAND4_X1  g0619(.A1(new_n803), .A2(new_n809), .A3(new_n816), .A4(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n808), .A2(G159), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT32), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n818), .A2(G97), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n260), .B1(new_n799), .B2(new_n202), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n790), .A2(new_n455), .B1(new_n801), .B2(new_n201), .ZN(new_n825));
  INV_X1    g0625(.A(new_n795), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n824), .B(new_n825), .C1(G77), .C2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n813), .A2(G107), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n815), .A2(G87), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n823), .A2(new_n827), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n820), .B1(new_n822), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n787), .B1(new_n831), .B2(new_n778), .ZN(new_n832));
  INV_X1    g0632(.A(new_n777), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n832), .B1(new_n714), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n714), .A2(G330), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(KEYINPUT88), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n836), .B(new_n716), .C1(G330), .C2(new_n714), .ZN(new_n837));
  INV_X1    g0637(.A(new_n726), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n212), .A2(G20), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n209), .B1(new_n839), .B2(G45), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n838), .A2(KEYINPUT94), .A3(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT94), .ZN(new_n842));
  INV_X1    g0642(.A(new_n840), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n842), .B1(new_n726), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  MUX2_X1   g0645(.A(new_n834), .B(new_n837), .S(new_n845), .Z(new_n846));
  XOR2_X1   g0646(.A(new_n846), .B(KEYINPUT97), .Z(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(G396));
  OR2_X1    g0648(.A1(new_n701), .A2(new_n405), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n414), .A2(new_n849), .B1(new_n416), .B2(new_n418), .ZN(new_n850));
  AND3_X1   g0650(.A1(new_n416), .A2(new_n418), .A3(new_n701), .ZN(new_n851));
  OAI21_X1  g0651(.A(KEYINPUT100), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT100), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n416), .A2(new_n418), .A3(new_n701), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n701), .A2(new_n405), .ZN(new_n855));
  AND2_X1   g0655(.A1(new_n399), .A2(new_n405), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n415), .A2(G200), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n855), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n853), .B(new_n854), .C1(new_n858), .C2(new_n419), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n852), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n692), .A2(new_n701), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n753), .A2(new_n766), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n861), .B1(new_n862), .B2(new_n860), .ZN(new_n863));
  OR2_X1    g0663(.A1(new_n863), .A2(new_n749), .ZN(new_n864));
  INV_X1    g0664(.A(new_n845), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n865), .B1(new_n863), .B2(new_n749), .ZN(new_n866));
  AND2_X1   g0666(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n778), .A2(new_n775), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n865), .B1(G77), .B2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(G294), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n823), .B1(new_n871), .B2(new_n799), .ZN(new_n872));
  XOR2_X1   g0672(.A(new_n872), .B(KEYINPUT99), .Z(new_n873));
  OAI21_X1  g0673(.A(new_n262), .B1(new_n814), .B2(new_n206), .ZN(new_n874));
  XOR2_X1   g0674(.A(new_n874), .B(KEYINPUT98), .Z(new_n875));
  INV_X1    g0675(.A(G283), .ZN(new_n876));
  OAI22_X1  g0676(.A1(new_n790), .A2(new_n876), .B1(new_n795), .B2(new_n291), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n877), .B1(G303), .B2(new_n802), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n808), .A2(G311), .B1(new_n813), .B2(G87), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n875), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n813), .A2(G68), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n201), .B2(new_n814), .ZN(new_n882));
  AOI211_X1 g0682(.A(new_n262), .B(new_n882), .C1(G132), .C2(new_n808), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(new_n202), .B2(new_n817), .ZN(new_n884));
  INV_X1    g0684(.A(new_n799), .ZN(new_n885));
  AOI22_X1  g0685(.A1(G143), .A2(new_n885), .B1(new_n826), .B2(G159), .ZN(new_n886));
  INV_X1    g0686(.A(G137), .ZN(new_n887));
  OAI221_X1 g0687(.A(new_n886), .B1(new_n887), .B2(new_n801), .C1(new_n339), .C2(new_n790), .ZN(new_n888));
  XOR2_X1   g0688(.A(new_n888), .B(KEYINPUT34), .Z(new_n889));
  OAI22_X1  g0689(.A1(new_n873), .A2(new_n880), .B1(new_n884), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n870), .B1(new_n890), .B2(new_n778), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n891), .B1(new_n776), .B2(new_n860), .ZN(new_n892));
  XOR2_X1   g0692(.A(new_n892), .B(KEYINPUT101), .Z(new_n893));
  NOR2_X1   g0693(.A1(new_n867), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(G384));
  OR2_X1    g0695(.A1(new_n573), .A2(new_n575), .ZN(new_n896));
  OR2_X1    g0696(.A1(new_n896), .A2(KEYINPUT35), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(KEYINPUT35), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n897), .A2(G116), .A3(new_n221), .A4(new_n898), .ZN(new_n899));
  XOR2_X1   g0699(.A(new_n899), .B(KEYINPUT36), .Z(new_n900));
  OAI211_X1 g0700(.A(new_n219), .B(G77), .C1(new_n202), .C2(new_n455), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n201), .A2(G68), .ZN(new_n902));
  AOI211_X1 g0702(.A(new_n209), .B(G13), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n494), .A2(new_n498), .ZN(new_n905));
  INV_X1    g0705(.A(new_n479), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n905), .A2(new_n700), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT37), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n907), .A2(new_n908), .A3(new_n909), .A4(new_n507), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(KEYINPUT102), .ZN(new_n911));
  AND3_X1   g0711(.A1(new_n494), .A2(new_n498), .A3(new_n506), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n912), .A2(new_n499), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT102), .ZN(new_n914));
  NAND4_X1  g0714(.A1(new_n913), .A2(new_n914), .A3(new_n909), .A4(new_n908), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n507), .B1(new_n503), .B2(new_n479), .ZN(new_n916));
  INV_X1    g0716(.A(new_n700), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n503), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(KEYINPUT37), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n911), .A2(new_n915), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n511), .A2(new_n918), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT38), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n919), .A2(new_n910), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n925), .A2(new_n921), .A3(KEYINPUT38), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n702), .A2(new_n460), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n461), .A2(new_n465), .A3(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n465), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n460), .B(new_n702), .C1(new_n450), .C2(new_n930), .ZN(new_n931));
  AOI22_X1  g0731(.A1(new_n929), .A2(new_n931), .B1(new_n859), .B2(new_n852), .ZN(new_n932));
  AND3_X1   g0732(.A1(new_n932), .A2(new_n748), .A3(KEYINPUT40), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n927), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT40), .ZN(new_n935));
  AND3_X1   g0735(.A1(new_n925), .A2(new_n921), .A3(KEYINPUT38), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT38), .B1(new_n925), .B2(new_n921), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n932), .A2(new_n748), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n935), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n934), .A2(new_n940), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n512), .A2(new_n748), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n941), .A2(new_n942), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n943), .A2(G330), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n659), .A2(new_n701), .ZN(new_n946));
  AOI22_X1  g0746(.A1(new_n919), .A2(new_n910), .B1(new_n511), .B2(new_n918), .ZN(new_n947));
  AOI21_X1  g0747(.A(KEYINPUT39), .B1(new_n947), .B2(KEYINPUT38), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n924), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(KEYINPUT39), .B1(new_n936), .B2(new_n937), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n946), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n658), .A2(new_n700), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n861), .A2(new_n854), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n929), .A2(new_n931), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n953), .B1(new_n956), .B2(new_n938), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n951), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n767), .A2(new_n512), .A3(new_n772), .ZN(new_n959));
  AND2_X1   g0759(.A1(new_n959), .A2(new_n667), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n958), .B(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n945), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n209), .B2(new_n839), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n945), .A2(new_n961), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n904), .B1(new_n963), .B2(new_n964), .ZN(G367));
  INV_X1    g0765(.A(new_n710), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(new_n836), .B2(new_n716), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n611), .A2(new_n701), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT104), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n601), .B(new_n611), .C1(new_n578), .C2(new_n701), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n967), .A2(new_n971), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT103), .Z(new_n973));
  OR2_X1    g0773(.A1(new_n701), .A2(new_n642), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n690), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n676), .B2(new_n974), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n976), .A2(KEYINPUT43), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n973), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n971), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n979), .A2(new_n722), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n611), .B1(new_n979), .B2(new_n560), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n980), .A2(KEYINPUT42), .B1(new_n981), .B2(new_n701), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n980), .A2(KEYINPUT42), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n982), .A2(new_n983), .B1(KEYINPUT43), .B2(new_n976), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n972), .B(KEYINPUT103), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(KEYINPUT43), .B2(new_n976), .ZN(new_n986));
  AND3_X1   g0786(.A1(new_n978), .A2(new_n984), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n984), .B1(new_n978), .B2(new_n986), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n726), .B(KEYINPUT41), .Z(new_n990));
  NAND2_X1  g0790(.A1(new_n722), .A2(new_n720), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n979), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT44), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n991), .A2(KEYINPUT44), .A3(new_n979), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n722), .A2(new_n971), .A3(KEYINPUT45), .A4(new_n720), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n722), .A2(new_n971), .A3(new_n720), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT45), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n994), .A2(new_n995), .B1(new_n996), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT105), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n967), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n999), .A2(new_n996), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n995), .ZN(new_n1004));
  AOI21_X1  g0804(.A(KEYINPUT44), .B1(new_n991), .B2(new_n979), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1003), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1006), .A2(KEYINPUT105), .ZN(new_n1007));
  OAI21_X1  g0807(.A(KEYINPUT106), .B1(new_n1002), .B2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n719), .B1(new_n1006), .B2(KEYINPUT105), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT106), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n722), .B1(new_n710), .B2(new_n721), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n717), .B2(new_n718), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1013), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n836), .A2(new_n1015), .A3(new_n716), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n773), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n1006), .A2(new_n967), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1008), .A2(new_n1012), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n990), .B1(new_n1021), .B2(new_n773), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT107), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n840), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  AOI211_X1 g0824(.A(KEYINPUT107), .B(new_n990), .C1(new_n1021), .C2(new_n773), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n989), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n976), .A2(new_n833), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n780), .B1(new_n213), .B2(new_n612), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n240), .A2(new_n781), .ZN(new_n1029));
  AND2_X1   g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(G317), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n262), .B1(new_n812), .B2(new_n615), .C1(new_n807), .C2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT108), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(G303), .A2(new_n885), .B1(new_n826), .B2(G283), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1035), .B1(new_n871), .B2(new_n790), .C1(new_n796), .C2(new_n801), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n814), .A2(new_n291), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1036), .B1(KEYINPUT46), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1037), .A2(KEYINPUT46), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(G107), .B2(new_n818), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n1034), .A2(new_n1038), .A3(new_n1039), .A4(new_n1041), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n260), .B1(new_n795), .B2(new_n201), .C1(new_n790), .C2(new_n488), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n813), .A2(G77), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n887), .B2(new_n807), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n1043), .B(new_n1045), .C1(G58), .C2(new_n815), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT109), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n818), .A2(G68), .ZN(new_n1048));
  INV_X1    g0848(.A(G143), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1048), .B1(new_n1049), .B2(new_n801), .C1(new_n339), .C2(new_n799), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1046), .B1(new_n1047), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1050), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1052), .A2(KEYINPUT109), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1042), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT47), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n845), .B(new_n1030), .C1(new_n1055), .C2(new_n778), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1027), .B1(new_n1057), .B2(KEYINPUT110), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(KEYINPUT110), .B2(new_n1057), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1026), .A2(new_n1059), .ZN(G387));
  AOI21_X1  g0860(.A(new_n838), .B1(new_n1017), .B2(new_n773), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(new_n773), .B2(new_n1017), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n817), .A2(new_n876), .B1(new_n871), .B2(new_n814), .ZN(new_n1063));
  INV_X1    g0863(.A(G303), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n799), .A2(new_n1031), .B1(new_n795), .B2(new_n1064), .ZN(new_n1065));
  OR2_X1    g0865(.A1(new_n1065), .A2(KEYINPUT111), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1065), .A2(KEYINPUT111), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n790), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n1068), .A2(G311), .B1(new_n802), .B2(G322), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1066), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT48), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1063), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  OR2_X1    g0872(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1072), .A2(KEYINPUT49), .A3(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n260), .B1(new_n808), .B2(G326), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1074), .B(new_n1075), .C1(new_n291), .C2(new_n812), .ZN(new_n1076));
  AOI21_X1  g0876(.A(KEYINPUT49), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(G77), .A2(new_n815), .B1(new_n813), .B2(G97), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n339), .B2(new_n807), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n817), .A2(new_n403), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n260), .B1(new_n795), .B2(new_n455), .C1(new_n201), .C2(new_n799), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n488), .A2(new_n801), .B1(new_n790), .B2(new_n343), .ZN(new_n1083));
  NOR4_X1   g0883(.A1(new_n1080), .A2(new_n1081), .A3(new_n1082), .A4(new_n1083), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n778), .B1(new_n1078), .B2(new_n1084), .ZN(new_n1085));
  OR2_X1    g0885(.A1(new_n237), .A2(new_n280), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n1086), .A2(new_n781), .B1(new_n725), .B2(new_n785), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n495), .A2(new_n201), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT50), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n280), .B1(new_n455), .B2(new_n353), .ZN(new_n1090));
  NOR3_X1   g0890(.A1(new_n1089), .A2(new_n725), .A3(new_n1090), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n1087), .A2(new_n1091), .B1(G107), .B2(new_n214), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n845), .B1(new_n1092), .B2(new_n779), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1085), .A2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(new_n966), .B2(new_n777), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(new_n1017), .B2(new_n843), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1062), .A2(new_n1096), .ZN(G393));
  XNOR2_X1  g0897(.A(new_n1006), .B(new_n967), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n838), .B1(new_n1098), .B2(new_n1018), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1021), .A2(new_n1099), .ZN(new_n1100));
  OR2_X1    g0900(.A1(new_n1098), .A2(new_n840), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n779), .B1(new_n214), .B2(new_n615), .C1(new_n247), .C2(new_n782), .ZN(new_n1102));
  AND2_X1   g0902(.A1(new_n1102), .A2(new_n865), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n262), .B1(new_n813), .B2(G87), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n1104), .B1(new_n455), .B2(new_n814), .C1(new_n1049), .C2(new_n807), .ZN(new_n1105));
  XOR2_X1   g0905(.A(new_n1105), .B(KEYINPUT113), .Z(new_n1106));
  OAI22_X1  g0906(.A1(new_n790), .A2(new_n201), .B1(new_n795), .B2(new_n343), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n801), .A2(new_n339), .B1(new_n799), .B2(new_n488), .ZN(new_n1108));
  XOR2_X1   g0908(.A(KEYINPUT112), .B(KEYINPUT51), .Z(new_n1109));
  AOI21_X1  g0909(.A(new_n1107), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  OAI221_X1 g0910(.A(new_n1110), .B1(new_n1108), .B2(new_n1109), .C1(new_n817), .C2(new_n353), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n262), .B1(new_n795), .B2(new_n871), .C1(new_n790), .C2(new_n1064), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(new_n813), .B2(G107), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n1113), .B1(new_n876), .B2(new_n814), .C1(new_n797), .C2(new_n807), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT52), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n801), .A2(new_n1031), .B1(new_n799), .B2(new_n796), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n818), .A2(G116), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1117), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n1106), .A2(new_n1111), .B1(new_n1114), .B2(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT114), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n778), .ZN(new_n1121));
  OAI221_X1 g0921(.A(new_n1103), .B1(new_n833), .B2(new_n971), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1100), .A2(new_n1101), .A3(new_n1122), .ZN(G390));
  AOI21_X1  g0923(.A(new_n851), .B1(new_n765), .B2(new_n860), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n955), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n946), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1126), .A2(new_n950), .A3(new_n949), .ZN(new_n1127));
  AOI21_X1  g0927(.A(KEYINPUT38), .B1(new_n920), .B2(new_n921), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n851), .B1(new_n771), .B2(new_n860), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n946), .B1(new_n1128), .B2(new_n936), .C1(new_n1129), .C2(new_n1125), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1127), .A2(new_n1130), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n748), .A2(G330), .A3(new_n860), .A4(new_n955), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1132), .A2(KEYINPUT115), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1133), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1127), .A2(new_n1130), .A3(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n750), .A2(new_n512), .ZN(new_n1138));
  AND3_X1   g0938(.A1(new_n959), .A2(new_n667), .A3(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n748), .A2(G330), .A3(new_n860), .ZN(new_n1140));
  AND3_X1   g0940(.A1(new_n1140), .A2(KEYINPUT116), .A3(new_n1125), .ZN(new_n1141));
  AOI21_X1  g0941(.A(KEYINPUT116), .B1(new_n1140), .B2(new_n1125), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1132), .A2(new_n1129), .ZN(new_n1143));
  NOR3_X1   g0943(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1140), .A2(new_n1125), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1124), .B1(new_n1145), .B2(new_n1132), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1139), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n838), .B1(new_n1137), .B2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1148), .B1(new_n1137), .B2(new_n1147), .ZN(new_n1149));
  AND3_X1   g0949(.A1(new_n1127), .A2(new_n1135), .A3(new_n1130), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1135), .B1(new_n1127), .B2(new_n1130), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n843), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n949), .A2(new_n775), .A3(new_n950), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n845), .B1(new_n343), .B2(new_n868), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n829), .A2(new_n262), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1156), .B(KEYINPUT118), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n790), .A2(new_n206), .B1(new_n795), .B2(new_n615), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n818), .A2(G77), .B1(KEYINPUT117), .B2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1159), .B1(KEYINPUT117), .B2(new_n1158), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n802), .A2(G283), .B1(new_n885), .B2(G116), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n881), .B(new_n1161), .C1(new_n871), .C2(new_n807), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n808), .A2(G125), .B1(new_n813), .B2(G50), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(KEYINPUT54), .B(G143), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n795), .A2(new_n1165), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n262), .B(new_n1166), .C1(G132), .C2(new_n885), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n1068), .A2(G137), .B1(new_n802), .B2(G128), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1164), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(G159), .B2(new_n818), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n814), .A2(new_n339), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1171), .B(KEYINPUT53), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n1157), .A2(new_n1163), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1154), .B(new_n1155), .C1(new_n1121), .C2(new_n1173), .ZN(new_n1174));
  AND2_X1   g0974(.A1(new_n1153), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1149), .A2(new_n1175), .ZN(G378));
  AND3_X1   g0976(.A1(new_n934), .A2(G330), .A3(new_n940), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n946), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT39), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n926), .A2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1181), .A2(new_n1128), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n925), .A2(new_n921), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(new_n923), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1180), .B1(new_n1184), .B2(new_n926), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1179), .B1(new_n1182), .B2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1125), .B1(new_n854), .B2(new_n861), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1184), .A2(new_n926), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n952), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n917), .A2(new_n348), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n666), .B2(new_n386), .ZN(new_n1194));
  AND3_X1   g0994(.A1(new_n377), .A2(new_n382), .A3(KEYINPUT86), .ZN(new_n1195));
  AOI21_X1  g0995(.A(KEYINPUT86), .B1(new_n377), .B2(new_n382), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n386), .B(new_n1193), .C1(new_n1195), .C2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1191), .B1(new_n1194), .B2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n386), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(new_n1192), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1201), .A2(new_n1197), .A3(new_n1190), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1199), .A2(new_n1202), .ZN(new_n1203));
  AND3_X1   g1003(.A1(new_n1186), .A2(new_n1189), .A3(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1203), .B1(new_n1186), .B2(new_n1189), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1178), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  AND3_X1   g1006(.A1(new_n1201), .A2(new_n1197), .A3(new_n1190), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1190), .B1(new_n1201), .B2(new_n1197), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n951), .B2(new_n957), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1186), .A2(new_n1189), .A3(new_n1203), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1210), .A2(new_n1211), .A3(new_n1177), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n840), .B1(new_n1206), .B2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1209), .A2(new_n775), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n865), .B1(G50), .B2(new_n869), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(G58), .A2(new_n813), .B1(new_n815), .B2(G77), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n363), .B(new_n262), .C1(new_n799), .C2(new_n206), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n790), .A2(new_n205), .B1(new_n801), .B2(new_n291), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n1218), .B(new_n1219), .C1(new_n612), .C2(new_n826), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n808), .A2(G283), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1048), .A2(new_n1217), .A3(new_n1220), .A4(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT58), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n262), .A2(new_n363), .ZN(new_n1224));
  AOI21_X1  g1024(.A(G50), .B1(new_n257), .B2(new_n363), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n1222), .A2(new_n1223), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(G132), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n790), .A2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(G128), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n799), .A2(new_n1229), .B1(new_n795), .B2(new_n887), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n1228), .B(new_n1230), .C1(G125), .C2(new_n802), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1231), .B1(new_n339), .B2(new_n817), .C1(new_n814), .C2(new_n1165), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(KEYINPUT59), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n813), .A2(G159), .ZN(new_n1234));
  AOI211_X1 g1034(.A(G33), .B(G41), .C1(new_n808), .C2(G124), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1233), .A2(new_n1234), .A3(new_n1235), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1232), .A2(KEYINPUT59), .ZN(new_n1237));
  OAI221_X1 g1037(.A(new_n1226), .B1(new_n1223), .B2(new_n1222), .C1(new_n1236), .C2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1216), .B1(new_n1238), .B2(new_n778), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1215), .A2(new_n1239), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n1240), .B(KEYINPUT119), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1214), .A2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  AND3_X1   g1043(.A1(new_n1210), .A2(new_n1177), .A3(new_n1211), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1177), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1245));
  OAI21_X1  g1045(.A(KEYINPUT57), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1139), .ZN(new_n1247));
  OR2_X1    g1047(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1247), .B1(new_n1152), .B2(new_n1248), .ZN(new_n1249));
  OAI211_X1 g1049(.A(KEYINPUT120), .B(new_n726), .C1(new_n1246), .C2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT57), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1251), .B1(new_n1252), .B2(new_n1249), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1250), .A2(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1139), .B1(new_n1137), .B2(new_n1147), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1206), .A2(new_n1212), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1255), .A2(new_n1256), .A3(KEYINPUT57), .ZN(new_n1257));
  AOI21_X1  g1057(.A(KEYINPUT120), .B1(new_n1257), .B2(new_n726), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1243), .B1(new_n1254), .B2(new_n1258), .ZN(G375));
  NOR2_X1   g1059(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(new_n1247), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n990), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1261), .A2(new_n1262), .A3(new_n1147), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1125), .A2(new_n775), .ZN(new_n1264));
  XNOR2_X1  g1064(.A(new_n1264), .B(KEYINPUT121), .ZN(new_n1265));
  OAI221_X1 g1065(.A(new_n1044), .B1(new_n205), .B2(new_n814), .C1(new_n1064), .C2(new_n807), .ZN(new_n1266));
  OAI221_X1 g1066(.A(new_n262), .B1(new_n795), .B2(new_n206), .C1(new_n876), .C2(new_n799), .ZN(new_n1267));
  OAI22_X1  g1067(.A1(new_n790), .A2(new_n291), .B1(new_n801), .B2(new_n871), .ZN(new_n1268));
  NOR4_X1   g1068(.A1(new_n1266), .A2(new_n1081), .A3(new_n1267), .A4(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(KEYINPUT122), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(new_n808), .A2(G128), .B1(new_n813), .B2(G58), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n818), .A2(G50), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n260), .B1(new_n795), .B2(new_n339), .ZN(new_n1274));
  OAI22_X1  g1074(.A1(new_n1227), .A2(new_n801), .B1(new_n790), .B2(new_n1165), .ZN(new_n1275));
  AOI211_X1 g1075(.A(new_n1274), .B(new_n1275), .C1(G137), .C2(new_n885), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n815), .A2(G159), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1272), .A2(new_n1273), .A3(new_n1276), .A4(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1271), .A2(new_n1278), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1270), .A2(KEYINPUT122), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n778), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n845), .B1(new_n455), .B2(new_n868), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1265), .A2(new_n1281), .A3(new_n1282), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1283), .B1(new_n1260), .B2(new_n840), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1263), .A2(new_n1285), .ZN(new_n1286));
  XOR2_X1   g1086(.A(new_n1286), .B(KEYINPUT123), .Z(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(G381));
  NOR2_X1   g1088(.A1(G396), .A2(G393), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1290), .A2(G384), .ZN(new_n1291));
  INV_X1    g1091(.A(G378), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1287), .A2(new_n1291), .A3(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(G390), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1026), .A2(new_n1059), .A3(new_n1294), .ZN(new_n1295));
  NOR3_X1   g1095(.A1(new_n1293), .A2(new_n1295), .A3(G375), .ZN(new_n1296));
  XOR2_X1   g1096(.A(new_n1296), .B(KEYINPUT124), .Z(G407));
  OR2_X1    g1097(.A1(G378), .A2(G343), .ZN(new_n1298));
  OAI211_X1 g1098(.A(G407), .B(G213), .C1(G375), .C2(new_n1298), .ZN(G409));
  NAND2_X1  g1099(.A1(G396), .A2(G393), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1290), .A2(KEYINPUT126), .A3(new_n1300), .ZN(new_n1301));
  AND3_X1   g1101(.A1(new_n1026), .A2(new_n1059), .A3(new_n1294), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1294), .B1(new_n1026), .B2(new_n1059), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1301), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(G387), .A2(G390), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT126), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1300), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1306), .B1(new_n1307), .B2(new_n1289), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(new_n1301), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1305), .A2(new_n1295), .A3(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1304), .A2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(G213), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1313), .A2(G343), .ZN(new_n1314));
  OAI211_X1 g1114(.A(G378), .B(new_n1243), .C1(new_n1254), .C2(new_n1258), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1240), .ZN(new_n1316));
  OAI21_X1  g1116(.A(KEYINPUT125), .B1(new_n1213), .B2(new_n1316), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1255), .A2(new_n1256), .A3(new_n1262), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  NOR3_X1   g1119(.A1(new_n1213), .A2(KEYINPUT125), .A3(new_n1316), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1292), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1314), .B1(new_n1315), .B2(new_n1321), .ZN(new_n1322));
  XNOR2_X1  g1122(.A(new_n1261), .B(KEYINPUT60), .ZN(new_n1323));
  AND2_X1   g1123(.A1(new_n1147), .A2(new_n726), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1325), .A2(G384), .A3(new_n1285), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1326), .ZN(new_n1327));
  AOI21_X1  g1127(.A(G384), .B1(new_n1325), .B2(new_n1285), .ZN(new_n1328));
  NOR2_X1   g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  AOI21_X1  g1129(.A(KEYINPUT62), .B1(new_n1322), .B2(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1315), .A2(new_n1321), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1314), .ZN(new_n1332));
  AOI21_X1  g1132(.A(KEYINPUT127), .B1(new_n1331), .B2(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT127), .ZN(new_n1334));
  AOI211_X1 g1134(.A(new_n1334), .B(new_n1314), .C1(new_n1315), .C2(new_n1321), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1333), .A2(new_n1335), .ZN(new_n1336));
  AND2_X1   g1136(.A1(new_n1329), .A2(KEYINPUT62), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1330), .B1(new_n1336), .B2(new_n1337), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1328), .ZN(new_n1339));
  NAND4_X1  g1139(.A1(new_n1339), .A2(G2897), .A3(new_n1314), .A4(new_n1326), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1314), .A2(G2897), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1341), .B1(new_n1327), .B2(new_n1328), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1340), .A2(new_n1342), .ZN(new_n1343));
  OAI21_X1  g1143(.A(new_n1343), .B1(new_n1333), .B2(new_n1335), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT61), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1344), .A2(new_n1345), .ZN(new_n1346));
  OAI21_X1  g1146(.A(new_n1312), .B1(new_n1338), .B2(new_n1346), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1336), .A2(KEYINPUT63), .A3(new_n1329), .ZN(new_n1348));
  INV_X1    g1148(.A(KEYINPUT63), .ZN(new_n1349));
  INV_X1    g1149(.A(new_n1322), .ZN(new_n1350));
  INV_X1    g1150(.A(new_n1329), .ZN(new_n1351));
  OAI21_X1  g1151(.A(new_n1349), .B1(new_n1350), .B2(new_n1351), .ZN(new_n1352));
  AOI21_X1  g1152(.A(KEYINPUT61), .B1(new_n1343), .B2(new_n1350), .ZN(new_n1353));
  NAND4_X1  g1153(.A1(new_n1348), .A2(new_n1311), .A3(new_n1352), .A4(new_n1353), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1347), .A2(new_n1354), .ZN(G405));
  NAND3_X1  g1155(.A1(new_n1304), .A2(new_n1310), .A3(new_n1351), .ZN(new_n1356));
  INV_X1    g1156(.A(new_n1356), .ZN(new_n1357));
  AOI21_X1  g1157(.A(new_n1351), .B1(new_n1304), .B2(new_n1310), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(G375), .A2(new_n1292), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1359), .A2(new_n1315), .ZN(new_n1360));
  NOR3_X1   g1160(.A1(new_n1357), .A2(new_n1358), .A3(new_n1360), .ZN(new_n1361));
  INV_X1    g1161(.A(new_n1360), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1311), .A2(new_n1329), .ZN(new_n1363));
  AOI21_X1  g1163(.A(new_n1362), .B1(new_n1363), .B2(new_n1356), .ZN(new_n1364));
  NOR2_X1   g1164(.A1(new_n1361), .A2(new_n1364), .ZN(G402));
endmodule


