//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 1 0 1 1 1 0 1 1 1 0 1 0 0 1 0 0 1 1 1 0 1 1 0 1 1 0 0 0 1 1 0 0 1 0 1 1 1 0 1 1 1 0 1 0 1 1 1 0 1 1 0 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:18 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n557,
    new_n558, new_n559, new_n560, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n580, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n623,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT64), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT65), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n453), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  AND2_X1   g035(.A1(KEYINPUT66), .A2(G2105), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT66), .A2(G2105), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n468));
  AND3_X1   g043(.A1(new_n466), .A2(new_n468), .A3(G125), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT67), .ZN(new_n470));
  INV_X1    g045(.A(G113), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n470), .B1(new_n471), .B2(new_n467), .ZN(new_n472));
  NAND3_X1  g047(.A1(KEYINPUT67), .A2(G113), .A3(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n464), .B1(new_n469), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n465), .A2(KEYINPUT68), .A3(G2104), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n476), .A2(new_n468), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT68), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n478), .B1(new_n467), .B2(KEYINPUT3), .ZN(new_n479));
  NAND4_X1  g054(.A1(new_n477), .A2(G137), .A3(new_n479), .A4(new_n463), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n467), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G101), .ZN(new_n482));
  AND3_X1   g057(.A1(new_n475), .A2(new_n480), .A3(new_n482), .ZN(G160));
  OAI21_X1  g058(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(G112), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n484), .B1(new_n464), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n479), .A2(new_n468), .A3(new_n476), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n487), .A2(new_n463), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n486), .B1(new_n488), .B2(G124), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n487), .A2(G2105), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G136), .ZN(new_n491));
  AND2_X1   g066(.A1(new_n489), .A2(new_n491), .ZN(G162));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT66), .ZN(new_n494));
  INV_X1    g069(.A(G2105), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(KEYINPUT66), .A2(G2105), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n496), .A2(G138), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n466), .A2(new_n468), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n493), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n481), .A2(G102), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n463), .A2(KEYINPUT4), .A3(G138), .ZN(new_n502));
  OAI211_X1 g077(.A(new_n500), .B(new_n501), .C1(new_n487), .C2(new_n502), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n479), .A2(new_n476), .A3(G126), .A4(new_n468), .ZN(new_n504));
  NAND2_X1  g079(.A1(G114), .A2(G2104), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n495), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n503), .A2(new_n506), .ZN(G164));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT5), .B(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G62), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT70), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n510), .A2(new_n511), .B1(G75), .B2(G543), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n509), .A2(KEYINPUT70), .A3(G62), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n508), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n508), .A2(KEYINPUT6), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT6), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G651), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  AND2_X1   g093(.A1(G50), .A2(G543), .ZN(new_n519));
  AND3_X1   g094(.A1(new_n518), .A2(KEYINPUT69), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g095(.A(KEYINPUT69), .B1(new_n518), .B2(new_n519), .ZN(new_n521));
  INV_X1    g096(.A(G88), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n509), .A2(new_n515), .A3(new_n517), .ZN(new_n523));
  OAI22_X1  g098(.A1(new_n520), .A2(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n514), .A2(new_n524), .ZN(G166));
  NAND3_X1  g100(.A1(new_n509), .A2(G63), .A3(G651), .ZN(new_n526));
  AND3_X1   g101(.A1(new_n515), .A2(new_n517), .A3(G543), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(G51), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n526), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT7), .ZN(new_n532));
  INV_X1    g107(.A(G89), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n523), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n530), .A2(new_n534), .ZN(G168));
  AOI22_X1  g110(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n536), .A2(new_n508), .ZN(new_n537));
  INV_X1    g112(.A(new_n523), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G90), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT71), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n527), .A2(G52), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n537), .A2(new_n539), .A3(new_n540), .A4(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(G90), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n541), .B1(new_n543), .B2(new_n523), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n536), .A2(new_n508), .ZN(new_n545));
  OAI21_X1  g120(.A(KEYINPUT71), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n542), .A2(new_n546), .ZN(G171));
  NAND2_X1  g122(.A1(new_n527), .A2(G43), .ZN(new_n548));
  INV_X1    g123(.A(G81), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n549), .B2(new_n523), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n509), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n551), .A2(new_n508), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT72), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT73), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT74), .ZN(G188));
  INV_X1    g136(.A(KEYINPUT75), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G53), .ZN(new_n563));
  OAI21_X1  g138(.A(KEYINPUT9), .B1(new_n528), .B2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT9), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n527), .A2(new_n562), .A3(new_n565), .A4(G53), .ZN(new_n566));
  INV_X1    g141(.A(G91), .ZN(new_n567));
  OAI21_X1  g142(.A(KEYINPUT76), .B1(new_n523), .B2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT76), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n518), .A2(new_n569), .A3(G91), .A4(new_n509), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n564), .A2(new_n566), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n509), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n572));
  OR2_X1    g147(.A1(new_n572), .A2(KEYINPUT77), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(KEYINPUT77), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n573), .A2(G651), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n571), .A2(new_n575), .ZN(G299));
  INV_X1    g151(.A(G171), .ZN(G301));
  INV_X1    g152(.A(G168), .ZN(G286));
  INV_X1    g153(.A(G166), .ZN(G303));
  NAND2_X1  g154(.A1(new_n527), .A2(G49), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n582), .B1(G87), .B2(new_n538), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G288));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  XOR2_X1   g160(.A(KEYINPUT5), .B(G543), .Z(new_n586));
  INV_X1    g161(.A(G61), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n588), .A2(KEYINPUT78), .A3(G651), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT78), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n509), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n591), .B2(new_n508), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT79), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n589), .A2(new_n592), .A3(KEYINPUT79), .ZN(new_n596));
  NAND4_X1  g171(.A1(new_n515), .A2(new_n517), .A3(G48), .A4(G543), .ZN(new_n597));
  INV_X1    g172(.A(G86), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n523), .B2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n595), .A2(new_n596), .A3(new_n600), .ZN(G305));
  XOR2_X1   g176(.A(KEYINPUT80), .B(G47), .Z(new_n602));
  INV_X1    g177(.A(G85), .ZN(new_n603));
  OAI22_X1  g178(.A1(new_n528), .A2(new_n602), .B1(new_n523), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n605), .A2(new_n508), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(G290));
  NAND3_X1  g183(.A1(new_n538), .A2(KEYINPUT10), .A3(G92), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT10), .ZN(new_n610));
  INV_X1    g185(.A(G92), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n523), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(G79), .A2(G543), .ZN(new_n614));
  INV_X1    g189(.A(G66), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n586), .B2(new_n615), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n616), .A2(G651), .B1(G54), .B2(new_n527), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n618), .A2(G868), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n619), .B1(G868), .B2(G171), .ZN(G284));
  AOI21_X1  g195(.A(new_n619), .B1(G868), .B2(G171), .ZN(G321));
  NAND2_X1  g196(.A1(G286), .A2(G868), .ZN(new_n622));
  AND2_X1   g197(.A1(new_n571), .A2(new_n575), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(G868), .ZN(G297));
  OAI21_X1  g199(.A(new_n622), .B1(new_n623), .B2(G868), .ZN(G280));
  INV_X1    g200(.A(new_n618), .ZN(new_n626));
  INV_X1    g201(.A(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(G860), .ZN(G148));
  OR2_X1    g203(.A1(new_n550), .A2(new_n552), .ZN(new_n629));
  INV_X1    g204(.A(G868), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g206(.A1(new_n618), .A2(G559), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n631), .B1(new_n632), .B2(new_n630), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(KEYINPUT81), .Z(G323));
  XNOR2_X1  g209(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g210(.A(KEYINPUT3), .B(G2104), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(new_n481), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(KEYINPUT12), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT13), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2100), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n488), .A2(G123), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(KEYINPUT82), .Z(new_n642));
  OAI21_X1  g217(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n643));
  INV_X1    g218(.A(G111), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n643), .B1(new_n464), .B2(new_n644), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n645), .B1(new_n490), .B2(G135), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(G2096), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n640), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n650), .B1(new_n649), .B2(new_n648), .ZN(G156));
  XNOR2_X1  g226(.A(G2451), .B(G2454), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT16), .ZN(new_n653));
  XOR2_X1   g228(.A(G2443), .B(G2446), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT83), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n655), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2427), .B(G2438), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2430), .ZN(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT15), .B(G2435), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n660), .A2(new_n661), .ZN(new_n663));
  AND3_X1   g238(.A1(new_n662), .A2(new_n663), .A3(KEYINPUT14), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n658), .A2(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(G14), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n666), .B1(new_n658), .B2(new_n664), .ZN(new_n667));
  AND2_X1   g242(.A1(new_n665), .A2(new_n667), .ZN(G401));
  XOR2_X1   g243(.A(G2084), .B(G2090), .Z(new_n669));
  XNOR2_X1  g244(.A(G2067), .B(G2678), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2072), .B(G2078), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT18), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n671), .B(KEYINPUT17), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n670), .B(KEYINPUT84), .ZN(new_n675));
  AND2_X1   g250(.A1(new_n675), .A2(new_n669), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n673), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(new_n671), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n669), .B1(new_n675), .B2(new_n678), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n679), .B1(new_n675), .B2(new_n674), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n677), .A2(KEYINPUT85), .A3(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  AOI21_X1  g257(.A(KEYINPUT85), .B1(new_n677), .B2(new_n680), .ZN(new_n683));
  OAI21_X1  g258(.A(G2096), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(new_n683), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n685), .A2(new_n649), .A3(new_n681), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(G2100), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n684), .A2(new_n686), .A3(G2100), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(G227));
  INV_X1    g267(.A(G1986), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1971), .B(G1976), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT19), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(G1956), .B(G2474), .Z(new_n697));
  XOR2_X1   g272(.A(G1961), .B(G1966), .Z(new_n698));
  AND2_X1   g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT20), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n697), .A2(new_n698), .ZN(new_n702));
  NOR3_X1   g277(.A1(new_n696), .A2(new_n699), .A3(new_n702), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(new_n696), .B2(new_n702), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n693), .B1(new_n701), .B2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n701), .A2(new_n704), .A3(new_n693), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n706), .A2(new_n707), .A3(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(new_n707), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n708), .B1(new_n711), .B2(new_n705), .ZN(new_n712));
  XNOR2_X1  g287(.A(G1991), .B(G1996), .ZN(new_n713));
  INV_X1    g288(.A(G1981), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n710), .A2(new_n712), .A3(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n715), .B1(new_n710), .B2(new_n712), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n717), .A2(new_n718), .ZN(G229));
  INV_X1    g294(.A(G29), .ZN(new_n720));
  NOR2_X1   g295(.A1(G160), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n720), .B1(KEYINPUT24), .B2(G34), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(KEYINPUT24), .B2(G34), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G2084), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT93), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n720), .A2(G32), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n490), .A2(G141), .ZN(new_n729));
  NAND3_X1  g304(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT26), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n730), .A2(new_n731), .ZN(new_n733));
  AOI22_X1  g308(.A1(new_n732), .A2(new_n733), .B1(G105), .B2(new_n481), .ZN(new_n734));
  INV_X1    g309(.A(new_n488), .ZN(new_n735));
  INV_X1    g310(.A(G129), .ZN(new_n736));
  OAI211_X1 g311(.A(new_n729), .B(new_n734), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n728), .B1(new_n738), .B2(new_n720), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT90), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT27), .B(G1996), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(G16), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(G5), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G171), .B2(new_n744), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n727), .B(new_n743), .C1(G1961), .C2(new_n746), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT94), .ZN(new_n748));
  NOR2_X1   g323(.A1(G168), .A2(new_n744), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(new_n744), .B2(G21), .ZN(new_n750));
  INV_X1    g325(.A(G1966), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(KEYINPUT92), .ZN(new_n753));
  INV_X1    g328(.A(G2072), .ZN(new_n754));
  AND2_X1   g329(.A1(new_n720), .A2(G33), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT25), .Z(new_n757));
  NAND2_X1  g332(.A1(new_n490), .A2(G139), .ZN(new_n758));
  AOI22_X1  g333(.A1(new_n636), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n759), .A2(new_n463), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n757), .A2(new_n758), .A3(new_n760), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n755), .B1(new_n761), .B2(G29), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n753), .B1(new_n754), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n754), .B2(new_n762), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n744), .A2(G4), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(new_n626), .B2(new_n744), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G1348), .ZN(new_n767));
  OAI22_X1  g342(.A1(new_n752), .A2(KEYINPUT92), .B1(new_n720), .B2(new_n647), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n724), .A2(new_n725), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT89), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n720), .A2(G26), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT28), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n490), .A2(G140), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n488), .A2(G128), .ZN(new_n775));
  OR2_X1    g350(.A1(G104), .A2(G2105), .ZN(new_n776));
  OAI211_X1 g351(.A(G2104), .B(new_n776), .C1(new_n463), .C2(G116), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n777), .A2(KEYINPUT88), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n777), .A2(KEYINPUT88), .ZN(new_n779));
  OAI211_X1 g354(.A(new_n774), .B(new_n775), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n773), .B1(new_n781), .B2(new_n720), .ZN(new_n782));
  INV_X1    g357(.A(G2067), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n764), .A2(new_n769), .A3(new_n771), .A4(new_n784), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT29), .B(G2090), .Z(new_n786));
  INV_X1    g361(.A(G162), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n787), .A2(G29), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n720), .A2(G35), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT95), .Z(new_n790));
  AOI21_X1  g365(.A(new_n786), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(G2078), .ZN(new_n792));
  NAND2_X1  g367(.A1(G164), .A2(G29), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G27), .B2(G29), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n791), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n788), .A2(new_n790), .A3(new_n786), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT31), .B(G11), .ZN(new_n797));
  INV_X1    g372(.A(G28), .ZN(new_n798));
  AOI21_X1  g373(.A(G29), .B1(new_n798), .B2(KEYINPUT30), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT91), .ZN(new_n800));
  OAI22_X1  g375(.A1(new_n799), .A2(new_n800), .B1(KEYINPUT30), .B2(new_n798), .ZN(new_n801));
  AND2_X1   g376(.A1(new_n799), .A2(new_n800), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n797), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(new_n750), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n803), .B1(new_n804), .B2(G1966), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n744), .A2(G19), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(new_n553), .B2(new_n744), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(G1341), .Z(new_n808));
  NAND4_X1  g383(.A1(new_n795), .A2(new_n796), .A3(new_n805), .A4(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n744), .A2(G20), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT23), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n623), .B2(new_n744), .ZN(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT96), .B(G1956), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n794), .A2(new_n792), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n812), .A2(new_n814), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n746), .A2(G1961), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n815), .A2(new_n816), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n809), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(new_n742), .B2(new_n740), .ZN(new_n821));
  NOR3_X1   g396(.A1(new_n748), .A2(new_n785), .A3(new_n821), .ZN(new_n822));
  AND2_X1   g397(.A1(new_n744), .A2(G6), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(G305), .B2(G16), .ZN(new_n824));
  XNOR2_X1  g399(.A(KEYINPUT32), .B(G1981), .ZN(new_n825));
  INV_X1    g400(.A(new_n825), .ZN(new_n826));
  OR2_X1    g401(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n744), .A2(G22), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(G166), .B2(new_n744), .ZN(new_n829));
  INV_X1    g404(.A(G1971), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n824), .A2(new_n826), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n744), .A2(G23), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(new_n583), .B2(new_n744), .ZN(new_n834));
  XNOR2_X1  g409(.A(KEYINPUT33), .B(G1976), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  NAND4_X1  g411(.A1(new_n827), .A2(new_n831), .A3(new_n832), .A4(new_n836), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n837), .A2(KEYINPUT34), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(KEYINPUT34), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n490), .A2(G131), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n488), .A2(G119), .ZN(new_n841));
  OAI221_X1 g416(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n463), .C2(G107), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n843), .A2(KEYINPUT86), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT86), .ZN(new_n845));
  NAND4_X1  g420(.A1(new_n840), .A2(new_n841), .A3(new_n845), .A4(new_n842), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(G29), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n849), .B1(G25), .B2(G29), .ZN(new_n850));
  XOR2_X1   g425(.A(KEYINPUT35), .B(G1991), .Z(new_n851));
  AND2_X1   g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n850), .A2(new_n851), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n744), .A2(G24), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n854), .B1(new_n607), .B2(new_n744), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(G1986), .ZN(new_n856));
  NOR3_X1   g431(.A1(new_n852), .A2(new_n853), .A3(new_n856), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n838), .A2(new_n839), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(KEYINPUT87), .A2(KEYINPUT36), .ZN(new_n859));
  OR2_X1    g434(.A1(KEYINPUT87), .A2(KEYINPUT36), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  OAI211_X1 g436(.A(new_n822), .B(new_n861), .C1(new_n858), .C2(new_n859), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT97), .ZN(G311));
  XNOR2_X1  g438(.A(new_n862), .B(KEYINPUT98), .ZN(G150));
  AOI22_X1  g439(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n865), .A2(new_n508), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n527), .A2(G55), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n538), .A2(G93), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n629), .A2(KEYINPUT99), .A3(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT99), .ZN(new_n871));
  NAND4_X1  g446(.A1(new_n866), .A2(new_n871), .A3(new_n867), .A4(new_n868), .ZN(new_n872));
  INV_X1    g447(.A(G93), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n867), .B1(new_n873), .B2(new_n523), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n865), .A2(new_n508), .ZN(new_n875));
  OAI21_X1  g450(.A(KEYINPUT99), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n872), .A2(new_n876), .A3(new_n553), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n870), .A2(new_n877), .ZN(new_n878));
  XOR2_X1   g453(.A(new_n878), .B(KEYINPUT38), .Z(new_n879));
  NAND2_X1  g454(.A1(new_n626), .A2(G559), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n879), .B(new_n880), .ZN(new_n881));
  AND2_X1   g456(.A1(new_n881), .A2(KEYINPUT39), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n881), .A2(KEYINPUT39), .ZN(new_n883));
  NOR3_X1   g458(.A1(new_n882), .A2(new_n883), .A3(G860), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n869), .A2(G860), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(KEYINPUT37), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n884), .A2(new_n886), .ZN(G145));
  NAND2_X1  g462(.A1(new_n490), .A2(G142), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT100), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n490), .A2(KEYINPUT100), .A3(G142), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n638), .ZN(new_n893));
  OAI21_X1  g468(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n894));
  INV_X1    g469(.A(G118), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n894), .B1(new_n464), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n896), .B1(new_n488), .B2(G130), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n892), .A2(new_n893), .A3(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n893), .B1(new_n892), .B2(new_n897), .ZN(new_n900));
  NOR3_X1   g475(.A1(new_n899), .A2(new_n900), .A3(new_n847), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n847), .B1(new_n899), .B2(new_n900), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n902), .A2(KEYINPUT101), .A3(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT101), .ZN(new_n905));
  INV_X1    g480(.A(new_n900), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n848), .B1(new_n906), .B2(new_n898), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n905), .B1(new_n907), .B2(new_n901), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n504), .A2(new_n505), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(G2105), .ZN(new_n910));
  INV_X1    g485(.A(new_n501), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n463), .A2(new_n636), .A3(G138), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n911), .B1(new_n912), .B2(new_n493), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n498), .A2(new_n493), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n914), .A2(new_n479), .A3(new_n477), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n910), .A2(new_n913), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n781), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n780), .A2(G164), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n761), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n917), .A2(new_n918), .A3(new_n761), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n737), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n917), .A2(new_n918), .A3(new_n761), .ZN(new_n923));
  NOR3_X1   g498(.A1(new_n923), .A2(new_n919), .A3(new_n738), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n904), .B(new_n908), .C1(new_n922), .C2(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(KEYINPUT101), .B1(new_n902), .B2(new_n903), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n920), .A2(new_n737), .A3(new_n921), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n738), .B1(new_n923), .B2(new_n919), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n647), .B(G160), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n930), .B(G162), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n925), .A2(new_n929), .A3(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(G37), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n925), .A2(new_n929), .ZN(new_n935));
  INV_X1    g510(.A(new_n931), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n938), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g514(.A(G299), .B(new_n618), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT41), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(KEYINPUT102), .B1(new_n623), .B2(new_n618), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n626), .A2(G299), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n618), .A2(new_n575), .A3(new_n571), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n943), .B1(new_n946), .B2(KEYINPUT102), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n942), .B1(new_n941), .B2(new_n947), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n878), .B(new_n632), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OR2_X1    g525(.A1(new_n950), .A2(KEYINPUT103), .ZN(new_n951));
  OR2_X1    g526(.A1(new_n949), .A2(new_n940), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n950), .A2(KEYINPUT103), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  OR2_X1    g529(.A1(new_n954), .A2(KEYINPUT42), .ZN(new_n955));
  XNOR2_X1  g530(.A(G305), .B(G166), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT105), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OR2_X1    g533(.A1(new_n583), .A2(KEYINPUT104), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n583), .A2(KEYINPUT104), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(new_n607), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n959), .A2(G290), .A3(new_n960), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AND2_X1   g539(.A1(G305), .A2(G303), .ZN(new_n965));
  NOR2_X1   g540(.A1(G305), .A2(G303), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT105), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n958), .A2(new_n964), .A3(new_n967), .ZN(new_n968));
  OR2_X1    g543(.A1(new_n967), .A2(new_n964), .ZN(new_n969));
  AND2_X1   g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n954), .A2(KEYINPUT42), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n955), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n970), .B1(new_n955), .B2(new_n971), .ZN(new_n973));
  OAI21_X1  g548(.A(G868), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n869), .A2(new_n630), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(G295));
  NAND2_X1  g551(.A1(new_n974), .A2(new_n975), .ZN(G331));
  NAND3_X1  g552(.A1(G286), .A2(new_n542), .A3(new_n546), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(G286), .B1(new_n542), .B2(new_n546), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n878), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(G171), .A2(G168), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n982), .A2(new_n870), .A3(new_n877), .A4(new_n978), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n981), .A2(new_n946), .A3(new_n983), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n984), .A2(KEYINPUT106), .ZN(new_n985));
  AND2_X1   g560(.A1(new_n984), .A2(KEYINPUT106), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT102), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n987), .B1(new_n626), .B2(G299), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n941), .B(new_n988), .C1(new_n940), .C2(new_n987), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n946), .A2(KEYINPUT41), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n981), .A2(new_n983), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n985), .B1(new_n986), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n968), .A2(new_n969), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n933), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT43), .ZN(new_n996));
  OAI211_X1 g571(.A(KEYINPUT41), .B(new_n988), .C1(new_n940), .C2(new_n987), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT107), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n947), .A2(KEYINPUT107), .A3(KEYINPUT41), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n999), .A2(new_n991), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n946), .A2(new_n941), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n984), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(new_n994), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  NOR3_X1   g581(.A1(new_n995), .A2(new_n996), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n995), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n986), .A2(new_n992), .ZN(new_n1009));
  INV_X1    g584(.A(new_n985), .ZN(new_n1010));
  AND3_X1   g585(.A1(new_n1009), .A2(new_n994), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(KEYINPUT43), .B1(new_n1008), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT44), .B1(new_n1007), .B2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(KEYINPUT43), .B1(new_n995), .B2(new_n1011), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n984), .A2(KEYINPUT106), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1016), .B1(new_n948), .B2(new_n991), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n970), .B1(new_n1017), .B2(new_n985), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1005), .A2(new_n1018), .A3(new_n996), .A4(new_n933), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1015), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1014), .B1(KEYINPUT44), .B2(new_n1021), .ZN(G397));
  INV_X1    g597(.A(KEYINPUT123), .ZN(new_n1023));
  INV_X1    g598(.A(G1384), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1024), .B1(new_n503), .B2(new_n506), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT45), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n475), .A2(new_n480), .A3(G40), .A4(new_n482), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1026), .A2(G1384), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1028), .B1(new_n916), .B2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1027), .A2(new_n1030), .A3(new_n792), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  XOR2_X1   g607(.A(KEYINPUT121), .B(KEYINPUT53), .Z(new_n1033));
  NOR2_X1   g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1025), .A2(KEYINPUT50), .ZN(new_n1036));
  NOR2_X1   g611(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1028), .B1(new_n916), .B2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(G1961), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT53), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1040), .B1(new_n1031), .B2(KEYINPUT119), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT119), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1027), .A2(new_n1030), .A3(new_n1042), .A4(new_n792), .ZN(new_n1043));
  AOI211_X1 g618(.A(KEYINPUT120), .B(new_n1039), .C1(new_n1041), .C2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT120), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1031), .A2(KEYINPUT119), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1046), .A2(KEYINPUT53), .A3(new_n1043), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1039), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1045), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1035), .B1(new_n1044), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT122), .ZN(new_n1051));
  AND3_X1   g626(.A1(new_n1050), .A2(new_n1051), .A3(G171), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1051), .B1(new_n1050), .B2(G171), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT51), .ZN(new_n1055));
  INV_X1    g630(.A(G8), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(new_n751), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1036), .A2(new_n1038), .A3(new_n725), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1056), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(G286), .A2(G8), .ZN(new_n1061));
  XNOR2_X1  g636(.A(new_n1061), .B(KEYINPUT117), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1055), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1059), .ZN(new_n1064));
  AOI21_X1  g639(.A(G1966), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1065));
  OAI21_X1  g640(.A(G8), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  XOR2_X1   g641(.A(new_n1061), .B(KEYINPUT117), .Z(new_n1067));
  NAND3_X1  g642(.A1(new_n1066), .A2(KEYINPUT51), .A3(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1062), .B1(new_n1065), .B2(new_n1064), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1063), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(KEYINPUT118), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT62), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT118), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1063), .A2(new_n1068), .A3(new_n1073), .A4(new_n1069), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1071), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n600), .A2(new_n589), .A3(new_n592), .ZN(new_n1076));
  AOI21_X1  g651(.A(KEYINPUT109), .B1(new_n1076), .B2(G1981), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n595), .A2(new_n714), .A3(new_n596), .A4(new_n600), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1076), .A2(KEYINPUT109), .A3(G1981), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1078), .A2(new_n1079), .A3(KEYINPUT49), .A4(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT111), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  AND3_X1   g658(.A1(new_n1076), .A2(KEYINPUT109), .A3(G1981), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1084), .A2(new_n1077), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1085), .A2(KEYINPUT111), .A3(KEYINPUT49), .A4(new_n1079), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1083), .A2(new_n1086), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1025), .A2(new_n1028), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(G8), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1085), .A2(new_n1079), .ZN(new_n1091));
  XOR2_X1   g666(.A(KEYINPUT110), .B(KEYINPUT49), .Z(new_n1092));
  AOI21_X1  g667(.A(new_n1090), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(G1976), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1089), .A2(G8), .A3(new_n1094), .A4(G288), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT52), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT108), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n583), .A2(G1976), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1098), .B(G8), .C1(new_n1025), .C2(new_n1028), .ZN(new_n1099));
  OAI211_X1 g674(.A(new_n1095), .B(new_n1096), .C1(new_n1097), .C2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1099), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n583), .A2(G1976), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n1101), .B(KEYINPUT108), .C1(KEYINPUT52), .C2(new_n1102), .ZN(new_n1103));
  AOI22_X1  g678(.A1(new_n1087), .A2(new_n1093), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1057), .A2(new_n830), .ZN(new_n1105));
  INV_X1    g680(.A(G2090), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1036), .A2(new_n1038), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(KEYINPUT55), .B1(G166), .B2(new_n1056), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT55), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1110), .B(G8), .C1(new_n514), .C2(new_n524), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  AND3_X1   g687(.A1(new_n1108), .A2(G8), .A3(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1112), .B1(new_n1108), .B2(G8), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  AND2_X1   g690(.A1(new_n1104), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1075), .A2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1023), .B1(new_n1054), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(KEYINPUT120), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1047), .A2(new_n1045), .A3(new_n1048), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1034), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(KEYINPUT122), .B1(new_n1122), .B2(G301), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1050), .A2(new_n1051), .A3(G171), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1125), .A2(KEYINPUT123), .A3(new_n1116), .A4(new_n1075), .ZN(new_n1126));
  AND2_X1   g701(.A1(new_n1070), .A2(KEYINPUT118), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1074), .ZN(new_n1128));
  OAI21_X1  g703(.A(KEYINPUT62), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1118), .A2(new_n1126), .A3(new_n1129), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n1079), .B(KEYINPUT112), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1087), .A2(new_n1093), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n583), .A2(new_n1094), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1131), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1090), .ZN(new_n1135));
  AOI22_X1  g710(.A1(new_n1134), .A2(new_n1135), .B1(new_n1104), .B2(new_n1113), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT113), .ZN(new_n1137));
  OAI21_X1  g712(.A(G168), .B1(new_n1137), .B2(KEYINPUT63), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1066), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1104), .A2(new_n1115), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1137), .A2(KEYINPUT63), .ZN(new_n1141));
  AND2_X1   g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1136), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  AOI211_X1 g719(.A(new_n1039), .B(new_n1034), .C1(KEYINPUT53), .C2(new_n1032), .ZN(new_n1145));
  AOI21_X1  g720(.A(KEYINPUT54), .B1(new_n1145), .B2(G301), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1123), .A2(new_n1124), .A3(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1145), .A2(G171), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n1148), .B(KEYINPUT54), .C1(new_n1122), .C2(G171), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(G1348), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1151));
  NOR3_X1   g726(.A1(new_n1025), .A2(G2067), .A3(new_n1028), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1155));
  INV_X1    g730(.A(G1956), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT57), .ZN(new_n1158));
  NAND2_X1  g733(.A1(G299), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n571), .A2(new_n575), .A3(KEYINPUT57), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  XNOR2_X1  g736(.A(KEYINPUT56), .B(G2072), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1027), .A2(new_n1030), .A3(new_n1162), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1157), .A2(new_n1161), .A3(new_n1163), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1154), .A2(new_n626), .A3(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1163), .ZN(new_n1166));
  AOI21_X1  g741(.A(G1956), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1167));
  OAI211_X1 g742(.A(new_n1159), .B(new_n1160), .C1(new_n1166), .C2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1165), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT61), .ZN(new_n1170));
  AND3_X1   g745(.A1(new_n1157), .A2(new_n1161), .A3(new_n1163), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1161), .B1(new_n1157), .B2(new_n1163), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1170), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1168), .A2(KEYINPUT61), .A3(new_n1164), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(G1996), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1027), .A2(new_n1030), .A3(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT114), .ZN(new_n1178));
  XOR2_X1   g753(.A(KEYINPUT58), .B(G1341), .Z(new_n1179));
  AOI22_X1  g754(.A1(new_n1177), .A2(new_n1178), .B1(new_n1089), .B2(new_n1179), .ZN(new_n1180));
  OR2_X1    g755(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n553), .A2(KEYINPUT115), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1183), .ZN(new_n1184));
  AND3_X1   g759(.A1(new_n1182), .A2(KEYINPUT59), .A3(new_n1184), .ZN(new_n1185));
  AOI21_X1  g760(.A(KEYINPUT59), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1186));
  NOR3_X1   g761(.A1(new_n1175), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT116), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT60), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1189), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1188), .B1(new_n1190), .B2(new_n626), .ZN(new_n1191));
  INV_X1    g766(.A(new_n1191), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1190), .A2(new_n1188), .A3(new_n626), .ZN(new_n1193));
  NAND4_X1  g768(.A1(new_n1192), .A2(KEYINPUT60), .A3(new_n1153), .A4(new_n1193), .ZN(new_n1194));
  INV_X1    g769(.A(new_n1193), .ZN(new_n1195));
  OAI22_X1  g770(.A1(new_n1195), .A2(new_n1191), .B1(new_n1189), .B2(new_n1154), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1169), .B1(new_n1187), .B2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1116), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1199));
  NOR2_X1   g774(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1144), .B1(new_n1150), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1130), .A2(new_n1201), .ZN(new_n1202));
  NOR2_X1   g777(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1203));
  OR2_X1    g778(.A1(new_n848), .A2(new_n851), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n848), .A2(new_n851), .ZN(new_n1205));
  XNOR2_X1  g780(.A(new_n780), .B(new_n783), .ZN(new_n1206));
  XNOR2_X1  g781(.A(new_n737), .B(new_n1176), .ZN(new_n1207));
  NAND4_X1  g782(.A1(new_n1204), .A2(new_n1205), .A3(new_n1206), .A4(new_n1207), .ZN(new_n1208));
  XNOR2_X1  g783(.A(new_n607), .B(new_n693), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n1203), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1202), .A2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1206), .A2(new_n738), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1212), .A2(new_n1203), .ZN(new_n1213));
  NOR3_X1   g788(.A1(new_n1027), .A2(G1996), .A3(new_n1028), .ZN(new_n1214));
  OR2_X1    g789(.A1(new_n1214), .A2(KEYINPUT46), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1214), .A2(KEYINPUT46), .ZN(new_n1216));
  NAND3_X1  g791(.A1(new_n1213), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1217));
  XNOR2_X1  g792(.A(new_n1217), .B(KEYINPUT47), .ZN(new_n1218));
  OR2_X1    g793(.A1(new_n1218), .A2(KEYINPUT124), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n1218), .A2(KEYINPUT124), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1208), .A2(new_n1203), .ZN(new_n1221));
  NAND3_X1  g796(.A1(new_n1203), .A2(new_n693), .A3(new_n607), .ZN(new_n1222));
  XNOR2_X1  g797(.A(new_n1222), .B(KEYINPUT48), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1224));
  OAI22_X1  g799(.A1(new_n1224), .A2(new_n1205), .B1(G2067), .B2(new_n780), .ZN(new_n1225));
  AOI22_X1  g800(.A1(new_n1221), .A2(new_n1223), .B1(new_n1203), .B2(new_n1225), .ZN(new_n1226));
  AND3_X1   g801(.A1(new_n1219), .A2(new_n1220), .A3(new_n1226), .ZN(new_n1227));
  NAND2_X1  g802(.A1(new_n1211), .A2(new_n1227), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g803(.A(KEYINPUT127), .ZN(new_n1230));
  INV_X1    g804(.A(new_n718), .ZN(new_n1231));
  NAND2_X1  g805(.A1(new_n1231), .A2(new_n716), .ZN(new_n1232));
  AOI21_X1  g806(.A(new_n459), .B1(new_n665), .B2(new_n667), .ZN(new_n1233));
  NAND4_X1  g807(.A1(new_n691), .A2(new_n1232), .A3(KEYINPUT125), .A4(new_n1233), .ZN(new_n1234));
  INV_X1    g808(.A(KEYINPUT125), .ZN(new_n1235));
  NAND3_X1  g809(.A1(new_n689), .A2(new_n1233), .A3(new_n690), .ZN(new_n1236));
  OAI21_X1  g810(.A(new_n1235), .B1(G229), .B2(new_n1236), .ZN(new_n1237));
  AOI22_X1  g811(.A1(new_n934), .A2(new_n937), .B1(new_n1234), .B2(new_n1237), .ZN(new_n1238));
  INV_X1    g812(.A(KEYINPUT126), .ZN(new_n1239));
  AND3_X1   g813(.A1(new_n1020), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  AOI21_X1  g814(.A(new_n1239), .B1(new_n1020), .B2(new_n1238), .ZN(new_n1241));
  OAI21_X1  g815(.A(new_n1230), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g816(.A1(new_n1020), .A2(new_n1238), .ZN(new_n1243));
  NAND2_X1  g817(.A1(new_n1243), .A2(KEYINPUT126), .ZN(new_n1244));
  NAND3_X1  g818(.A1(new_n1020), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1245));
  NAND3_X1  g819(.A1(new_n1244), .A2(KEYINPUT127), .A3(new_n1245), .ZN(new_n1246));
  NAND2_X1  g820(.A1(new_n1242), .A2(new_n1246), .ZN(G308));
  NAND2_X1  g821(.A1(new_n1244), .A2(new_n1245), .ZN(G225));
endmodule


