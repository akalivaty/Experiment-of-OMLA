//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 0 0 0 1 0 1 0 1 0 1 0 1 0 0 0 1 0 0 0 1 1 0 0 0 1 0 1 0 1 0 0 1 0 1 1 0 0 1 1 1 1 0 0 0 0 1 0 0 0 0 0 0 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:08 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n608, new_n609, new_n610,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n616, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958;
  INV_X1    g000(.A(G125), .ZN(new_n187));
  OR3_X1    g001(.A1(new_n187), .A2(KEYINPUT16), .A3(G140), .ZN(new_n188));
  XOR2_X1   g002(.A(G125), .B(G140), .Z(new_n189));
  INV_X1    g003(.A(KEYINPUT16), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n188), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n191), .B(new_n192), .ZN(new_n193));
  XOR2_X1   g007(.A(KEYINPUT24), .B(G110), .Z(new_n194));
  INV_X1    g008(.A(G119), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G128), .ZN(new_n196));
  INV_X1    g010(.A(G128), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G119), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n194), .A2(new_n196), .A3(new_n198), .ZN(new_n199));
  XNOR2_X1  g013(.A(new_n198), .B(KEYINPUT23), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(new_n196), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G110), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n193), .A2(new_n199), .A3(new_n202), .ZN(new_n203));
  OR2_X1    g017(.A1(new_n191), .A2(new_n192), .ZN(new_n204));
  INV_X1    g018(.A(new_n189), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(new_n192), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n201), .A2(G110), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n194), .B1(new_n196), .B2(new_n198), .ZN(new_n208));
  OAI211_X1 g022(.A(new_n204), .B(new_n206), .C1(new_n207), .C2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n203), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G953), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n211), .A2(G221), .A3(G234), .ZN(new_n212));
  XNOR2_X1  g026(.A(new_n212), .B(KEYINPUT22), .ZN(new_n213));
  XNOR2_X1  g027(.A(new_n213), .B(G137), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n210), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G902), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n203), .A2(new_n209), .A3(new_n214), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  OR2_X1    g033(.A1(new_n219), .A2(KEYINPUT25), .ZN(new_n220));
  XNOR2_X1  g034(.A(KEYINPUT74), .B(G217), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n217), .A2(G234), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n219), .A2(KEYINPUT25), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n220), .A2(new_n221), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  AND2_X1   g038(.A1(new_n216), .A2(new_n218), .ZN(new_n225));
  AOI21_X1  g039(.A(G902), .B1(new_n221), .B2(new_n222), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT70), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n229), .B1(new_n195), .B2(G116), .ZN(new_n230));
  INV_X1    g044(.A(G116), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n231), .A2(KEYINPUT70), .A3(G119), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n195), .A2(G116), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(KEYINPUT2), .B(G113), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n236), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n238), .A2(new_n233), .A3(new_n234), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G131), .ZN(new_n242));
  INV_X1    g056(.A(G137), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n243), .A2(G134), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT11), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n246), .B1(G134), .B2(new_n243), .ZN(new_n247));
  INV_X1    g061(.A(G134), .ZN(new_n248));
  NOR3_X1   g062(.A1(new_n248), .A2(KEYINPUT11), .A3(G137), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n242), .B(new_n245), .C1(new_n247), .C2(new_n249), .ZN(new_n250));
  OAI21_X1  g064(.A(KEYINPUT66), .B1(new_n243), .B2(G134), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT66), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n252), .A2(new_n248), .A3(G137), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n243), .A2(G134), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n251), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  AOI22_X1  g069(.A1(new_n250), .A2(KEYINPUT67), .B1(G131), .B2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n255), .A2(KEYINPUT67), .A3(G131), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  OAI21_X1  g072(.A(KEYINPUT68), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G143), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n260), .B(G146), .C1(new_n197), .C2(KEYINPUT1), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n197), .A2(new_n192), .A3(G143), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT69), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n261), .A2(KEYINPUT69), .A3(new_n262), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n197), .A2(KEYINPUT1), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n192), .A2(G143), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n260), .A2(G146), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n265), .A2(new_n266), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT68), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT67), .ZN(new_n273));
  OAI21_X1  g087(.A(KEYINPUT11), .B1(new_n248), .B2(G137), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n246), .A2(new_n243), .A3(G134), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n244), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n273), .B1(new_n276), .B2(new_n242), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n255), .A2(G131), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n272), .B(new_n257), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n259), .A2(new_n271), .A3(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n245), .B1(new_n247), .B2(new_n249), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n281), .A2(KEYINPUT65), .A3(G131), .ZN(new_n282));
  AOI21_X1  g096(.A(KEYINPUT65), .B1(new_n276), .B2(new_n242), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n281), .A2(G131), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n268), .A2(new_n269), .ZN(new_n286));
  OR2_X1    g100(.A1(KEYINPUT0), .A2(G128), .ZN(new_n287));
  NAND2_X1  g101(.A1(KEYINPUT0), .A2(G128), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  XNOR2_X1  g103(.A(G143), .B(G146), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n290), .A2(KEYINPUT0), .A3(G128), .ZN(new_n291));
  AND2_X1   g105(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT64), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AND3_X1   g108(.A1(new_n289), .A2(new_n291), .A3(new_n293), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n282), .B(new_n285), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n241), .B1(new_n280), .B2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n285), .A2(new_n292), .A3(new_n282), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n271), .B(new_n257), .C1(new_n278), .C2(new_n277), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT71), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n240), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n237), .A2(KEYINPUT71), .A3(new_n239), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n298), .A2(new_n299), .A3(new_n301), .A4(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(KEYINPUT28), .B1(new_n297), .B2(new_n304), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n304), .A2(KEYINPUT28), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n309));
  XNOR2_X1  g123(.A(new_n309), .B(G101), .ZN(new_n310));
  INV_X1    g124(.A(G237), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT72), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT72), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G237), .ZN(new_n314));
  AOI21_X1  g128(.A(G953), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G210), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n310), .B(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n308), .A2(new_n318), .ZN(new_n319));
  AND3_X1   g133(.A1(new_n298), .A2(new_n299), .A3(KEYINPUT30), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n280), .A2(new_n296), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT30), .ZN(new_n322));
  AOI211_X1 g136(.A(new_n241), .B(new_n320), .C1(new_n321), .C2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n303), .A2(new_n317), .ZN(new_n324));
  OAI21_X1  g138(.A(KEYINPUT31), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n240), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT31), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n327), .A2(new_n328), .A3(new_n303), .A4(new_n317), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n319), .A2(new_n325), .A3(new_n329), .ZN(new_n330));
  NOR2_X1   g144(.A1(G472), .A2(G902), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT32), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT32), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n330), .A2(new_n334), .A3(new_n331), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n318), .B1(new_n305), .B2(new_n307), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n327), .A2(new_n303), .A3(new_n318), .ZN(new_n339));
  AOI21_X1  g153(.A(KEYINPUT29), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n298), .A2(new_n299), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n301), .A2(new_n302), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n303), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(KEYINPUT28), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(KEYINPUT73), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT73), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n344), .A2(new_n347), .A3(KEYINPUT28), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n346), .A2(KEYINPUT29), .A3(new_n307), .A4(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n217), .B1(new_n349), .B2(new_n318), .ZN(new_n350));
  OAI21_X1  g164(.A(G472), .B1(new_n340), .B2(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n228), .B1(new_n336), .B2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(G469), .ZN(new_n353));
  XNOR2_X1  g167(.A(G110), .B(G140), .ZN(new_n354));
  AND2_X1   g168(.A1(new_n211), .A2(G227), .ZN(new_n355));
  XOR2_X1   g169(.A(new_n354), .B(new_n355), .Z(new_n356));
  INV_X1    g170(.A(G107), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n357), .A2(G104), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT3), .ZN(new_n359));
  INV_X1    g173(.A(G104), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n360), .A2(G107), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n358), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(KEYINPUT3), .B1(new_n360), .B2(G107), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(KEYINPUT75), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT75), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n365), .B(KEYINPUT3), .C1(new_n360), .C2(G107), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n362), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G101), .ZN(new_n368));
  INV_X1    g182(.A(G101), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n362), .A2(new_n369), .A3(new_n364), .A4(new_n366), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n368), .A2(KEYINPUT4), .A3(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT4), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n367), .A2(new_n372), .A3(G101), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n371), .A2(new_n292), .A3(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(G101), .B1(new_n358), .B2(new_n361), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n370), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT77), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n376), .A2(new_n377), .A3(KEYINPUT10), .A4(new_n271), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n271), .A2(KEYINPUT10), .A3(new_n375), .A4(new_n370), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(KEYINPUT77), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT76), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n270), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n290), .A2(KEYINPUT76), .A3(new_n267), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n375), .B(new_n370), .C1(new_n384), .C2(new_n263), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT10), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n374), .A2(new_n378), .A3(new_n380), .A4(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n285), .A2(new_n282), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(KEYINPUT80), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT80), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n388), .A2(new_n393), .A3(new_n390), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n389), .B(KEYINPUT78), .ZN(new_n396));
  AND2_X1   g210(.A1(new_n378), .A2(new_n380), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n396), .A2(new_n397), .A3(new_n374), .A4(new_n387), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n356), .B1(new_n395), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT12), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT79), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n400), .B1(new_n389), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n385), .B1(new_n376), .B2(new_n271), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n390), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n402), .A2(new_n390), .A3(new_n404), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AND3_X1   g222(.A1(new_n408), .A2(new_n398), .A3(new_n356), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n353), .B(new_n217), .C1(new_n399), .C2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT78), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n389), .B(new_n411), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n388), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n356), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n408), .A2(new_n398), .ZN(new_n416));
  AOI22_X1  g230(.A1(new_n395), .A2(new_n415), .B1(new_n416), .B2(new_n414), .ZN(new_n417));
  OAI21_X1  g231(.A(G469), .B1(new_n417), .B2(G902), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n410), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(G214), .B1(G237), .B2(G902), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT81), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n422), .B1(new_n271), .B2(G125), .ZN(new_n423));
  AOI22_X1  g237(.A1(new_n263), .A2(new_n264), .B1(new_n290), .B2(new_n267), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n424), .A2(KEYINPUT81), .A3(new_n187), .A4(new_n266), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(KEYINPUT85), .ZN(new_n427));
  OR2_X1    g241(.A1(new_n292), .A2(new_n187), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT85), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n423), .A2(new_n429), .A3(new_n425), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n427), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n211), .A2(G224), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(KEYINPUT7), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n371), .A2(new_n240), .A3(new_n373), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT5), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n235), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(G113), .B1(new_n234), .B2(KEYINPUT5), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n376), .B(new_n239), .C1(new_n437), .C2(new_n438), .ZN(new_n439));
  XOR2_X1   g253(.A(G110), .B(G122), .Z(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n435), .A2(new_n439), .A3(new_n441), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n426), .A2(KEYINPUT7), .A3(new_n432), .A4(new_n428), .ZN(new_n443));
  AND2_X1   g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n438), .B(KEYINPUT83), .ZN(new_n445));
  OAI21_X1  g259(.A(KEYINPUT82), .B1(new_n235), .B2(new_n436), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT82), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n233), .A2(new_n447), .A3(KEYINPUT5), .A4(new_n234), .ZN(new_n448));
  AND3_X1   g262(.A1(new_n445), .A2(new_n446), .A3(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n239), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n376), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n239), .B1(new_n437), .B2(new_n438), .ZN(new_n452));
  OR2_X1    g266(.A1(new_n452), .A2(new_n376), .ZN(new_n453));
  XOR2_X1   g267(.A(new_n440), .B(KEYINPUT8), .Z(new_n454));
  NAND3_X1  g268(.A1(new_n451), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT84), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n451), .A2(KEYINPUT84), .A3(new_n453), .A4(new_n454), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n434), .A2(new_n444), .A3(new_n457), .A4(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n435), .A2(new_n439), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n440), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n461), .A2(KEYINPUT6), .A3(new_n442), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT6), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n460), .A2(new_n463), .A3(new_n440), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n426), .A2(new_n428), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n465), .A2(G224), .A3(new_n211), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n426), .A2(new_n432), .A3(new_n428), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n462), .A2(new_n464), .A3(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n459), .A2(new_n469), .A3(new_n217), .ZN(new_n470));
  OAI21_X1  g284(.A(G210), .B1(G237), .B2(G902), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n459), .A2(new_n469), .A3(new_n217), .A4(new_n471), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n421), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(G221), .ZN(new_n476));
  XOR2_X1   g290(.A(KEYINPUT9), .B(G234), .Z(new_n477));
  AOI21_X1  g291(.A(new_n476), .B1(new_n477), .B2(new_n217), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  AND3_X1   g293(.A1(new_n419), .A2(new_n475), .A3(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(G128), .B(G143), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(KEYINPUT13), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n260), .A2(G128), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n482), .B(G134), .C1(KEYINPUT13), .C2(new_n483), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n484), .B(KEYINPUT88), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n481), .A2(new_n248), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT87), .ZN(new_n487));
  INV_X1    g301(.A(G122), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n487), .B1(new_n488), .B2(G116), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n231), .A2(KEYINPUT87), .A3(G122), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n491), .B1(new_n231), .B2(G122), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n492), .B(G107), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n485), .A2(new_n486), .A3(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n481), .B(new_n248), .ZN(new_n495));
  OR2_X1    g309(.A1(new_n492), .A2(G107), .ZN(new_n496));
  AND3_X1   g310(.A1(new_n491), .A2(KEYINPUT89), .A3(KEYINPUT14), .ZN(new_n497));
  OAI22_X1  g311(.A1(new_n491), .A2(KEYINPUT14), .B1(new_n231), .B2(G122), .ZN(new_n498));
  AOI21_X1  g312(.A(KEYINPUT89), .B1(new_n491), .B2(KEYINPUT14), .ZN(new_n499));
  NOR3_X1   g313(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n495), .B(new_n496), .C1(new_n500), .C2(new_n357), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n494), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n477), .A2(new_n211), .A3(new_n221), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n503), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n494), .A2(new_n505), .A3(new_n501), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n217), .ZN(new_n508));
  INV_X1    g322(.A(G478), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n509), .A2(KEYINPUT15), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n508), .B(new_n511), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n315), .A2(G143), .A3(G214), .ZN(new_n513));
  AOI21_X1  g327(.A(G143), .B1(new_n315), .B2(G214), .ZN(new_n514));
  OAI21_X1  g328(.A(G131), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n315), .A2(G214), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n260), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n315), .A2(G143), .A3(G214), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n517), .A2(new_n242), .A3(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT17), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n515), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n191), .B(G146), .ZN(new_n522));
  OAI211_X1 g336(.A(KEYINPUT17), .B(G131), .C1(new_n513), .C2(new_n514), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  XNOR2_X1  g338(.A(G113), .B(G122), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n525), .B(new_n360), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT18), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n517), .B(new_n518), .C1(new_n527), .C2(new_n242), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n189), .A2(G146), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n206), .A2(new_n529), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n528), .B(new_n530), .C1(new_n527), .C2(new_n515), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n524), .A2(new_n526), .A3(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT86), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n524), .A2(KEYINPUT86), .A3(new_n526), .A4(new_n531), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n515), .A2(new_n519), .ZN(new_n537));
  XOR2_X1   g351(.A(new_n189), .B(KEYINPUT19), .Z(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(new_n192), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n537), .A2(new_n204), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(new_n531), .ZN(new_n541));
  INV_X1    g355(.A(new_n526), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n536), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(G475), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n544), .A2(new_n545), .A3(new_n217), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT20), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n524), .A2(new_n531), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n542), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n536), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n217), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(G475), .ZN(new_n553));
  AOI21_X1  g367(.A(G475), .B1(new_n536), .B2(new_n543), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n554), .A2(KEYINPUT20), .A3(new_n217), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n512), .A2(new_n548), .A3(new_n553), .A4(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(G234), .A2(G237), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n557), .A2(G952), .A3(new_n211), .ZN(new_n558));
  XOR2_X1   g372(.A(new_n558), .B(KEYINPUT90), .Z(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  XOR2_X1   g374(.A(KEYINPUT21), .B(G898), .Z(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n557), .A2(G902), .A3(G953), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n560), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n556), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n352), .A2(new_n480), .A3(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n567), .B(G101), .ZN(G3));
  NAND3_X1  g382(.A1(new_n548), .A2(new_n553), .A3(new_n555), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n506), .A2(KEYINPUT92), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT92), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n494), .A2(new_n571), .A3(new_n505), .A4(new_n501), .ZN(new_n572));
  XOR2_X1   g386(.A(new_n503), .B(KEYINPUT91), .Z(new_n573));
  NAND2_X1  g387(.A1(new_n502), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n570), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(KEYINPUT33), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT33), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n504), .A2(new_n577), .A3(new_n506), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n579), .A2(G478), .A3(new_n217), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n508), .A2(new_n509), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n565), .ZN(new_n583));
  AND4_X1   g397(.A1(new_n475), .A2(new_n569), .A3(new_n582), .A4(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n330), .A2(new_n217), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(G472), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n332), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  AOI211_X1 g402(.A(new_n478), .B(new_n228), .C1(new_n410), .C2(new_n418), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n584), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  XOR2_X1   g404(.A(KEYINPUT34), .B(G104), .Z(new_n591));
  XNOR2_X1  g405(.A(new_n590), .B(new_n591), .ZN(G6));
  NAND2_X1  g406(.A1(new_n473), .A2(new_n474), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n593), .A2(new_n420), .A3(new_n583), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n508), .B(new_n510), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n595), .A2(new_n548), .A3(new_n553), .A4(new_n555), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n589), .A2(new_n588), .A3(new_n597), .ZN(new_n598));
  XOR2_X1   g412(.A(KEYINPUT35), .B(G107), .Z(new_n599));
  XNOR2_X1  g413(.A(new_n598), .B(new_n599), .ZN(G9));
  NOR2_X1   g414(.A1(new_n215), .A2(KEYINPUT36), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n210), .B(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n226), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n224), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n480), .A2(new_n588), .A3(new_n566), .A4(new_n604), .ZN(new_n605));
  XOR2_X1   g419(.A(new_n605), .B(KEYINPUT37), .Z(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(G110), .ZN(G12));
  INV_X1    g421(.A(new_n335), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n334), .B1(new_n330), .B2(new_n331), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n351), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n610), .A2(new_n604), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n611), .A2(new_n480), .ZN(new_n612));
  INV_X1    g426(.A(G900), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n560), .B1(new_n613), .B2(new_n564), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n596), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(G128), .ZN(G30));
  AOI21_X1  g431(.A(new_n478), .B1(new_n410), .B2(new_n418), .ZN(new_n618));
  XOR2_X1   g432(.A(new_n614), .B(KEYINPUT39), .Z(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  XOR2_X1   g434(.A(new_n620), .B(KEYINPUT40), .Z(new_n621));
  XNOR2_X1  g435(.A(new_n593), .B(KEYINPUT38), .ZN(new_n622));
  AOI21_X1  g436(.A(KEYINPUT20), .B1(new_n554), .B2(new_n217), .ZN(new_n623));
  AOI22_X1  g437(.A1(new_n534), .A2(new_n535), .B1(new_n542), .B2(new_n541), .ZN(new_n624));
  NOR4_X1   g438(.A1(new_n624), .A2(new_n547), .A3(G475), .A4(G902), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n545), .B1(new_n551), .B2(new_n217), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n623), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NOR3_X1   g441(.A1(new_n627), .A2(new_n421), .A3(new_n512), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n318), .B1(new_n327), .B2(new_n303), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n217), .B1(new_n344), .B2(new_n317), .ZN(new_n630));
  OAI21_X1  g444(.A(G472), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(KEYINPUT93), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n336), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n633), .A2(new_n604), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n621), .A2(new_n622), .A3(new_n628), .A4(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G143), .ZN(G45));
  AND2_X1   g450(.A1(new_n569), .A2(new_n582), .ZN(new_n637));
  INV_X1    g451(.A(new_n614), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n612), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(G146), .ZN(G48));
  INV_X1    g456(.A(new_n394), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n393), .B1(new_n388), .B2(new_n390), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n398), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n409), .B1(new_n645), .B2(new_n414), .ZN(new_n646));
  OAI21_X1  g460(.A(G469), .B1(new_n646), .B2(G902), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n647), .A2(new_n479), .A3(new_n410), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(KEYINPUT94), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT94), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n647), .A2(new_n650), .A3(new_n479), .A4(new_n410), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n652), .A2(new_n352), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n584), .ZN(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT41), .B(G113), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G15));
  NAND2_X1  g470(.A1(new_n653), .A2(new_n597), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G116), .ZN(G18));
  INV_X1    g472(.A(new_n648), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n659), .A2(KEYINPUT95), .A3(new_n475), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT95), .ZN(new_n661));
  INV_X1    g475(.A(new_n475), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n661), .B1(new_n648), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n664), .A2(new_n566), .A3(new_n611), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G119), .ZN(G21));
  AOI21_X1  g480(.A(new_n347), .B1(new_n344), .B2(KEYINPUT28), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT28), .ZN(new_n668));
  AOI211_X1 g482(.A(KEYINPUT73), .B(new_n668), .C1(new_n343), .C2(new_n303), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n667), .A2(new_n669), .A3(new_n306), .ZN(new_n670));
  OAI211_X1 g484(.A(KEYINPUT96), .B(new_n325), .C1(new_n670), .C2(new_n317), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n329), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n346), .A2(new_n307), .A3(new_n348), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n318), .ZN(new_n674));
  AOI21_X1  g488(.A(KEYINPUT96), .B1(new_n674), .B2(new_n325), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n331), .B1(new_n672), .B2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT97), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n324), .B1(new_n326), .B2(new_n240), .ZN(new_n678));
  AOI22_X1  g492(.A1(new_n318), .A2(new_n308), .B1(new_n678), .B2(new_n328), .ZN(new_n679));
  AOI21_X1  g493(.A(G902), .B1(new_n679), .B2(new_n325), .ZN(new_n680));
  INV_X1    g494(.A(G472), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n677), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n585), .A2(KEYINPUT97), .A3(G472), .ZN(new_n683));
  AND3_X1   g497(.A1(new_n676), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n228), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n569), .A2(new_n420), .A3(new_n593), .A4(new_n595), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n686), .A2(new_n565), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n684), .A2(new_n652), .A3(new_n685), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(KEYINPUT98), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(new_n488), .ZN(G24));
  NAND4_X1  g504(.A1(new_n676), .A2(new_n604), .A3(new_n682), .A4(new_n683), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(KEYINPUT99), .ZN(new_n692));
  AOI21_X1  g506(.A(KEYINPUT97), .B1(new_n585), .B2(G472), .ZN(new_n693));
  AOI211_X1 g507(.A(new_n677), .B(new_n681), .C1(new_n330), .C2(new_n217), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT99), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n695), .A2(new_n696), .A3(new_n604), .A4(new_n676), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n692), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n639), .B1(new_n660), .B2(new_n663), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(KEYINPUT100), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT100), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n698), .A2(new_n699), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G125), .ZN(G27));
  INV_X1    g519(.A(KEYINPUT101), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT29), .ZN(new_n707));
  AOI211_X1 g521(.A(new_n304), .B(new_n317), .C1(new_n326), .C2(new_n240), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n707), .B1(new_n708), .B2(new_n337), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n670), .A2(KEYINPUT29), .A3(new_n317), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n709), .A2(new_n710), .A3(new_n217), .ZN(new_n711));
  AOI22_X1  g525(.A1(new_n333), .A2(new_n335), .B1(G472), .B2(new_n711), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n706), .B1(new_n712), .B2(new_n228), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n473), .A2(new_n420), .A3(new_n474), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n715), .A2(new_n569), .A3(new_n582), .A4(new_n638), .ZN(new_n716));
  INV_X1    g530(.A(new_n618), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n610), .A2(KEYINPUT101), .A3(new_n685), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n713), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n716), .A2(new_n717), .A3(KEYINPUT42), .ZN(new_n721));
  AOI22_X1  g535(.A1(new_n720), .A2(KEYINPUT42), .B1(new_n352), .B2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G131), .ZN(G33));
  OAI21_X1  g537(.A(KEYINPUT102), .B1(new_n596), .B2(new_n614), .ZN(new_n724));
  AND3_X1   g538(.A1(new_n724), .A2(new_n618), .A3(new_n715), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT102), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n627), .A2(new_n726), .A3(new_n595), .A4(new_n638), .ZN(new_n727));
  AND3_X1   g541(.A1(new_n727), .A2(new_n610), .A3(new_n685), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT103), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n725), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n724), .A2(new_n618), .A3(new_n715), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n727), .A2(new_n610), .A3(new_n685), .ZN(new_n732));
  OAI21_X1  g546(.A(KEYINPUT103), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G134), .ZN(G36));
  AOI21_X1  g549(.A(new_n569), .B1(new_n581), .B2(new_n580), .ZN(new_n736));
  NAND2_X1  g550(.A1(KEYINPUT106), .A2(KEYINPUT43), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g553(.A1(KEYINPUT106), .A2(KEYINPUT43), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n739), .B1(new_n736), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n587), .A2(new_n604), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(KEYINPUT107), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n746), .A2(KEYINPUT44), .ZN(new_n747));
  OR2_X1    g561(.A1(new_n747), .A2(KEYINPUT108), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n714), .B1(new_n746), .B2(KEYINPUT44), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n747), .A2(KEYINPUT108), .ZN(new_n750));
  AND3_X1   g564(.A1(new_n748), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  XOR2_X1   g565(.A(new_n417), .B(KEYINPUT45), .Z(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(G469), .ZN(new_n753));
  NAND2_X1  g567(.A1(G469), .A2(G902), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT46), .ZN(new_n756));
  OR3_X1    g570(.A1(new_n755), .A2(KEYINPUT104), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n755), .A2(new_n756), .ZN(new_n758));
  OAI21_X1  g572(.A(KEYINPUT104), .B1(new_n755), .B2(new_n756), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n757), .A2(new_n410), .A3(new_n758), .A4(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n760), .A2(new_n479), .A3(new_n619), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(KEYINPUT105), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n751), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G137), .ZN(G39));
  NAND2_X1  g578(.A1(new_n760), .A2(new_n479), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT47), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n760), .A2(KEYINPUT47), .A3(new_n479), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n716), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n769), .A2(new_n712), .A3(new_n228), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G140), .ZN(G42));
  NOR4_X1   g585(.A1(new_n743), .A2(new_n559), .A3(new_n648), .A4(new_n714), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n698), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n633), .A2(new_n560), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  NOR3_X1   g589(.A1(new_n648), .A2(new_n228), .A3(new_n714), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  OR3_X1    g591(.A1(new_n777), .A2(new_n569), .A3(new_n582), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n773), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n743), .A2(new_n559), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n684), .A2(new_n685), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n622), .A2(new_n420), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n780), .A2(new_n659), .A3(new_n781), .A4(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT115), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n783), .A2(new_n784), .A3(KEYINPUT50), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n784), .A2(KEYINPUT50), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n784), .A2(KEYINPUT50), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n783), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT116), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  OAI21_X1  g605(.A(KEYINPUT116), .B1(new_n785), .B2(new_n788), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n779), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT117), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n647), .A2(new_n410), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n767), .B(new_n768), .C1(new_n479), .C2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n780), .A2(new_n781), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n797), .A2(new_n715), .A3(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(KEYINPUT51), .B1(new_n795), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n799), .A2(new_n664), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n772), .A2(new_n713), .A3(new_n719), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(KEYINPUT48), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n804), .A2(G952), .A3(new_n211), .ZN(new_n805));
  INV_X1    g619(.A(new_n779), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(KEYINPUT118), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n800), .A2(new_n807), .A3(new_n789), .ZN(new_n808));
  OAI21_X1  g622(.A(KEYINPUT51), .B1(new_n806), .B2(KEYINPUT118), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n802), .B(new_n805), .C1(new_n808), .C2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n775), .A2(new_n637), .A3(new_n776), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT114), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n612), .B1(new_n615), .B2(new_n640), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n717), .A2(new_n686), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n634), .A2(new_n638), .A3(new_n815), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n698), .A2(new_n699), .A3(new_n702), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n702), .B1(new_n698), .B2(new_n699), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n814), .B(new_n816), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(KEYINPUT52), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT52), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n704), .A2(new_n821), .A3(new_n814), .A4(new_n816), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n652), .B(new_n352), .C1(new_n584), .C2(new_n597), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n688), .A2(new_n823), .ZN(new_n824));
  AOI211_X1 g638(.A(new_n421), .B(new_n565), .C1(new_n473), .C2(new_n474), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n825), .A2(KEYINPUT111), .A3(new_n595), .A4(new_n627), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT111), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n827), .B1(new_n594), .B2(new_n596), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n826), .A2(new_n828), .A3(new_n588), .A4(new_n589), .ZN(new_n829));
  AND4_X1   g643(.A1(new_n567), .A2(new_n829), .A3(new_n590), .A4(new_n605), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT112), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n831), .B1(new_n556), .B2(new_n614), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n627), .A2(KEYINPUT112), .A3(new_n512), .A4(new_n638), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n832), .A2(new_n833), .A3(new_n715), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT113), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n832), .A2(new_n833), .A3(KEYINPUT113), .A4(new_n715), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n836), .A2(new_n618), .A3(new_n611), .A4(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n824), .A2(new_n830), .A3(new_n665), .A4(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n698), .A2(new_n718), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n722), .A2(new_n734), .A3(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n820), .A2(new_n822), .A3(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n820), .A2(new_n822), .A3(new_n842), .A4(KEYINPUT53), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n845), .A2(KEYINPUT54), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(KEYINPUT54), .B1(new_n845), .B2(new_n846), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n813), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n845), .A2(new_n846), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT54), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n845), .A2(KEYINPUT54), .A3(new_n846), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n852), .A2(KEYINPUT114), .A3(new_n853), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n811), .A2(new_n812), .A3(new_n849), .A4(new_n854), .ZN(new_n855));
  OAI22_X1  g669(.A1(new_n801), .A2(new_n855), .B1(G952), .B2(G953), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n228), .A2(new_n421), .A3(new_n478), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n857), .B(KEYINPUT109), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n796), .A2(KEYINPUT49), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n858), .A2(new_n736), .A3(new_n859), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n860), .B(KEYINPUT110), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n796), .A2(KEYINPUT49), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n622), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n861), .A2(new_n633), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n856), .A2(new_n864), .ZN(G75));
  AOI21_X1  g679(.A(new_n217), .B1(new_n845), .B2(new_n846), .ZN(new_n866));
  AOI21_X1  g680(.A(KEYINPUT56), .B1(new_n866), .B2(G210), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT120), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n462), .A2(new_n464), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n869), .B(new_n468), .ZN(new_n870));
  XNOR2_X1  g684(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n870), .B(new_n871), .Z(new_n872));
  AND3_X1   g686(.A1(new_n867), .A2(new_n868), .A3(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n211), .A2(G952), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n875), .B1(new_n867), .B2(new_n868), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n872), .B1(new_n867), .B2(new_n868), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n873), .A2(new_n876), .A3(new_n877), .ZN(G51));
  XOR2_X1   g692(.A(new_n646), .B(KEYINPUT121), .Z(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n847), .A2(new_n848), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n754), .B(KEYINPUT57), .Z(new_n882));
  AOI21_X1  g696(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  AOI211_X1 g697(.A(new_n217), .B(new_n753), .C1(new_n845), .C2(new_n846), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n875), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(KEYINPUT122), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT122), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n887), .B(new_n875), .C1(new_n883), .C2(new_n884), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n886), .A2(new_n888), .ZN(G54));
  NAND3_X1  g703(.A1(new_n866), .A2(KEYINPUT58), .A3(G475), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(new_n624), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n891), .A2(new_n874), .ZN(G60));
  NAND2_X1  g706(.A1(G478), .A2(G902), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT59), .Z(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n847), .A2(new_n848), .A3(new_n813), .ZN(new_n896));
  AOI21_X1  g710(.A(KEYINPUT114), .B1(new_n852), .B2(new_n853), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(new_n579), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n898), .A2(KEYINPUT123), .A3(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT123), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n894), .B1(new_n849), .B2(new_n854), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n901), .B1(new_n902), .B2(new_n579), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n899), .A2(new_n894), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n874), .B1(new_n881), .B2(new_n904), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n900), .A2(new_n903), .A3(new_n905), .ZN(G63));
  NAND2_X1  g720(.A1(G217), .A2(G902), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n907), .B(KEYINPUT60), .Z(new_n908));
  NAND2_X1  g722(.A1(new_n850), .A2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(new_n225), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n850), .A2(new_n602), .A3(new_n908), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n911), .A2(KEYINPUT61), .A3(new_n875), .A4(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT124), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n850), .A2(KEYINPUT124), .A3(new_n602), .A4(new_n908), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n915), .A2(new_n911), .A3(new_n875), .A4(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT61), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n917), .A2(KEYINPUT125), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT125), .B1(new_n917), .B2(new_n918), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n913), .B1(new_n919), .B2(new_n920), .ZN(G66));
  INV_X1    g735(.A(G224), .ZN(new_n922));
  OAI21_X1  g736(.A(G953), .B1(new_n562), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n824), .A2(new_n830), .A3(new_n665), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT126), .Z(new_n925));
  OAI21_X1  g739(.A(new_n923), .B1(new_n925), .B2(G953), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n869), .B1(G898), .B2(new_n211), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n926), .B(new_n927), .ZN(G69));
  XNOR2_X1  g742(.A(new_n326), .B(new_n538), .ZN(new_n929));
  NAND2_X1  g743(.A1(G900), .A2(G953), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n722), .A2(new_n734), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n770), .A2(new_n931), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n704), .A2(new_n814), .ZN(new_n933));
  AND4_X1   g747(.A1(new_n593), .A2(new_n713), .A3(new_n628), .A4(new_n719), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n762), .B1(new_n751), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n932), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  OAI211_X1 g750(.A(new_n929), .B(new_n930), .C1(new_n936), .C2(G953), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n933), .A2(new_n635), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT62), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n938), .B(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n569), .A2(new_n512), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n352), .B1(new_n637), .B2(new_n941), .ZN(new_n942));
  NOR3_X1   g756(.A1(new_n942), .A2(new_n620), .A3(new_n714), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n943), .B1(new_n751), .B2(new_n762), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n940), .A2(new_n770), .A3(new_n944), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n945), .A2(new_n211), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n937), .B1(new_n946), .B2(new_n929), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n211), .B1(G227), .B2(G900), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n947), .B(new_n948), .ZN(G72));
  XNOR2_X1  g763(.A(new_n708), .B(KEYINPUT127), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n932), .A2(new_n935), .A3(new_n925), .A4(new_n933), .ZN(new_n951));
  NAND2_X1  g765(.A1(G472), .A2(G902), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT63), .Z(new_n953));
  AOI21_X1  g767(.A(new_n950), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n629), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n940), .A2(new_n944), .A3(new_n770), .A4(new_n925), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n955), .B1(new_n956), .B2(new_n953), .ZN(new_n957));
  AND4_X1   g771(.A1(new_n339), .A2(new_n850), .A3(new_n955), .A4(new_n953), .ZN(new_n958));
  NOR4_X1   g772(.A1(new_n954), .A2(new_n957), .A3(new_n874), .A4(new_n958), .ZN(G57));
endmodule


