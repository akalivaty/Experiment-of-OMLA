

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753;

  BUF_X1 U366 ( .A(n700), .Z(n346) );
  XNOR2_X1 U367 ( .A(n453), .B(n452), .ZN(n366) );
  XNOR2_X1 U368 ( .A(n554), .B(n553), .ZN(n700) );
  NOR2_X1 U369 ( .A1(n675), .A2(n674), .ZN(n554) );
  XNOR2_X1 U370 ( .A(n575), .B(n345), .ZN(n671) );
  XNOR2_X1 U371 ( .A(KEYINPUT38), .B(KEYINPUT75), .ZN(n345) );
  XNOR2_X1 U372 ( .A(n687), .B(n467), .ZN(n608) );
  XNOR2_X1 U373 ( .A(n579), .B(n578), .ZN(n617) );
  OR2_X1 U374 ( .A1(n646), .A2(G902), .ZN(n440) );
  NAND2_X1 U375 ( .A1(n429), .A2(n428), .ZN(n542) );
  XNOR2_X1 U376 ( .A(n403), .B(n401), .ZN(n732) );
  XNOR2_X1 U377 ( .A(n522), .B(n521), .ZN(n403) );
  XNOR2_X1 U378 ( .A(G107), .B(KEYINPUT77), .ZN(n404) );
  NOR2_X2 U379 ( .A1(n684), .A2(n605), .ZN(n606) );
  AND2_X2 U380 ( .A1(n400), .A2(n611), .ZN(n581) );
  OR2_X2 U381 ( .A1(n710), .A2(n421), .ZN(n420) );
  XNOR2_X2 U382 ( .A(n506), .B(n471), .ZN(n717) );
  INV_X2 U383 ( .A(KEYINPUT3), .ZN(n406) );
  INV_X2 U384 ( .A(G953), .ZN(n741) );
  BUF_X1 U385 ( .A(G128), .Z(n392) );
  OR2_X1 U386 ( .A1(n569), .A2(n660), .ZN(n435) );
  NOR2_X1 U387 ( .A1(n661), .A2(n676), .ZN(n568) );
  INV_X1 U388 ( .A(n570), .ZN(n687) );
  INV_X1 U389 ( .A(KEYINPUT16), .ZN(n402) );
  INV_X1 U390 ( .A(KEYINPUT4), .ZN(n465) );
  NOR2_X1 U391 ( .A1(n641), .A2(n347), .ZN(n469) );
  AND2_X1 U392 ( .A1(n350), .A2(n665), .ZN(n445) );
  NOR2_X1 U393 ( .A1(n623), .A2(n608), .ZN(n407) );
  XNOR2_X1 U394 ( .A(n560), .B(n365), .ZN(n753) );
  NOR2_X1 U395 ( .A1(n690), .A2(n605), .ZN(n394) );
  OR2_X1 U396 ( .A1(n579), .A2(n559), .ZN(n565) );
  XNOR2_X1 U397 ( .A(n551), .B(KEYINPUT106), .ZN(n611) );
  NAND2_X1 U398 ( .A1(n416), .A2(n424), .ZN(n584) );
  XNOR2_X1 U399 ( .A(n530), .B(n402), .ZN(n401) );
  XNOR2_X1 U400 ( .A(n465), .B(G146), .ZN(n513) );
  INV_X1 U401 ( .A(KEYINPUT31), .ZN(n393) );
  XNOR2_X2 U402 ( .A(n437), .B(KEYINPUT39), .ZN(n587) );
  XNOR2_X1 U403 ( .A(n590), .B(n589), .ZN(n601) );
  XNOR2_X1 U404 ( .A(n463), .B(n462), .ZN(n738) );
  INV_X1 U405 ( .A(G140), .ZN(n462) );
  XNOR2_X1 U406 ( .A(KEYINPUT10), .B(G125), .ZN(n463) );
  NOR2_X1 U407 ( .A1(G237), .A2(G953), .ZN(n507) );
  NAND2_X1 U408 ( .A1(n422), .A2(n636), .ZN(n421) );
  INV_X1 U409 ( .A(n526), .ZN(n422) );
  XNOR2_X1 U410 ( .A(n459), .B(n457), .ZN(n562) );
  XNOR2_X1 U411 ( .A(n550), .B(n458), .ZN(n457) );
  NOR2_X1 U412 ( .A1(n724), .A2(G902), .ZN(n459) );
  INV_X1 U413 ( .A(G478), .ZN(n458) );
  OR2_X2 U414 ( .A1(n384), .A2(n381), .ZN(n579) );
  NAND2_X1 U415 ( .A1(n386), .A2(n385), .ZN(n384) );
  NAND2_X1 U416 ( .A1(n387), .A2(G902), .ZN(n385) );
  NAND2_X1 U417 ( .A1(n436), .A2(n669), .ZN(n740) );
  XNOR2_X1 U418 ( .A(n738), .B(G146), .ZN(n535) );
  NAND2_X1 U419 ( .A1(n430), .A2(n481), .ZN(n429) );
  AND2_X1 U420 ( .A1(n608), .A2(n574), .ZN(n400) );
  NOR2_X1 U421 ( .A1(n666), .A2(n613), .ZN(n614) );
  XNOR2_X1 U422 ( .A(n513), .B(n427), .ZN(n426) );
  XNOR2_X1 U423 ( .A(n482), .B(G137), .ZN(n427) );
  INV_X1 U424 ( .A(G131), .ZN(n482) );
  INV_X1 U425 ( .A(n584), .ZN(n575) );
  NAND2_X1 U426 ( .A1(n380), .A2(n379), .ZN(n374) );
  NOR2_X1 U427 ( .A1(n605), .A2(KEYINPUT34), .ZN(n379) );
  AND2_X1 U428 ( .A1(n376), .A2(n377), .ZN(n375) );
  AND2_X1 U429 ( .A1(n378), .A2(n597), .ZN(n377) );
  INV_X1 U430 ( .A(n556), .ZN(n439) );
  NAND2_X1 U431 ( .A1(n420), .A2(n418), .ZN(n417) );
  NOR2_X1 U432 ( .A1(n572), .A2(n419), .ZN(n418) );
  NOR2_X1 U433 ( .A1(n410), .A2(n425), .ZN(n409) );
  XNOR2_X1 U434 ( .A(n577), .B(n576), .ZN(n578) );
  NOR2_X2 U435 ( .A1(n579), .A2(n681), .ZN(n604) );
  XOR2_X1 U436 ( .A(KEYINPUT72), .B(KEYINPUT8), .Z(n492) );
  XOR2_X1 U437 ( .A(KEYINPUT85), .B(KEYINPUT24), .Z(n487) );
  XNOR2_X1 U438 ( .A(n392), .B(G110), .ZN(n486) );
  XNOR2_X1 U439 ( .A(n363), .B(n490), .ZN(n494) );
  XNOR2_X1 U440 ( .A(n489), .B(n364), .ZN(n363) );
  INV_X1 U441 ( .A(KEYINPUT94), .ZN(n364) );
  XOR2_X1 U442 ( .A(KEYINPUT9), .B(G107), .Z(n545) );
  XNOR2_X1 U443 ( .A(G116), .B(G122), .ZN(n544) );
  XNOR2_X1 U444 ( .A(KEYINPUT101), .B(KEYINPUT103), .ZN(n539) );
  XOR2_X1 U445 ( .A(KEYINPUT7), .B(KEYINPUT102), .Z(n540) );
  XNOR2_X1 U446 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U447 ( .A(n367), .B(n532), .ZN(n537) );
  INV_X1 U448 ( .A(KEYINPUT66), .ZN(n450) );
  INV_X1 U449 ( .A(G125), .ZN(n360) );
  NOR2_X1 U450 ( .A1(n567), .A2(n566), .ZN(n551) );
  XNOR2_X1 U451 ( .A(n501), .B(n500), .ZN(n626) );
  XNOR2_X1 U452 ( .A(n361), .B(KEYINPUT22), .ZN(n623) );
  BUF_X1 U453 ( .A(n687), .Z(n362) );
  INV_X1 U454 ( .A(n682), .ZN(n454) );
  NAND2_X1 U455 ( .A1(n348), .A2(n461), .ZN(n444) );
  XNOR2_X1 U456 ( .A(KEYINPUT96), .B(KEYINPUT12), .ZN(n370) );
  OR2_X1 U457 ( .A1(G237), .A2(G902), .ZN(n525) );
  NAND2_X1 U458 ( .A1(G469), .A2(n383), .ZN(n382) );
  INV_X1 U459 ( .A(G902), .ZN(n383) );
  NAND2_X1 U460 ( .A1(n626), .A2(n464), .ZN(n681) );
  XNOR2_X1 U461 ( .A(n369), .B(n368), .ZN(n367) );
  XNOR2_X1 U462 ( .A(n531), .B(KEYINPUT11), .ZN(n368) );
  XNOR2_X1 U463 ( .A(n530), .B(n370), .ZN(n369) );
  XNOR2_X1 U464 ( .A(G113), .B(G143), .ZN(n531) );
  XNOR2_X1 U465 ( .A(G131), .B(KEYINPUT98), .ZN(n528) );
  XOR2_X1 U466 ( .A(KEYINPUT97), .B(KEYINPUT99), .Z(n529) );
  XNOR2_X1 U467 ( .A(n371), .B(G104), .ZN(n530) );
  INV_X1 U468 ( .A(G122), .ZN(n371) );
  NAND2_X1 U469 ( .A1(G234), .A2(G237), .ZN(n475) );
  NAND2_X1 U470 ( .A1(n601), .A2(n608), .ZN(n466) );
  NAND2_X1 U471 ( .A1(n526), .A2(n524), .ZN(n423) );
  XNOR2_X1 U472 ( .A(n506), .B(n441), .ZN(n646) );
  XNOR2_X1 U473 ( .A(n508), .B(KEYINPUT5), .ZN(n509) );
  XOR2_X1 U474 ( .A(G104), .B(G140), .Z(n484) );
  BUF_X1 U475 ( .A(n699), .Z(n396) );
  NAND2_X1 U476 ( .A1(n448), .A2(n357), .ZN(n447) );
  XNOR2_X1 U477 ( .A(n600), .B(n599), .ZN(n628) );
  NAND2_X1 U478 ( .A1(n375), .A2(n374), .ZN(n600) );
  AND2_X1 U479 ( .A1(n420), .A2(n423), .ZN(n416) );
  AND2_X1 U480 ( .A1(n512), .A2(n438), .ZN(n563) );
  NOR2_X1 U481 ( .A1(n572), .A2(n570), .ZN(n511) );
  XNOR2_X1 U482 ( .A(n373), .B(n372), .ZN(n566) );
  XNOR2_X1 U483 ( .A(n538), .B(G475), .ZN(n372) );
  OR2_X1 U484 ( .A1(n720), .A2(G902), .ZN(n373) );
  NAND2_X1 U485 ( .A1(n411), .A2(n409), .ZN(n408) );
  AND2_X1 U486 ( .A1(n413), .A2(n415), .ZN(n412) );
  INV_X1 U487 ( .A(n417), .ZN(n411) );
  XNOR2_X1 U488 ( .A(n495), .B(n496), .ZN(n643) );
  XNOR2_X1 U489 ( .A(n549), .B(n548), .ZN(n724) );
  XNOR2_X1 U490 ( .A(n547), .B(n546), .ZN(n548) );
  NAND2_X1 U491 ( .A1(n524), .A2(KEYINPUT2), .ZN(n470) );
  XNOR2_X1 U492 ( .A(n732), .B(n523), .ZN(n710) );
  XNOR2_X1 U493 ( .A(n520), .B(n359), .ZN(n523) );
  XNOR2_X1 U494 ( .A(n519), .B(n360), .ZN(n359) );
  INV_X1 U495 ( .A(KEYINPUT42), .ZN(n365) );
  XNOR2_X1 U496 ( .A(n358), .B(n552), .ZN(n752) );
  INV_X1 U497 ( .A(KEYINPUT114), .ZN(n452) );
  NAND2_X1 U498 ( .A1(n455), .A2(n454), .ZN(n453) );
  XNOR2_X1 U499 ( .A(n456), .B(n352), .ZN(n455) );
  BUF_X1 U500 ( .A(n628), .Z(n750) );
  NOR2_X1 U501 ( .A1(n626), .A2(n625), .ZN(n655) );
  NOR2_X1 U502 ( .A1(n705), .A2(G953), .ZN(n460) );
  NAND2_X1 U503 ( .A1(n669), .A2(n524), .ZN(n347) );
  XOR2_X1 U504 ( .A(G902), .B(KEYINPUT15), .Z(n524) );
  XOR2_X1 U505 ( .A(n447), .B(KEYINPUT83), .Z(n348) );
  AND2_X1 U506 ( .A1(n391), .A2(n390), .ZN(n349) );
  AND2_X1 U507 ( .A1(n446), .A2(n653), .ZN(n350) );
  XOR2_X1 U508 ( .A(n510), .B(KEYINPUT73), .Z(n351) );
  INV_X1 U509 ( .A(G469), .ZN(n387) );
  INV_X1 U510 ( .A(KEYINPUT19), .ZN(n425) );
  XNOR2_X1 U511 ( .A(KEYINPUT113), .B(KEYINPUT36), .ZN(n352) );
  XOR2_X1 U512 ( .A(KEYINPUT108), .B(KEYINPUT33), .Z(n353) );
  XOR2_X1 U513 ( .A(n720), .B(n719), .Z(n354) );
  XOR2_X1 U514 ( .A(n646), .B(n645), .Z(n355) );
  XOR2_X1 U515 ( .A(n643), .B(KEYINPUT124), .Z(n356) );
  XOR2_X1 U516 ( .A(KEYINPUT84), .B(KEYINPUT2), .Z(n357) );
  NOR2_X1 U517 ( .A1(G952), .A2(n741), .ZN(n726) );
  INV_X1 U518 ( .A(n726), .ZN(n390) );
  NAND2_X1 U519 ( .A1(n617), .A2(n588), .ZN(n590) );
  NAND2_X1 U520 ( .A1(n587), .A2(n611), .ZN(n358) );
  AND2_X1 U521 ( .A1(n474), .A2(n439), .ZN(n438) );
  NAND2_X1 U522 ( .A1(n612), .A2(n611), .ZN(n665) );
  XNOR2_X1 U523 ( .A(n394), .B(n393), .ZN(n612) );
  NAND2_X1 U524 ( .A1(n601), .A2(n362), .ZN(n690) );
  NAND2_X1 U525 ( .A1(n606), .A2(n607), .ZN(n361) );
  NOR2_X1 U526 ( .A1(n580), .A2(n435), .ZN(n434) );
  XNOR2_X2 U527 ( .A(n405), .B(n505), .ZN(n522) );
  NAND2_X1 U528 ( .A1(n752), .A2(n753), .ZN(n395) );
  XNOR2_X1 U529 ( .A(n366), .B(n751), .ZN(G27) );
  XNOR2_X1 U530 ( .A(n366), .B(KEYINPUT88), .ZN(n580) );
  NAND2_X1 U531 ( .A1(n699), .A2(KEYINPUT34), .ZN(n376) );
  NAND2_X1 U532 ( .A1(n605), .A2(KEYINPUT34), .ZN(n378) );
  INV_X1 U533 ( .A(n699), .ZN(n380) );
  XNOR2_X2 U534 ( .A(n466), .B(n353), .ZN(n699) );
  NOR2_X1 U535 ( .A1(n717), .A2(n382), .ZN(n381) );
  NAND2_X1 U536 ( .A1(n717), .A2(n387), .ZN(n386) );
  INV_X1 U537 ( .A(n388), .ZN(n399) );
  NAND2_X1 U538 ( .A1(n389), .A2(n390), .ZN(n388) );
  XNOR2_X1 U539 ( .A(n721), .B(n354), .ZN(n389) );
  XNOR2_X1 U540 ( .A(n647), .B(n355), .ZN(n391) );
  INV_X1 U541 ( .A(G134), .ZN(n481) );
  AND2_X2 U542 ( .A1(n722), .A2(G210), .ZN(n712) );
  XNOR2_X1 U543 ( .A(n395), .B(n561), .ZN(n433) );
  XNOR2_X1 U544 ( .A(n397), .B(n356), .ZN(n473) );
  NAND2_X1 U545 ( .A1(n722), .A2(G217), .ZN(n397) );
  NAND2_X1 U546 ( .A1(n727), .A2(n469), .ZN(n468) );
  XNOR2_X2 U547 ( .A(n635), .B(n634), .ZN(n727) );
  XNOR2_X1 U548 ( .A(n715), .B(n398), .ZN(n718) );
  XNOR2_X1 U549 ( .A(n717), .B(n716), .ZN(n398) );
  XNOR2_X1 U550 ( .A(n399), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U551 ( .A(n537), .B(n536), .ZN(n720) );
  XNOR2_X2 U552 ( .A(n404), .B(G110), .ZN(n521) );
  XNOR2_X2 U553 ( .A(n406), .B(G119), .ZN(n405) );
  NAND2_X1 U554 ( .A1(n407), .A2(n619), .ZN(n622) );
  NAND2_X1 U555 ( .A1(n407), .A2(n609), .ZN(n649) );
  NAND2_X1 U556 ( .A1(n412), .A2(n408), .ZN(n591) );
  INV_X1 U557 ( .A(n424), .ZN(n410) );
  INV_X1 U558 ( .A(n414), .ZN(n413) );
  NOR2_X1 U559 ( .A1(n424), .A2(KEYINPUT19), .ZN(n414) );
  NAND2_X1 U560 ( .A1(n417), .A2(n425), .ZN(n415) );
  INV_X1 U561 ( .A(n423), .ZN(n419) );
  NAND2_X1 U562 ( .A1(n710), .A2(n526), .ZN(n424) );
  XNOR2_X2 U563 ( .A(n542), .B(n426), .ZN(n739) );
  NAND2_X1 U564 ( .A1(n515), .A2(G134), .ZN(n428) );
  INV_X1 U565 ( .A(n515), .ZN(n430) );
  XNOR2_X1 U566 ( .A(n432), .B(n431), .ZN(n586) );
  INV_X1 U567 ( .A(KEYINPUT48), .ZN(n431) );
  NAND2_X1 U568 ( .A1(n434), .A2(n433), .ZN(n432) );
  INV_X1 U569 ( .A(n641), .ZN(n436) );
  NAND2_X1 U570 ( .A1(n563), .A2(n671), .ZN(n437) );
  XNOR2_X2 U571 ( .A(n440), .B(n351), .ZN(n570) );
  XNOR2_X1 U572 ( .A(n509), .B(n522), .ZN(n441) );
  XNOR2_X1 U573 ( .A(n442), .B(n706), .ZN(G75) );
  NAND2_X1 U574 ( .A1(n443), .A2(n460), .ZN(n442) );
  XNOR2_X1 U575 ( .A(n444), .B(KEYINPUT86), .ZN(n443) );
  INV_X1 U576 ( .A(n591), .ZN(n595) );
  NAND2_X1 U577 ( .A1(n649), .A2(n445), .ZN(n613) );
  INV_X1 U578 ( .A(n650), .ZN(n446) );
  NAND2_X1 U579 ( .A1(n449), .A2(n727), .ZN(n448) );
  INV_X1 U580 ( .A(n740), .ZN(n449) );
  XNOR2_X2 U581 ( .A(n451), .B(n450), .ZN(n515) );
  XNOR2_X2 U582 ( .A(G143), .B(G128), .ZN(n451) );
  NAND2_X1 U583 ( .A1(n581), .A2(n575), .ZN(n456) );
  INV_X1 U584 ( .A(n704), .ZN(n461) );
  INV_X1 U585 ( .A(n626), .ZN(n555) );
  INV_X1 U586 ( .A(n681), .ZN(n588) );
  INV_X1 U587 ( .A(n684), .ZN(n464) );
  INV_X1 U588 ( .A(KEYINPUT6), .ZN(n467) );
  NAND2_X1 U589 ( .A1(n468), .A2(n470), .ZN(n637) );
  XNOR2_X1 U590 ( .A(n485), .B(n521), .ZN(n471) );
  XNOR2_X2 U591 ( .A(n739), .B(n514), .ZN(n506) );
  OR2_X1 U592 ( .A1(n594), .A2(n593), .ZN(n472) );
  XNOR2_X1 U593 ( .A(KEYINPUT110), .B(n604), .ZN(n474) );
  INV_X1 U594 ( .A(KEYINPUT44), .ZN(n627) );
  INV_X1 U595 ( .A(KEYINPUT76), .ZN(n589) );
  XNOR2_X1 U596 ( .A(n494), .B(n493), .ZN(n495) );
  AND2_X1 U597 ( .A1(n573), .A2(n672), .ZN(n574) );
  XNOR2_X1 U598 ( .A(n710), .B(n709), .ZN(n711) );
  XNOR2_X1 U599 ( .A(n598), .B(KEYINPUT87), .ZN(n599) );
  XOR2_X1 U600 ( .A(KEYINPUT40), .B(KEYINPUT111), .Z(n552) );
  XNOR2_X1 U601 ( .A(n475), .B(KEYINPUT14), .ZN(n476) );
  XNOR2_X1 U602 ( .A(KEYINPUT74), .B(n476), .ZN(n478) );
  NAND2_X1 U603 ( .A1(G952), .A2(n478), .ZN(n698) );
  NOR2_X1 U604 ( .A1(G953), .A2(n698), .ZN(n477) );
  XOR2_X1 U605 ( .A(KEYINPUT93), .B(n477), .Z(n594) );
  AND2_X1 U606 ( .A1(n478), .A2(G953), .ZN(n479) );
  NAND2_X1 U607 ( .A1(G902), .A2(n479), .ZN(n592) );
  NOR2_X1 U608 ( .A1(G900), .A2(n592), .ZN(n480) );
  NOR2_X1 U609 ( .A1(n594), .A2(n480), .ZN(n556) );
  XOR2_X2 U610 ( .A(KEYINPUT71), .B(G101), .Z(n514) );
  NAND2_X1 U611 ( .A1(G227), .A2(n741), .ZN(n483) );
  XNOR2_X1 U612 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U613 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U614 ( .A(n535), .B(n488), .ZN(n496) );
  XOR2_X1 U615 ( .A(KEYINPUT23), .B(KEYINPUT95), .Z(n490) );
  XNOR2_X1 U616 ( .A(G119), .B(G137), .ZN(n489) );
  NAND2_X1 U617 ( .A1(G234), .A2(n741), .ZN(n491) );
  XNOR2_X1 U618 ( .A(n492), .B(n491), .ZN(n543) );
  NAND2_X1 U619 ( .A1(G221), .A2(n543), .ZN(n493) );
  NOR2_X1 U620 ( .A1(n643), .A2(G902), .ZN(n501) );
  XOR2_X1 U621 ( .A(KEYINPUT25), .B(KEYINPUT79), .Z(n499) );
  INV_X1 U622 ( .A(n524), .ZN(n636) );
  NAND2_X1 U623 ( .A1(G234), .A2(n636), .ZN(n497) );
  XNOR2_X1 U624 ( .A(KEYINPUT20), .B(n497), .ZN(n502) );
  NAND2_X1 U625 ( .A1(n502), .A2(G217), .ZN(n498) );
  XNOR2_X1 U626 ( .A(n499), .B(n498), .ZN(n500) );
  NAND2_X1 U627 ( .A1(n502), .A2(G221), .ZN(n503) );
  XNOR2_X1 U628 ( .A(KEYINPUT21), .B(n503), .ZN(n684) );
  NAND2_X1 U629 ( .A1(G214), .A2(n525), .ZN(n504) );
  XOR2_X1 U630 ( .A(KEYINPUT92), .B(n504), .Z(n572) );
  XNOR2_X2 U631 ( .A(G113), .B(G116), .ZN(n505) );
  XNOR2_X1 U632 ( .A(n507), .B(KEYINPUT78), .ZN(n533) );
  NAND2_X1 U633 ( .A1(n533), .A2(G210), .ZN(n508) );
  INV_X1 U634 ( .A(G472), .ZN(n510) );
  XNOR2_X1 U635 ( .A(KEYINPUT30), .B(n511), .ZN(n512) );
  XNOR2_X1 U636 ( .A(n514), .B(n513), .ZN(n516) );
  XNOR2_X1 U637 ( .A(n516), .B(n515), .ZN(n520) );
  XOR2_X1 U638 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n518) );
  NAND2_X1 U639 ( .A1(G224), .A2(n741), .ZN(n517) );
  XNOR2_X1 U640 ( .A(n518), .B(n517), .ZN(n519) );
  NAND2_X1 U641 ( .A1(G210), .A2(n525), .ZN(n526) );
  XNOR2_X1 U642 ( .A(n529), .B(n528), .ZN(n532) );
  NAND2_X1 U643 ( .A1(G214), .A2(n533), .ZN(n534) );
  XNOR2_X1 U644 ( .A(KEYINPUT100), .B(KEYINPUT13), .ZN(n538) );
  XNOR2_X1 U645 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U646 ( .A(n542), .B(n541), .Z(n549) );
  NAND2_X1 U647 ( .A1(G217), .A2(n543), .ZN(n547) );
  XNOR2_X1 U648 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U649 ( .A(KEYINPUT104), .B(KEYINPUT105), .ZN(n550) );
  INV_X1 U650 ( .A(n562), .ZN(n567) );
  INV_X1 U651 ( .A(n572), .ZN(n672) );
  NAND2_X1 U652 ( .A1(n672), .A2(n671), .ZN(n675) );
  NAND2_X1 U653 ( .A1(n566), .A2(n562), .ZN(n674) );
  XNOR2_X1 U654 ( .A(KEYINPUT112), .B(KEYINPUT41), .ZN(n553) );
  NOR2_X1 U655 ( .A1(n556), .A2(n684), .ZN(n557) );
  NAND2_X1 U656 ( .A1(n555), .A2(n557), .ZN(n571) );
  NOR2_X1 U657 ( .A1(n571), .A2(n570), .ZN(n558) );
  XOR2_X1 U658 ( .A(KEYINPUT28), .B(n558), .Z(n559) );
  NOR2_X1 U659 ( .A1(n700), .A2(n565), .ZN(n560) );
  XOR2_X1 U660 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n561) );
  NOR2_X1 U661 ( .A1(n566), .A2(n562), .ZN(n597) );
  NAND2_X1 U662 ( .A1(n563), .A2(n597), .ZN(n564) );
  NOR2_X1 U663 ( .A1(n584), .A2(n564), .ZN(n660) );
  OR2_X1 U664 ( .A1(n565), .A2(n591), .ZN(n661) );
  NAND2_X1 U665 ( .A1(n567), .A2(n566), .ZN(n657) );
  INV_X1 U666 ( .A(n657), .ZN(n602) );
  NOR2_X1 U667 ( .A1(n602), .A2(n611), .ZN(n676) );
  XOR2_X1 U668 ( .A(KEYINPUT47), .B(n568), .Z(n569) );
  INV_X1 U669 ( .A(n571), .ZN(n573) );
  INV_X1 U670 ( .A(KEYINPUT69), .ZN(n577) );
  INV_X1 U671 ( .A(KEYINPUT1), .ZN(n576) );
  INV_X1 U672 ( .A(n617), .ZN(n682) );
  XOR2_X1 U673 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n583) );
  NAND2_X1 U674 ( .A1(n682), .A2(n581), .ZN(n582) );
  XNOR2_X1 U675 ( .A(n583), .B(n582), .ZN(n585) );
  NAND2_X1 U676 ( .A1(n585), .A2(n584), .ZN(n670) );
  NAND2_X1 U677 ( .A1(n586), .A2(n670), .ZN(n641) );
  NAND2_X1 U678 ( .A1(n587), .A2(n602), .ZN(n669) );
  NOR2_X1 U679 ( .A1(G898), .A2(n592), .ZN(n593) );
  NAND2_X1 U680 ( .A1(n595), .A2(n472), .ZN(n596) );
  XNOR2_X2 U681 ( .A(n596), .B(KEYINPUT0), .ZN(n605) );
  XOR2_X1 U682 ( .A(KEYINPUT35), .B(KEYINPUT80), .Z(n598) );
  NAND2_X1 U683 ( .A1(n628), .A2(KEYINPUT44), .ZN(n615) );
  AND2_X1 U684 ( .A1(n602), .A2(n612), .ZN(n666) );
  INV_X1 U685 ( .A(n611), .ZN(n662) );
  NOR2_X1 U686 ( .A1(n362), .A2(n605), .ZN(n603) );
  NAND2_X1 U687 ( .A1(n604), .A2(n603), .ZN(n610) );
  NOR2_X1 U688 ( .A1(n662), .A2(n610), .ZN(n650) );
  INV_X1 U689 ( .A(n674), .ZN(n607) );
  NOR2_X1 U690 ( .A1(n555), .A2(n454), .ZN(n609) );
  OR2_X1 U691 ( .A1(n657), .A2(n610), .ZN(n653) );
  NAND2_X1 U692 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U693 ( .A(n616), .B(KEYINPUT89), .ZN(n633) );
  NAND2_X1 U694 ( .A1(n555), .A2(n454), .ZN(n618) );
  XNOR2_X1 U695 ( .A(KEYINPUT107), .B(n618), .ZN(n619) );
  XNOR2_X1 U696 ( .A(KEYINPUT81), .B(KEYINPUT68), .ZN(n620) );
  XNOR2_X1 U697 ( .A(n620), .B(KEYINPUT32), .ZN(n621) );
  XNOR2_X1 U698 ( .A(n622), .B(n621), .ZN(n749) );
  NOR2_X1 U699 ( .A1(n362), .A2(n623), .ZN(n624) );
  NAND2_X1 U700 ( .A1(n682), .A2(n624), .ZN(n625) );
  NOR2_X2 U701 ( .A1(n749), .A2(n655), .ZN(n629) );
  XNOR2_X1 U702 ( .A(n629), .B(n627), .ZN(n631) );
  NAND2_X1 U703 ( .A1(n629), .A2(n750), .ZN(n630) );
  NAND2_X1 U704 ( .A1(n631), .A2(n630), .ZN(n632) );
  NAND2_X1 U705 ( .A1(n633), .A2(n632), .ZN(n635) );
  XOR2_X1 U706 ( .A(KEYINPUT45), .B(KEYINPUT65), .Z(n634) );
  XNOR2_X1 U707 ( .A(n637), .B(KEYINPUT67), .ZN(n642) );
  NAND2_X1 U708 ( .A1(KEYINPUT2), .A2(n669), .ZN(n638) );
  XOR2_X1 U709 ( .A(KEYINPUT82), .B(n638), .Z(n639) );
  NAND2_X1 U710 ( .A1(n727), .A2(n639), .ZN(n640) );
  NOR2_X1 U711 ( .A1(n641), .A2(n640), .ZN(n704) );
  NOR2_X2 U712 ( .A1(n642), .A2(n704), .ZN(n722) );
  NAND2_X1 U713 ( .A1(n473), .A2(n390), .ZN(n644) );
  XNOR2_X1 U714 ( .A(n644), .B(KEYINPUT125), .ZN(G66) );
  NAND2_X1 U715 ( .A1(n722), .A2(G472), .ZN(n647) );
  XOR2_X1 U716 ( .A(KEYINPUT62), .B(KEYINPUT91), .Z(n645) );
  INV_X1 U717 ( .A(KEYINPUT63), .ZN(n648) );
  XNOR2_X1 U718 ( .A(n349), .B(n648), .ZN(G57) );
  XNOR2_X1 U719 ( .A(G101), .B(n649), .ZN(G3) );
  XOR2_X1 U720 ( .A(G104), .B(n650), .Z(G6) );
  XOR2_X1 U721 ( .A(KEYINPUT27), .B(KEYINPUT115), .Z(n652) );
  XNOR2_X1 U722 ( .A(G107), .B(KEYINPUT26), .ZN(n651) );
  XNOR2_X1 U723 ( .A(n652), .B(n651), .ZN(n654) );
  XOR2_X1 U724 ( .A(n654), .B(n653), .Z(G9) );
  XOR2_X1 U725 ( .A(G110), .B(n655), .Z(n656) );
  XNOR2_X1 U726 ( .A(KEYINPUT116), .B(n656), .ZN(G12) );
  NOR2_X1 U727 ( .A1(n657), .A2(n661), .ZN(n659) );
  XNOR2_X1 U728 ( .A(n392), .B(KEYINPUT29), .ZN(n658) );
  XNOR2_X1 U729 ( .A(n659), .B(n658), .ZN(G30) );
  XOR2_X1 U730 ( .A(G143), .B(n660), .Z(G45) );
  NOR2_X1 U731 ( .A1(n662), .A2(n661), .ZN(n663) );
  XOR2_X1 U732 ( .A(G146), .B(n663), .Z(G48) );
  XOR2_X1 U733 ( .A(G113), .B(KEYINPUT117), .Z(n664) );
  XNOR2_X1 U734 ( .A(n665), .B(n664), .ZN(G15) );
  XOR2_X1 U735 ( .A(G116), .B(n666), .Z(n667) );
  XNOR2_X1 U736 ( .A(KEYINPUT118), .B(n667), .ZN(G18) );
  XOR2_X1 U737 ( .A(G134), .B(KEYINPUT119), .Z(n668) );
  XNOR2_X1 U738 ( .A(n669), .B(n668), .ZN(G36) );
  XNOR2_X1 U739 ( .A(G140), .B(n670), .ZN(G42) );
  XOR2_X1 U740 ( .A(KEYINPUT53), .B(KEYINPUT122), .Z(n706) );
  NOR2_X1 U741 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U742 ( .A1(n674), .A2(n673), .ZN(n679) );
  NOR2_X1 U743 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U744 ( .A(n677), .B(KEYINPUT120), .ZN(n678) );
  NOR2_X1 U745 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U746 ( .A1(n396), .A2(n680), .ZN(n695) );
  NAND2_X1 U747 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U748 ( .A(n683), .B(KEYINPUT50), .ZN(n689) );
  AND2_X1 U749 ( .A1(n684), .A2(n555), .ZN(n685) );
  XOR2_X1 U750 ( .A(KEYINPUT49), .B(n685), .Z(n686) );
  NOR2_X1 U751 ( .A1(n362), .A2(n686), .ZN(n688) );
  NAND2_X1 U752 ( .A1(n689), .A2(n688), .ZN(n691) );
  NAND2_X1 U753 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U754 ( .A(KEYINPUT51), .B(n692), .ZN(n693) );
  NOR2_X1 U755 ( .A1(n346), .A2(n693), .ZN(n694) );
  NOR2_X1 U756 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U757 ( .A(n696), .B(KEYINPUT52), .ZN(n697) );
  NOR2_X1 U758 ( .A1(n698), .A2(n697), .ZN(n702) );
  NOR2_X1 U759 ( .A1(n346), .A2(n396), .ZN(n701) );
  NOR2_X1 U760 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U761 ( .A(KEYINPUT121), .B(n703), .ZN(n705) );
  XOR2_X1 U762 ( .A(KEYINPUT54), .B(KEYINPUT123), .Z(n708) );
  XNOR2_X1 U763 ( .A(KEYINPUT90), .B(KEYINPUT55), .ZN(n707) );
  XNOR2_X1 U764 ( .A(n708), .B(n707), .ZN(n709) );
  XNOR2_X1 U765 ( .A(n712), .B(n711), .ZN(n713) );
  NOR2_X1 U766 ( .A1(n713), .A2(n726), .ZN(n714) );
  XNOR2_X1 U767 ( .A(n714), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U768 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n716) );
  NAND2_X1 U769 ( .A1(n722), .A2(G469), .ZN(n715) );
  NOR2_X1 U770 ( .A1(n726), .A2(n718), .ZN(G54) );
  NAND2_X1 U771 ( .A1(n722), .A2(G475), .ZN(n721) );
  XOR2_X1 U772 ( .A(KEYINPUT59), .B(KEYINPUT70), .Z(n719) );
  NAND2_X1 U773 ( .A1(G478), .A2(n722), .ZN(n723) );
  XNOR2_X1 U774 ( .A(n724), .B(n723), .ZN(n725) );
  NOR2_X1 U775 ( .A1(n726), .A2(n725), .ZN(G63) );
  NAND2_X1 U776 ( .A1(n741), .A2(n727), .ZN(n731) );
  NAND2_X1 U777 ( .A1(G953), .A2(G224), .ZN(n728) );
  XNOR2_X1 U778 ( .A(KEYINPUT61), .B(n728), .ZN(n729) );
  NAND2_X1 U779 ( .A1(n729), .A2(G898), .ZN(n730) );
  NAND2_X1 U780 ( .A1(n731), .A2(n730), .ZN(n736) );
  XNOR2_X1 U781 ( .A(n732), .B(G101), .ZN(n734) );
  NOR2_X1 U782 ( .A1(n741), .A2(G898), .ZN(n733) );
  NOR2_X1 U783 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U784 ( .A(n736), .B(n735), .ZN(n737) );
  XNOR2_X1 U785 ( .A(KEYINPUT126), .B(n737), .ZN(G69) );
  XNOR2_X1 U786 ( .A(n739), .B(n738), .ZN(n743) );
  XOR2_X1 U787 ( .A(n743), .B(n740), .Z(n742) );
  NAND2_X1 U788 ( .A1(n742), .A2(n741), .ZN(n748) );
  XNOR2_X1 U789 ( .A(G227), .B(n743), .ZN(n744) );
  XNOR2_X1 U790 ( .A(n744), .B(KEYINPUT127), .ZN(n745) );
  NAND2_X1 U791 ( .A1(n745), .A2(G900), .ZN(n746) );
  NAND2_X1 U792 ( .A1(G953), .A2(n746), .ZN(n747) );
  NAND2_X1 U793 ( .A1(n748), .A2(n747), .ZN(G72) );
  XOR2_X1 U794 ( .A(n749), .B(G119), .Z(G21) );
  XOR2_X1 U795 ( .A(n750), .B(G122), .Z(G24) );
  XNOR2_X1 U796 ( .A(G125), .B(KEYINPUT37), .ZN(n751) );
  XNOR2_X1 U797 ( .A(n752), .B(G131), .ZN(G33) );
  XNOR2_X1 U798 ( .A(n753), .B(G137), .ZN(G39) );
endmodule

