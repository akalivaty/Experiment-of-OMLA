//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 0 1 1 0 1 1 1 0 1 1 0 0 1 1 1 1 1 0 1 1 0 0 1 1 0 1 0 0 1 1 1 0 1 0 0 0 1 1 1 0 1 1 0 1 1 1 1 1 1 0 1 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n868, new_n869, new_n870,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n978, new_n979;
  XOR2_X1   g000(.A(G78gat), .B(G106gat), .Z(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT84), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT31), .B(G50gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G228gat), .A2(G233gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208));
  AND2_X1   g007(.A1(KEYINPUT74), .A2(KEYINPUT2), .ZN(new_n209));
  NOR2_X1   g008(.A1(KEYINPUT74), .A2(KEYINPUT2), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT75), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  OAI211_X1 g012(.A(KEYINPUT75), .B(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n214));
  INV_X1    g013(.A(G148gat), .ZN(new_n215));
  OR2_X1    g014(.A1(new_n215), .A2(G141gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(G141gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n213), .A2(new_n214), .A3(new_n218), .ZN(new_n219));
  AND2_X1   g018(.A1(G155gat), .A2(G162gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(G155gat), .A2(G162gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT73), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(KEYINPUT73), .B1(G155gat), .B2(G162gat), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n220), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT77), .B1(new_n220), .B2(new_n221), .ZN(new_n226));
  INV_X1    g025(.A(G155gat), .ZN(new_n227));
  INV_X1    g026(.A(G162gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT77), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n229), .A2(new_n230), .A3(new_n208), .ZN(new_n231));
  AOI22_X1  g030(.A1(new_n226), .A2(new_n231), .B1(KEYINPUT2), .B2(new_n208), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n215), .A2(KEYINPUT76), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT76), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(G148gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n233), .A2(new_n235), .A3(G141gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(new_n216), .ZN(new_n237));
  AOI22_X1  g036(.A1(new_n219), .A2(new_n225), .B1(new_n232), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G211gat), .ZN(new_n239));
  INV_X1    g038(.A(G218gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(G211gat), .A2(G218gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(KEYINPUT70), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT70), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n241), .A2(new_n245), .A3(new_n242), .ZN(new_n246));
  AND2_X1   g045(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(G197gat), .ZN(new_n248));
  INV_X1    g047(.A(G204gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(G197gat), .A2(G204gat), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT22), .ZN(new_n252));
  AOI22_X1  g051(.A1(new_n250), .A2(new_n251), .B1(new_n252), .B2(new_n242), .ZN(new_n253));
  AOI21_X1  g052(.A(KEYINPUT29), .B1(new_n247), .B2(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n254), .B1(new_n247), .B2(new_n253), .ZN(new_n255));
  XOR2_X1   g054(.A(KEYINPUT78), .B(KEYINPUT3), .Z(new_n256));
  AOI21_X1  g055(.A(new_n238), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT69), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n244), .A2(new_n258), .A3(new_n246), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n259), .B(new_n253), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n238), .A2(new_n256), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT29), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n207), .B1(new_n257), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(KEYINPUT85), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n219), .A2(new_n225), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n226), .A2(new_n231), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n208), .A2(KEYINPUT2), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n268), .A2(new_n237), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n207), .B1(new_n271), .B2(KEYINPUT3), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n260), .A2(new_n262), .A3(new_n271), .ZN(new_n273));
  OAI211_X1 g072(.A(new_n272), .B(new_n273), .C1(new_n263), .C2(KEYINPUT85), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n264), .B1(new_n266), .B2(new_n274), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n275), .A2(G22gat), .ZN(new_n276));
  INV_X1    g075(.A(G22gat), .ZN(new_n277));
  OR2_X1    g076(.A1(new_n263), .A2(KEYINPUT85), .ZN(new_n278));
  AND2_X1   g077(.A1(new_n273), .A2(new_n272), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n278), .A2(new_n279), .A3(new_n265), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n277), .B1(new_n280), .B2(new_n264), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n206), .B1(new_n276), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n275), .A2(G22gat), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n280), .A2(new_n277), .A3(new_n264), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n283), .A2(new_n284), .A3(new_n205), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT32), .ZN(new_n287));
  XNOR2_X1  g086(.A(G127gat), .B(G134gat), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(G113gat), .B(G120gat), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n289), .B1(KEYINPUT1), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n290), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT1), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n292), .A2(new_n288), .A3(new_n293), .ZN(new_n294));
  AND2_X1   g093(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT24), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n297), .A2(G183gat), .A3(G190gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(G183gat), .B(G190gat), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n298), .B1(new_n299), .B2(new_n297), .ZN(new_n300));
  INV_X1    g099(.A(G169gat), .ZN(new_n301));
  INV_X1    g100(.A(G176gat), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n301), .A2(new_n302), .A3(KEYINPUT23), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT23), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n304), .B1(G169gat), .B2(G176gat), .ZN(new_n305));
  NOR2_X1   g104(.A1(G169gat), .A2(G176gat), .ZN(new_n306));
  OAI211_X1 g105(.A(KEYINPUT25), .B(new_n303), .C1(new_n305), .C2(new_n306), .ZN(new_n307));
  OAI21_X1  g106(.A(KEYINPUT65), .B1(new_n300), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(G169gat), .A2(G176gat), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n306), .B1(KEYINPUT23), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n303), .A2(KEYINPUT25), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT65), .ZN(new_n313));
  AND3_X1   g112(.A1(new_n297), .A2(G183gat), .A3(G190gat), .ZN(new_n314));
  INV_X1    g113(.A(G183gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(G190gat), .ZN(new_n316));
  INV_X1    g115(.A(G190gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G183gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n314), .B1(new_n319), .B2(KEYINPUT24), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n312), .A2(new_n313), .A3(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n310), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n301), .A2(KEYINPUT64), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT64), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(G169gat), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n323), .A2(new_n325), .A3(KEYINPUT23), .A4(new_n302), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n320), .A2(new_n322), .A3(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT25), .ZN(new_n328));
  AOI22_X1  g127(.A1(new_n308), .A2(new_n321), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n315), .A2(KEYINPUT27), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT27), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(G183gat), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n330), .A2(new_n332), .A3(new_n317), .ZN(new_n333));
  AOI22_X1  g132(.A1(new_n333), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n306), .A2(KEYINPUT66), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(KEYINPUT26), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT26), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n306), .A2(KEYINPUT66), .A3(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n336), .A2(new_n309), .A3(new_n338), .ZN(new_n339));
  AND2_X1   g138(.A1(new_n330), .A2(new_n332), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT28), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n340), .A2(new_n341), .A3(new_n317), .ZN(new_n342));
  AND3_X1   g141(.A1(new_n334), .A2(new_n339), .A3(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n296), .B1(new_n329), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n322), .A2(new_n326), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n328), .B1(new_n345), .B2(new_n300), .ZN(new_n346));
  NOR3_X1   g145(.A1(new_n300), .A2(new_n307), .A3(KEYINPUT65), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n313), .B1(new_n312), .B2(new_n320), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n346), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n343), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n349), .A2(new_n295), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n344), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(G227gat), .ZN(new_n353));
  INV_X1    g152(.A(G233gat), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n287), .B1(new_n352), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n352), .A2(new_n355), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT33), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  XOR2_X1   g159(.A(G71gat), .B(G99gat), .Z(new_n361));
  XNOR2_X1  g160(.A(G15gat), .B(G43gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n361), .B(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n357), .A2(new_n360), .A3(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n352), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT68), .ZN(new_n366));
  INV_X1    g165(.A(new_n355), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n365), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT67), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n363), .A2(KEYINPUT33), .ZN(new_n370));
  AND4_X1   g169(.A1(new_n369), .A2(new_n358), .A3(KEYINPUT32), .A4(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n369), .B1(new_n356), .B2(new_n370), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n364), .B(new_n368), .C1(new_n371), .C2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n358), .A2(KEYINPUT32), .A3(new_n370), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT67), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n356), .A2(new_n369), .A3(new_n370), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n368), .B1(new_n378), .B2(new_n364), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n366), .B1(new_n365), .B2(new_n367), .ZN(new_n380));
  OAI22_X1  g179(.A1(new_n374), .A2(new_n379), .B1(KEYINPUT34), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n364), .B1(new_n371), .B2(new_n372), .ZN(new_n382));
  INV_X1    g181(.A(new_n368), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n380), .A2(KEYINPUT34), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n384), .A2(new_n373), .A3(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n286), .B1(new_n381), .B2(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(G8gat), .B(G36gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(G64gat), .B(G92gat), .ZN(new_n389));
  XOR2_X1   g188(.A(new_n388), .B(new_n389), .Z(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(G226gat), .A2(G233gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n308), .A2(new_n321), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n343), .B1(new_n393), .B2(new_n346), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n392), .B1(new_n394), .B2(KEYINPUT29), .ZN(new_n395));
  INV_X1    g194(.A(new_n392), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n396), .B1(new_n329), .B2(new_n343), .ZN(new_n397));
  AND3_X1   g196(.A1(new_n395), .A2(new_n260), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n260), .B1(new_n395), .B2(new_n397), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n391), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT29), .B1(new_n349), .B2(new_n350), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n397), .B1(new_n401), .B2(new_n396), .ZN(new_n402));
  INV_X1    g201(.A(new_n260), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n395), .A2(new_n260), .A3(new_n397), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n404), .A2(KEYINPUT30), .A3(new_n390), .A4(new_n405), .ZN(new_n406));
  AND3_X1   g205(.A1(new_n400), .A2(new_n406), .A3(KEYINPUT71), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT71), .B1(new_n400), .B2(new_n406), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n404), .A2(new_n390), .A3(new_n405), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT30), .ZN(new_n410));
  AND3_X1   g209(.A1(new_n409), .A2(KEYINPUT72), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT72), .B1(new_n409), .B2(new_n410), .ZN(new_n412));
  OAI22_X1  g211(.A1(new_n407), .A2(new_n408), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT79), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT3), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n296), .B1(new_n238), .B2(new_n415), .ZN(new_n416));
  AND3_X1   g215(.A1(new_n267), .A2(new_n270), .A3(new_n256), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n414), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n225), .ZN(new_n419));
  AOI22_X1  g218(.A1(new_n211), .A2(new_n212), .B1(new_n216), .B2(new_n217), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n419), .B1(new_n420), .B2(new_n214), .ZN(new_n421));
  INV_X1    g220(.A(new_n270), .ZN(new_n422));
  OAI21_X1  g221(.A(KEYINPUT3), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n423), .A2(new_n261), .A3(KEYINPUT79), .A4(new_n296), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n418), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n270), .A2(new_n294), .A3(new_n291), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n426), .A2(new_n421), .ZN(new_n427));
  XNOR2_X1  g226(.A(KEYINPUT80), .B(KEYINPUT4), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT81), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n430), .B1(new_n426), .B2(new_n421), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n295), .A2(new_n267), .A3(KEYINPUT81), .A4(new_n270), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT4), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n429), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n425), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(G225gat), .A2(G233gat), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  NOR3_X1   g237(.A1(new_n436), .A2(KEYINPUT5), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n433), .A2(new_n434), .ZN(new_n441));
  OR2_X1    g240(.A1(new_n427), .A2(new_n428), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n443), .A2(new_n425), .A3(new_n437), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT5), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT82), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n271), .A2(new_n296), .A3(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(KEYINPUT82), .B1(new_n238), .B2(new_n295), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n449), .A2(new_n431), .A3(new_n432), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n445), .B1(new_n450), .B2(new_n438), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT83), .ZN(new_n452));
  AND3_X1   g251(.A1(new_n444), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n452), .B1(new_n444), .B2(new_n451), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n440), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  XNOR2_X1  g254(.A(G1gat), .B(G29gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n456), .B(KEYINPUT0), .ZN(new_n457));
  XNOR2_X1  g256(.A(G57gat), .B(G85gat), .ZN(new_n458));
  XOR2_X1   g257(.A(new_n457), .B(new_n458), .Z(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(KEYINPUT6), .ZN(new_n460));
  INV_X1    g259(.A(new_n459), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT6), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n455), .A2(new_n460), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n444), .A2(new_n451), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(KEYINPUT83), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n444), .A2(new_n451), .A3(new_n452), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n468), .A2(new_n462), .A3(new_n440), .A4(new_n461), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n413), .B1(new_n464), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n387), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT35), .ZN(new_n472));
  AND2_X1   g271(.A1(new_n400), .A2(new_n406), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n473), .B1(new_n411), .B2(new_n412), .ZN(new_n474));
  AOI211_X1 g273(.A(new_n286), .B(new_n474), .C1(new_n381), .C2(new_n386), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n464), .A2(new_n469), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n476), .A2(KEYINPUT35), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n472), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n381), .A2(new_n386), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT36), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n381), .A2(KEYINPUT36), .A3(new_n386), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n464), .A2(new_n469), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT37), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n404), .A2(new_n486), .A3(new_n405), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT88), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT88), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n404), .A2(new_n489), .A3(new_n486), .A4(new_n405), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  OAI211_X1 g290(.A(KEYINPUT87), .B(KEYINPUT37), .C1(new_n398), .C2(new_n399), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT38), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n391), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(KEYINPUT37), .B1(new_n398), .B2(new_n399), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT87), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n491), .A2(new_n492), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n495), .A2(new_n391), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n499), .B1(new_n488), .B2(new_n490), .ZN(new_n500));
  OAI211_X1 g299(.A(new_n498), .B(new_n409), .C1(new_n500), .C2(new_n493), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n485), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n286), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n439), .B1(new_n466), .B2(new_n467), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n474), .B1(new_n504), .B2(new_n459), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n437), .B1(new_n425), .B2(new_n435), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT39), .ZN(new_n508));
  INV_X1    g307(.A(new_n450), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n508), .B1(new_n509), .B2(new_n437), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n461), .B1(new_n506), .B2(new_n508), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT40), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n511), .A2(new_n512), .A3(KEYINPUT40), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n503), .B1(new_n505), .B2(new_n517), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n282), .A2(KEYINPUT86), .A3(new_n285), .ZN(new_n519));
  AOI21_X1  g318(.A(KEYINPUT86), .B1(new_n282), .B2(new_n285), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI22_X1  g320(.A1(new_n502), .A2(new_n518), .B1(new_n470), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n479), .B1(new_n484), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(G29gat), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n524), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n525));
  XOR2_X1   g324(.A(KEYINPUT14), .B(G29gat), .Z(new_n526));
  OAI21_X1  g325(.A(new_n525), .B1(new_n526), .B2(G36gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(G43gat), .B(G50gat), .ZN(new_n528));
  AOI22_X1  g327(.A1(new_n527), .A2(KEYINPUT90), .B1(KEYINPUT15), .B2(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n527), .B1(KEYINPUT15), .B2(new_n528), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(G15gat), .B(G22gat), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT16), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n533), .B1(new_n534), .B2(G1gat), .ZN(new_n535));
  INV_X1    g334(.A(G8gat), .ZN(new_n536));
  OAI221_X1 g335(.A(new_n535), .B1(KEYINPUT91), .B2(new_n536), .C1(G1gat), .C2(new_n533), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(KEYINPUT91), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  OR2_X1    g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n537), .A2(new_n539), .ZN(new_n541));
  AND3_X1   g340(.A1(new_n540), .A2(KEYINPUT92), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g341(.A(KEYINPUT92), .B1(new_n540), .B2(new_n541), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n532), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n540), .A2(new_n541), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT92), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n540), .A2(KEYINPUT92), .A3(new_n541), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n547), .A2(new_n531), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n544), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(G229gat), .A2(G233gat), .ZN(new_n551));
  XOR2_X1   g350(.A(new_n551), .B(KEYINPUT13), .Z(new_n552));
  NAND2_X1  g351(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT93), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n550), .A2(KEYINPUT93), .A3(new_n552), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT18), .ZN(new_n557));
  AND2_X1   g356(.A1(new_n531), .A2(KEYINPUT17), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n545), .B1(new_n531), .B2(KEYINPUT17), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n544), .B(new_n551), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  AOI22_X1  g359(.A1(new_n555), .A2(new_n556), .B1(new_n557), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT94), .ZN(new_n562));
  OR2_X1    g361(.A1(new_n558), .A2(new_n559), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n563), .A2(KEYINPUT18), .A3(new_n551), .A4(new_n544), .ZN(new_n564));
  XOR2_X1   g363(.A(G113gat), .B(G141gat), .Z(new_n565));
  XNOR2_X1  g364(.A(G169gat), .B(G197gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n565), .B(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n568));
  XOR2_X1   g367(.A(new_n567), .B(new_n568), .Z(new_n569));
  XOR2_X1   g368(.A(new_n569), .B(KEYINPUT12), .Z(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n561), .A2(new_n562), .A3(new_n564), .A4(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n560), .A2(new_n557), .ZN(new_n573));
  AOI21_X1  g372(.A(KEYINPUT93), .B1(new_n550), .B2(new_n552), .ZN(new_n574));
  INV_X1    g373(.A(new_n552), .ZN(new_n575));
  AOI211_X1 g374(.A(new_n554), .B(new_n575), .C1(new_n544), .C2(new_n549), .ZN(new_n576));
  OAI211_X1 g375(.A(new_n564), .B(new_n573), .C1(new_n574), .C2(new_n576), .ZN(new_n577));
  OAI21_X1  g376(.A(KEYINPUT94), .B1(new_n577), .B2(new_n570), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n572), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n570), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AND2_X1   g380(.A1(new_n523), .A2(new_n581), .ZN(new_n582));
  OR2_X1    g381(.A1(G57gat), .A2(G64gat), .ZN(new_n583));
  NAND2_X1  g382(.A1(G57gat), .A2(G64gat), .ZN(new_n584));
  AND2_X1   g383(.A1(G71gat), .A2(G78gat), .ZN(new_n585));
  OAI211_X1 g384(.A(new_n583), .B(new_n584), .C1(new_n585), .C2(KEYINPUT9), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT95), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g387(.A1(G71gat), .A2(G78gat), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n588), .B(new_n590), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n591), .A2(KEYINPUT21), .ZN(new_n592));
  NAND2_X1  g391(.A1(G231gat), .A2(G233gat), .ZN(new_n593));
  XOR2_X1   g392(.A(new_n592), .B(new_n593), .Z(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(G127gat), .ZN(new_n595));
  AOI211_X1 g394(.A(new_n543), .B(new_n542), .C1(KEYINPUT21), .C2(new_n591), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(G155gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(G183gat), .B(G211gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  OR2_X1    g400(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n597), .A2(new_n601), .ZN(new_n603));
  AND2_X1   g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n605));
  NAND2_X1  g404(.A1(G85gat), .A2(G92gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(KEYINPUT7), .ZN(new_n607));
  NOR2_X1   g406(.A1(G85gat), .A2(G92gat), .ZN(new_n608));
  NAND2_X1  g407(.A1(G99gat), .A2(G106gat), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n608), .B1(KEYINPUT8), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G99gat), .B(G106gat), .ZN(new_n612));
  XOR2_X1   g411(.A(new_n611), .B(new_n612), .Z(new_n613));
  OAI21_X1  g412(.A(new_n605), .B1(new_n531), .B2(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(KEYINPUT96), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n613), .B1(new_n531), .B2(KEYINPUT17), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n615), .B1(new_n558), .B2(new_n616), .ZN(new_n617));
  XOR2_X1   g416(.A(G190gat), .B(G218gat), .Z(new_n618));
  OR2_X1    g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(G134gat), .B(G162gat), .ZN(new_n620));
  AOI21_X1  g419(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n617), .A2(new_n618), .ZN(new_n623));
  AND3_X1   g422(.A1(new_n619), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n622), .B1(new_n619), .B2(new_n623), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n604), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n590), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n588), .B(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n613), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n611), .B(new_n612), .ZN(new_n631));
  OAI21_X1  g430(.A(KEYINPUT97), .B1(new_n631), .B2(new_n591), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n630), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(G230gat), .A2(G233gat), .ZN(new_n634));
  OR2_X1    g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT10), .ZN(new_n636));
  NOR3_X1   g435(.A1(new_n613), .A2(new_n636), .A3(new_n629), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n637), .B1(new_n633), .B2(new_n636), .ZN(new_n638));
  XOR2_X1   g437(.A(new_n634), .B(KEYINPUT98), .Z(new_n639));
  OAI21_X1  g438(.A(new_n635), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(G120gat), .B(G148gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(G176gat), .B(G204gat), .ZN(new_n642));
  XOR2_X1   g441(.A(new_n641), .B(new_n642), .Z(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  OR2_X1    g444(.A1(new_n630), .A2(new_n632), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n632), .ZN(new_n647));
  AOI21_X1  g446(.A(KEYINPUT10), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n634), .B1(new_n648), .B2(new_n637), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n649), .A2(new_n635), .A3(new_n643), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n645), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n582), .A2(new_n627), .A3(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n653), .A2(new_n485), .ZN(new_n654));
  XOR2_X1   g453(.A(new_n654), .B(G1gat), .Z(G1324gat));
  INV_X1    g454(.A(new_n474), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g456(.A(KEYINPUT16), .B(G8gat), .Z(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n659), .B1(new_n536), .B2(new_n657), .ZN(new_n660));
  MUX2_X1   g459(.A(new_n659), .B(new_n660), .S(KEYINPUT42), .Z(G1325gat));
  AND3_X1   g460(.A1(new_n381), .A2(KEYINPUT36), .A3(new_n386), .ZN(new_n662));
  AOI21_X1  g461(.A(KEYINPUT36), .B1(new_n381), .B2(new_n386), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(G15gat), .B1(new_n653), .B2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n480), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n666), .A2(G15gat), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n665), .B1(new_n653), .B2(new_n667), .ZN(G1326gat));
  NOR2_X1   g467(.A1(new_n653), .A2(new_n521), .ZN(new_n669));
  XOR2_X1   g468(.A(KEYINPUT43), .B(G22gat), .Z(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(G1327gat));
  NAND2_X1  g470(.A1(new_n602), .A2(new_n603), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n672), .A2(new_n651), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(new_n626), .ZN(new_n674));
  XOR2_X1   g473(.A(new_n674), .B(KEYINPUT99), .Z(new_n675));
  NAND2_X1  g474(.A1(new_n582), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n677), .A2(new_n524), .A3(new_n476), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(KEYINPUT45), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT44), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n680), .B1(new_n523), .B2(new_n626), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n626), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT102), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n684), .B1(new_n522), .B2(new_n484), .ZN(new_n685));
  INV_X1    g484(.A(new_n412), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n409), .A2(KEYINPUT72), .A3(new_n410), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  AOI22_X1  g487(.A1(new_n688), .A2(new_n473), .B1(new_n455), .B2(new_n461), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n515), .A2(new_n516), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n286), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n409), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n491), .A2(new_n391), .A3(new_n495), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n692), .B1(new_n693), .B2(KEYINPUT38), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n694), .A2(new_n469), .A3(new_n464), .A4(new_n498), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n413), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n485), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n520), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n282), .A2(KEYINPUT86), .A3(new_n285), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n664), .A2(KEYINPUT102), .A3(new_n696), .A4(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n685), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n683), .B1(new_n704), .B2(new_n479), .ZN(new_n705));
  AOI21_X1  g504(.A(KEYINPUT103), .B1(new_n705), .B2(new_n680), .ZN(new_n706));
  AOI22_X1  g505(.A1(KEYINPUT35), .A2(new_n471), .B1(new_n475), .B2(new_n477), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n707), .B1(new_n685), .B2(new_n703), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT103), .ZN(new_n709));
  NOR4_X1   g508(.A1(new_n708), .A2(new_n709), .A3(KEYINPUT44), .A4(new_n683), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n682), .B1(new_n706), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n581), .A2(KEYINPUT100), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT100), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n579), .A2(new_n713), .A3(new_n580), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(new_n673), .ZN(new_n717));
  XOR2_X1   g516(.A(new_n717), .B(KEYINPUT101), .Z(new_n718));
  NAND2_X1  g517(.A1(new_n711), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(G29gat), .B1(new_n719), .B2(new_n485), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n679), .A2(new_n720), .ZN(G1328gat));
  AOI21_X1  g520(.A(G36gat), .B1(KEYINPUT104), .B2(KEYINPUT46), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n677), .A2(new_n474), .A3(new_n722), .ZN(new_n723));
  NOR2_X1   g522(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n723), .B(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(G36gat), .B1(new_n719), .B2(new_n656), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(G1329gat));
  NOR3_X1   g526(.A1(new_n676), .A2(G43gat), .A3(new_n666), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n711), .A2(new_n484), .A3(new_n718), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n728), .B1(new_n729), .B2(G43gat), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g530(.A(G50gat), .ZN(new_n732));
  INV_X1    g531(.A(new_n719), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n732), .B1(new_n733), .B2(new_n286), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n732), .B(new_n701), .C1(new_n676), .C2(KEYINPUT105), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n676), .A2(KEYINPUT105), .ZN(new_n736));
  OAI21_X1  g535(.A(KEYINPUT48), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n735), .A2(new_n736), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n711), .A2(new_n701), .A3(new_n718), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n738), .B1(new_n739), .B2(G50gat), .ZN(new_n740));
  OAI22_X1  g539(.A1(new_n734), .A2(new_n737), .B1(new_n740), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND3_X1  g540(.A1(new_n715), .A2(new_n627), .A3(new_n651), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT106), .ZN(new_n743));
  OR3_X1    g542(.A1(new_n743), .A2(KEYINPUT107), .A3(new_n708), .ZN(new_n744));
  OAI21_X1  g543(.A(KEYINPUT107), .B1(new_n743), .B2(new_n708), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(new_n476), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(G57gat), .ZN(G1332gat));
  OAI22_X1  g548(.A1(new_n746), .A2(new_n656), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT108), .ZN(new_n751));
  XNOR2_X1  g550(.A(KEYINPUT49), .B(G64gat), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n744), .A2(new_n474), .A3(new_n745), .A4(new_n752), .ZN(new_n753));
  AND3_X1   g552(.A1(new_n750), .A2(new_n751), .A3(new_n753), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n751), .B1(new_n750), .B2(new_n753), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n754), .A2(new_n755), .ZN(G1333gat));
  INV_X1    g555(.A(G71gat), .ZN(new_n757));
  XOR2_X1   g556(.A(new_n480), .B(KEYINPUT109), .Z(new_n758));
  OAI21_X1  g557(.A(new_n757), .B1(new_n746), .B2(new_n758), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n744), .A2(G71gat), .A3(new_n484), .A4(new_n745), .ZN(new_n760));
  XNOR2_X1  g559(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n761));
  AND3_X1   g560(.A1(new_n759), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n761), .B1(new_n759), .B2(new_n760), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n762), .A2(new_n763), .ZN(G1334gat));
  NAND2_X1  g563(.A1(new_n747), .A2(new_n701), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g565(.A1(new_n522), .A2(new_n484), .A3(new_n684), .ZN(new_n767));
  AOI22_X1  g566(.A1(new_n691), .A2(new_n695), .B1(new_n698), .B2(new_n701), .ZN(new_n768));
  AOI21_X1  g567(.A(KEYINPUT102), .B1(new_n768), .B2(new_n664), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n479), .B1(new_n767), .B2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT112), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n770), .A2(new_n771), .A3(new_n626), .ZN(new_n772));
  OAI21_X1  g571(.A(KEYINPUT112), .B1(new_n708), .B2(new_n683), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n715), .A2(new_n604), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT111), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n772), .A2(new_n773), .A3(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n772), .A2(new_n773), .A3(KEYINPUT51), .A4(new_n775), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n778), .A2(KEYINPUT113), .A3(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT113), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n776), .A2(new_n781), .A3(new_n777), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n485), .A2(G85gat), .A3(new_n652), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n780), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n775), .A2(new_n651), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n711), .A2(new_n476), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(G85gat), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n784), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(KEYINPUT114), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT114), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n784), .A2(new_n788), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n790), .A2(new_n792), .ZN(G1336gat));
  NAND3_X1  g592(.A1(new_n711), .A2(new_n474), .A3(new_n786), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(G92gat), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n652), .A2(new_n656), .A3(G92gat), .ZN(new_n798));
  AND3_X1   g597(.A1(new_n780), .A2(new_n782), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n778), .A2(new_n779), .ZN(new_n800));
  AOI22_X1  g599(.A1(new_n794), .A2(G92gat), .B1(new_n800), .B2(new_n798), .ZN(new_n801));
  OAI22_X1  g600(.A1(new_n797), .A2(new_n799), .B1(new_n801), .B2(new_n796), .ZN(G1337gat));
  INV_X1    g601(.A(G99gat), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n480), .A2(new_n803), .A3(new_n651), .ZN(new_n804));
  XOR2_X1   g603(.A(new_n804), .B(KEYINPUT115), .Z(new_n805));
  NAND3_X1  g604(.A1(new_n780), .A2(new_n782), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n705), .A2(new_n680), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n709), .ZN(new_n808));
  INV_X1    g607(.A(new_n710), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n681), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n810), .A2(new_n664), .A3(new_n785), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n806), .B1(new_n811), .B2(new_n803), .ZN(G1338gat));
  INV_X1    g611(.A(KEYINPUT53), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n810), .A2(new_n503), .A3(new_n785), .ZN(new_n814));
  INV_X1    g613(.A(G106gat), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n813), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n652), .A2(new_n503), .A3(G106gat), .ZN(new_n817));
  AND3_X1   g616(.A1(new_n780), .A2(new_n782), .A3(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n711), .A2(new_n701), .A3(new_n786), .ZN(new_n819));
  AOI22_X1  g618(.A1(new_n819), .A2(G106gat), .B1(new_n800), .B2(new_n817), .ZN(new_n820));
  OAI22_X1  g619(.A1(new_n816), .A2(new_n818), .B1(new_n813), .B2(new_n820), .ZN(G1339gat));
  NAND2_X1  g620(.A1(new_n638), .A2(new_n639), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n822), .A2(KEYINPUT54), .A3(new_n649), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n824));
  INV_X1    g623(.A(new_n639), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n824), .B(new_n825), .C1(new_n648), .C2(new_n637), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n823), .A2(KEYINPUT55), .A3(new_n644), .A4(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT116), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n827), .A2(new_n828), .A3(new_n650), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n823), .A2(new_n644), .A3(new_n826), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT55), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n828), .B1(new_n827), .B2(new_n650), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n712), .A2(new_n835), .A3(new_n714), .ZN(new_n836));
  INV_X1    g635(.A(new_n569), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n550), .A2(new_n552), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n838), .A2(KEYINPUT117), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n551), .B1(new_n563), .B2(new_n544), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n838), .A2(KEYINPUT117), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n837), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n579), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n845), .A2(new_n652), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n626), .B1(new_n836), .B2(new_n847), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n835), .A2(new_n626), .A3(new_n579), .A4(new_n844), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n604), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n627), .A2(new_n652), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n716), .A2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n701), .B1(new_n851), .B2(new_n854), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n855), .A2(new_n476), .A3(new_n480), .A4(new_n656), .ZN(new_n856));
  INV_X1    g655(.A(G113gat), .ZN(new_n857));
  INV_X1    g656(.A(new_n581), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n485), .B1(new_n851), .B2(new_n854), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n860), .A2(new_n475), .ZN(new_n861));
  AOI21_X1  g660(.A(G113gat), .B1(new_n861), .B2(new_n716), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n859), .A2(new_n862), .ZN(G1340gat));
  INV_X1    g662(.A(G120gat), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n856), .A2(new_n864), .A3(new_n652), .ZN(new_n865));
  AOI21_X1  g664(.A(G120gat), .B1(new_n861), .B2(new_n651), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n865), .A2(new_n866), .ZN(G1341gat));
  OAI21_X1  g666(.A(G127gat), .B1(new_n856), .B2(new_n604), .ZN(new_n868));
  INV_X1    g667(.A(G127gat), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n861), .A2(new_n869), .A3(new_n672), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n868), .A2(new_n870), .ZN(G1342gat));
  INV_X1    g670(.A(G134gat), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n861), .A2(new_n872), .A3(new_n626), .ZN(new_n873));
  OR2_X1    g672(.A1(new_n873), .A2(KEYINPUT56), .ZN(new_n874));
  OAI21_X1  g673(.A(G134gat), .B1(new_n856), .B2(new_n683), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n873), .A2(KEYINPUT56), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(G1343gat));
  NOR3_X1   g676(.A1(new_n484), .A2(new_n503), .A3(new_n474), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n860), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n858), .A2(G141gat), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT120), .ZN(new_n882));
  AOI21_X1  g681(.A(KEYINPUT58), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n851), .A2(new_n854), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT57), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n884), .A2(new_n885), .A3(new_n286), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n484), .A2(new_n485), .A3(new_n474), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n887), .B(KEYINPUT118), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n832), .A2(new_n650), .A3(new_n827), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n889), .B1(new_n580), .B2(new_n579), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n683), .B1(new_n846), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n672), .B1(new_n891), .B2(new_n849), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n701), .B1(new_n892), .B2(new_n853), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n888), .B1(new_n893), .B2(KEYINPUT57), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n886), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(G141gat), .B1(new_n895), .B2(new_n858), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n883), .B(new_n896), .C1(new_n882), .C2(new_n881), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT119), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n886), .A2(new_n894), .A3(new_n716), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(G141gat), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n881), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n898), .B1(new_n901), .B2(KEYINPUT58), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT58), .ZN(new_n903));
  AOI211_X1 g702(.A(KEYINPUT119), .B(new_n903), .C1(new_n900), .C2(new_n881), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n897), .B1(new_n902), .B2(new_n904), .ZN(G1344gat));
  NAND2_X1  g704(.A1(new_n233), .A2(new_n235), .ZN(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n879), .A2(new_n907), .A3(new_n651), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT121), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n908), .B(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT59), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n884), .A2(new_n286), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(KEYINPUT57), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n852), .A2(new_n581), .ZN(new_n914));
  OAI211_X1 g713(.A(new_n885), .B(new_n701), .C1(new_n892), .C2(new_n914), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n888), .A2(new_n652), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n913), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n911), .B1(new_n917), .B2(G148gat), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n895), .A2(new_n652), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n919), .A2(KEYINPUT59), .A3(new_n907), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n910), .B1(new_n918), .B2(new_n920), .ZN(G1345gat));
  OAI21_X1  g720(.A(G155gat), .B1(new_n895), .B2(new_n604), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n879), .A2(new_n227), .A3(new_n672), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(G1346gat));
  NOR3_X1   g723(.A1(new_n895), .A2(new_n228), .A3(new_n683), .ZN(new_n925));
  AOI21_X1  g724(.A(G162gat), .B1(new_n879), .B2(new_n626), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n925), .A2(new_n926), .ZN(G1347gat));
  NOR2_X1   g726(.A1(new_n476), .A2(new_n656), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n884), .A2(new_n928), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n929), .A2(new_n387), .ZN(new_n930));
  NAND4_X1  g729(.A1(new_n930), .A2(new_n323), .A3(new_n325), .A4(new_n716), .ZN(new_n931));
  XOR2_X1   g730(.A(new_n928), .B(KEYINPUT122), .Z(new_n932));
  NOR2_X1   g731(.A1(new_n932), .A2(new_n758), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n855), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g733(.A(G169gat), .B1(new_n934), .B2(new_n858), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n931), .A2(new_n935), .ZN(G1348gat));
  NAND3_X1  g735(.A1(new_n930), .A2(new_n302), .A3(new_n651), .ZN(new_n937));
  OAI21_X1  g736(.A(G176gat), .B1(new_n934), .B2(new_n652), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(G1349gat));
  INV_X1    g738(.A(KEYINPUT123), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n940), .A2(KEYINPUT60), .ZN(new_n941));
  NAND4_X1  g740(.A1(new_n929), .A2(new_n340), .A3(new_n387), .A4(new_n672), .ZN(new_n942));
  OAI21_X1  g741(.A(G183gat), .B1(new_n934), .B2(new_n604), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n941), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n940), .A2(KEYINPUT60), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n944), .B(new_n945), .ZN(G1350gat));
  NAND4_X1  g745(.A1(new_n929), .A2(new_n317), .A3(new_n387), .A4(new_n626), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n855), .A2(new_n626), .A3(new_n933), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT61), .ZN(new_n949));
  AND4_X1   g748(.A1(KEYINPUT124), .A2(new_n948), .A3(new_n949), .A4(G190gat), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT124), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n317), .B1(new_n951), .B2(KEYINPUT61), .ZN(new_n952));
  AOI22_X1  g751(.A1(new_n948), .A2(new_n952), .B1(KEYINPUT124), .B2(new_n949), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n947), .B1(new_n950), .B2(new_n953), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT125), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI211_X1 g755(.A(KEYINPUT125), .B(new_n947), .C1(new_n950), .C2(new_n953), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(G1351gat));
  AND3_X1   g757(.A1(new_n929), .A2(new_n664), .A3(new_n286), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n959), .A2(new_n248), .A3(new_n716), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n932), .A2(new_n484), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n913), .A2(new_n915), .A3(new_n961), .ZN(new_n962));
  OAI21_X1  g761(.A(KEYINPUT126), .B1(new_n962), .B2(new_n858), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(G197gat), .ZN(new_n964));
  NOR3_X1   g763(.A1(new_n962), .A2(KEYINPUT126), .A3(new_n858), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n960), .B1(new_n964), .B2(new_n965), .ZN(G1352gat));
  NAND3_X1  g765(.A1(new_n959), .A2(new_n249), .A3(new_n651), .ZN(new_n967));
  OR2_X1    g766(.A1(new_n967), .A2(KEYINPUT62), .ZN(new_n968));
  OAI21_X1  g767(.A(G204gat), .B1(new_n962), .B2(new_n652), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n967), .A2(KEYINPUT62), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(G1353gat));
  NAND3_X1  g770(.A1(new_n959), .A2(new_n239), .A3(new_n672), .ZN(new_n972));
  NAND4_X1  g771(.A1(new_n913), .A2(new_n672), .A3(new_n915), .A4(new_n961), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n973), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n974));
  INV_X1    g773(.A(new_n974), .ZN(new_n975));
  AOI21_X1  g774(.A(KEYINPUT63), .B1(new_n973), .B2(G211gat), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n972), .B1(new_n975), .B2(new_n976), .ZN(G1354gat));
  OAI21_X1  g776(.A(G218gat), .B1(new_n962), .B2(new_n683), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n959), .A2(new_n240), .A3(new_n626), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n978), .A2(new_n979), .ZN(G1355gat));
endmodule


