//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 0 0 1 0 1 0 1 1 0 1 0 0 1 0 0 0 0 1 1 1 1 1 1 0 0 1 0 1 0 0 0 1 1 0 1 1 0 1 1 1 0 0 1 0 1 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:09 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n774, new_n775, new_n776, new_n777, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n789, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT32), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT71), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT0), .B(G128), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  AND2_X1   g007(.A1(KEYINPUT64), .A2(G143), .ZN(new_n194));
  NOR2_X1   g008(.A1(KEYINPUT64), .A2(G143), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n193), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n193), .A2(G143), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n192), .B1(new_n196), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT64), .ZN(new_n200));
  INV_X1    g014(.A(G143), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(KEYINPUT64), .A2(G143), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n202), .A2(G146), .A3(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n193), .A2(G143), .ZN(new_n205));
  AND2_X1   g019(.A1(KEYINPUT0), .A2(G128), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n204), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT65), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n204), .A2(KEYINPUT65), .A3(new_n205), .A4(new_n206), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n199), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G137), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n212), .A2(KEYINPUT11), .A3(G134), .ZN(new_n213));
  INV_X1    g027(.A(G134), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G137), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(KEYINPUT68), .B(G131), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT11), .ZN(new_n219));
  OAI211_X1 g033(.A(KEYINPUT67), .B(new_n219), .C1(new_n214), .C2(G137), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n212), .A2(G134), .ZN(new_n222));
  AOI21_X1  g036(.A(KEYINPUT67), .B1(new_n222), .B2(new_n219), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n217), .B(new_n218), .C1(new_n221), .C2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G131), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n219), .B1(new_n214), .B2(G137), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n216), .B1(new_n228), .B2(new_n220), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n224), .B1(new_n225), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n211), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G128), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n232), .A2(KEYINPUT1), .ZN(new_n233));
  AND3_X1   g047(.A1(new_n204), .A2(new_n205), .A3(new_n233), .ZN(new_n234));
  OAI21_X1  g048(.A(KEYINPUT1), .B1(new_n201), .B2(G146), .ZN(new_n235));
  AOI22_X1  g049(.A1(new_n196), .A2(new_n198), .B1(G128), .B2(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(KEYINPUT70), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n225), .B1(new_n222), .B2(new_n215), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n238), .B1(new_n229), .B2(new_n218), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n204), .A2(new_n205), .A3(new_n233), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT70), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n202), .A2(new_n203), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n197), .B1(new_n242), .B2(new_n193), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n235), .A2(G128), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n240), .B(new_n241), .C1(new_n243), .C2(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n237), .A2(new_n239), .A3(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n231), .A2(new_n247), .A3(KEYINPUT30), .ZN(new_n248));
  XOR2_X1   g062(.A(KEYINPUT2), .B(G113), .Z(new_n249));
  XNOR2_X1  g063(.A(G116), .B(G119), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT2), .B(G113), .ZN(new_n252));
  INV_X1    g066(.A(G116), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n253), .A2(G119), .ZN(new_n254));
  INV_X1    g068(.A(G119), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n255), .A2(G116), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n252), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  AND3_X1   g071(.A1(new_n251), .A2(new_n257), .A3(KEYINPUT69), .ZN(new_n258));
  AOI21_X1  g072(.A(KEYINPUT69), .B1(new_n251), .B2(new_n257), .ZN(new_n259));
  OR2_X1    g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n248), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT30), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n239), .B1(new_n236), .B2(new_n234), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n230), .B1(new_n211), .B2(KEYINPUT66), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT66), .ZN(new_n265));
  AOI211_X1 g079(.A(new_n265), .B(new_n199), .C1(new_n209), .C2(new_n210), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n263), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n261), .B1(new_n262), .B2(new_n267), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n258), .A2(new_n259), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n231), .A2(new_n247), .A3(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G237), .ZN(new_n271));
  INV_X1    g085(.A(G953), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n271), .A2(new_n272), .A3(G210), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n273), .B(KEYINPUT27), .ZN(new_n274));
  XNOR2_X1  g088(.A(KEYINPUT26), .B(G101), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n274), .B(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n270), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n191), .B1(new_n268), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n267), .A2(new_n262), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n248), .A2(new_n260), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n277), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n281), .A2(KEYINPUT71), .A3(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n278), .A2(KEYINPUT31), .A3(new_n283), .ZN(new_n284));
  AND3_X1   g098(.A1(new_n231), .A2(new_n247), .A3(new_n269), .ZN(new_n285));
  OR2_X1    g099(.A1(new_n285), .A2(KEYINPUT28), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n285), .B1(new_n267), .B2(new_n260), .ZN(new_n287));
  XNOR2_X1  g101(.A(KEYINPUT73), .B(KEYINPUT28), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  XNOR2_X1  g103(.A(new_n276), .B(KEYINPUT72), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n277), .B1(new_n279), .B2(new_n280), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT31), .ZN(new_n292));
  AOI22_X1  g106(.A1(new_n289), .A2(new_n290), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  AND3_X1   g107(.A1(new_n284), .A2(new_n293), .A3(KEYINPUT74), .ZN(new_n294));
  AOI21_X1  g108(.A(KEYINPUT74), .B1(new_n284), .B2(new_n293), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n190), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n269), .B1(new_n231), .B2(new_n247), .ZN(new_n297));
  OR2_X1    g111(.A1(new_n285), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(KEYINPUT28), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(new_n286), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n276), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT29), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(G902), .B1(new_n301), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n281), .A2(new_n270), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(new_n302), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n307), .B(new_n303), .C1(new_n289), .C2(new_n290), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G472), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n284), .A2(new_n293), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT74), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n284), .A2(new_n293), .A3(KEYINPUT74), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n188), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n296), .B(new_n310), .C1(new_n315), .C2(KEYINPUT32), .ZN(new_n316));
  INV_X1    g130(.A(G217), .ZN(new_n317));
  INV_X1    g131(.A(G902), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n317), .B1(G234), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT16), .ZN(new_n321));
  INV_X1    g135(.A(G140), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n321), .A2(new_n322), .A3(G125), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(G125), .ZN(new_n324));
  INV_X1    g138(.A(G125), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G140), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n323), .B1(new_n327), .B2(new_n321), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n193), .ZN(new_n329));
  OAI211_X1 g143(.A(G146), .B(new_n323), .C1(new_n327), .C2(new_n321), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n255), .A2(G128), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n232), .A2(KEYINPUT23), .A3(G119), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n232), .A2(G119), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  OAI211_X1 g148(.A(new_n331), .B(new_n332), .C1(new_n334), .C2(KEYINPUT23), .ZN(new_n335));
  AOI22_X1  g149(.A1(new_n329), .A2(new_n330), .B1(G110), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n333), .A2(new_n331), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT75), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n333), .A2(new_n331), .A3(KEYINPUT75), .ZN(new_n340));
  XOR2_X1   g154(.A(KEYINPUT24), .B(G110), .Z(new_n341));
  NAND3_X1  g155(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT76), .ZN(new_n343));
  AND2_X1   g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n342), .A2(new_n343), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n336), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  AND2_X1   g160(.A1(new_n339), .A2(new_n340), .ZN(new_n347));
  OAI22_X1  g161(.A1(new_n347), .A2(new_n341), .B1(G110), .B2(new_n335), .ZN(new_n348));
  XNOR2_X1  g162(.A(G125), .B(G140), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n193), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n348), .A2(new_n330), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n346), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(KEYINPUT22), .B(G137), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n272), .A2(G221), .A3(G234), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n353), .B(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n352), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n346), .A2(new_n351), .A3(new_n355), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(new_n318), .A3(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT25), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n357), .A2(KEYINPUT25), .A3(new_n318), .A4(new_n358), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n320), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n358), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n355), .B1(new_n346), .B2(new_n351), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  XOR2_X1   g180(.A(new_n366), .B(KEYINPUT77), .Z(new_n367));
  NOR2_X1   g181(.A1(new_n319), .A2(G902), .ZN(new_n368));
  XOR2_X1   g182(.A(new_n368), .B(KEYINPUT78), .Z(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n363), .B1(new_n367), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(G214), .B1(G237), .B2(G902), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n372), .B(KEYINPUT81), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT80), .ZN(new_n375));
  XNOR2_X1  g189(.A(G104), .B(G107), .ZN(new_n376));
  INV_X1    g190(.A(G101), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n375), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G107), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G104), .ZN(new_n380));
  INV_X1    g194(.A(G104), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G107), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n383), .A2(KEYINPUT80), .A3(G101), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n378), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT3), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n386), .B(new_n382), .C1(new_n380), .C2(KEYINPUT79), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT79), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n388), .A2(new_n379), .A3(KEYINPUT3), .A4(G104), .ZN(new_n389));
  AOI21_X1  g203(.A(G101), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n385), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n250), .A2(KEYINPUT5), .ZN(new_n392));
  INV_X1    g206(.A(G113), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT5), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n393), .B1(new_n254), .B2(new_n394), .ZN(new_n395));
  AOI22_X1  g209(.A1(new_n392), .A2(new_n395), .B1(new_n249), .B2(new_n250), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n391), .A2(new_n396), .ZN(new_n397));
  XNOR2_X1  g211(.A(G110), .B(G122), .ZN(new_n398));
  NOR3_X1   g212(.A1(new_n381), .A2(KEYINPUT79), .A3(G107), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n386), .B1(new_n379), .B2(G104), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n389), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n377), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n387), .A2(G101), .A3(new_n389), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(KEYINPUT4), .A3(new_n403), .ZN(new_n404));
  OR3_X1    g218(.A1(new_n401), .A2(KEYINPUT4), .A3(new_n377), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n397), .B(new_n398), .C1(new_n269), .C2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT85), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n407), .B(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n392), .A2(KEYINPUT87), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n395), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n392), .A2(KEYINPUT87), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n251), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n391), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT88), .ZN(new_n415));
  XOR2_X1   g229(.A(new_n398), .B(KEYINPUT8), .Z(new_n416));
  NAND3_X1  g230(.A1(new_n402), .A2(new_n384), .A3(new_n378), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n416), .B1(new_n417), .B2(new_n396), .ZN(new_n418));
  AND3_X1   g232(.A1(new_n414), .A2(new_n415), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n415), .B1(new_n414), .B2(new_n418), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT7), .ZN(new_n421));
  INV_X1    g235(.A(new_n236), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n422), .A2(new_n325), .A3(new_n240), .ZN(new_n423));
  XNOR2_X1  g237(.A(KEYINPUT86), .B(G224), .ZN(new_n424));
  OAI221_X1 g238(.A(new_n423), .B1(G953), .B2(new_n424), .C1(new_n211), .C2(new_n325), .ZN(new_n425));
  OAI22_X1  g239(.A1(new_n419), .A2(new_n420), .B1(new_n421), .B2(new_n425), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n409), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n423), .B1(new_n211), .B2(new_n325), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n424), .A2(G953), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n428), .B1(new_n421), .B2(new_n429), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n430), .B(KEYINPUT89), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(G902), .B1(new_n427), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n397), .B1(new_n269), .B2(new_n406), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT82), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n397), .B(KEYINPUT82), .C1(new_n269), .C2(new_n406), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n398), .B(KEYINPUT83), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n436), .A2(new_n437), .A3(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT84), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT6), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n260), .A2(new_n405), .A3(new_n404), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n444), .A2(new_n397), .A3(new_n408), .A4(new_n398), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n407), .A2(KEYINPUT85), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n445), .A2(KEYINPUT6), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n438), .B1(new_n434), .B2(new_n435), .ZN(new_n448));
  INV_X1    g262(.A(new_n442), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n448), .A2(new_n449), .A3(new_n437), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n443), .A2(new_n447), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n428), .A2(new_n429), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(new_n425), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(G210), .B1(G237), .B2(G902), .ZN(new_n455));
  AND3_X1   g269(.A1(new_n433), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n455), .B1(new_n433), .B2(new_n454), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n374), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(KEYINPUT9), .B(G234), .ZN(new_n459));
  NOR3_X1   g273(.A1(new_n459), .A2(new_n317), .A3(G953), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(KEYINPUT94), .B1(new_n242), .B2(new_n232), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n194), .A2(new_n195), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT94), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n463), .A2(new_n464), .A3(G128), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n201), .A2(G128), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n214), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  AOI211_X1 g283(.A(G134), .B(new_n467), .C1(new_n462), .C2(new_n465), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(G122), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(G116), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n253), .A2(G122), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n473), .A2(new_n474), .A3(KEYINPUT93), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(KEYINPUT93), .B1(new_n473), .B2(new_n474), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n379), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n474), .A2(KEYINPUT14), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT14), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n480), .A2(new_n253), .A3(G122), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n479), .A2(new_n481), .A3(KEYINPUT95), .A4(new_n473), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT96), .ZN(new_n483));
  NOR3_X1   g297(.A1(new_n472), .A2(KEYINPUT14), .A3(G116), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT95), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n379), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n482), .A2(new_n483), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n483), .B1(new_n482), .B2(new_n486), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n478), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n471), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT93), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n253), .A2(G122), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n472), .A2(G116), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n495), .A2(G107), .A3(new_n475), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n478), .A2(new_n496), .ZN(new_n497));
  NOR3_X1   g311(.A1(new_n242), .A2(KEYINPUT94), .A3(new_n232), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n464), .B1(new_n463), .B2(G128), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n214), .B(new_n468), .C1(new_n498), .C2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT13), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n466), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n462), .A2(KEYINPUT13), .A3(new_n465), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n503), .A2(new_n504), .A3(new_n468), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n501), .B1(new_n505), .B2(G134), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n461), .B1(new_n491), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n489), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n487), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n509), .B(new_n478), .C1(new_n470), .C2(new_n469), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n467), .B1(new_n466), .B2(new_n502), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n214), .B1(new_n511), .B2(new_n504), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n510), .B(new_n460), .C1(new_n512), .C2(new_n501), .ZN(new_n513));
  AOI21_X1  g327(.A(G902), .B1(new_n507), .B2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(G478), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n515), .A2(KEYINPUT15), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n514), .B(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(G234), .A2(G237), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n519), .A2(G952), .A3(new_n272), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n520), .B(KEYINPUT97), .ZN(new_n521));
  AND3_X1   g335(.A1(new_n519), .A2(G902), .A3(G953), .ZN(new_n522));
  XNOR2_X1  g336(.A(KEYINPUT21), .B(G898), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AND2_X1   g338(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n271), .A2(new_n272), .A3(G214), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n463), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n271), .A2(new_n272), .A3(G143), .A4(G214), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n218), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT17), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n527), .A2(new_n218), .A3(new_n528), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  AND2_X1   g348(.A1(new_n329), .A2(new_n330), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n529), .A2(KEYINPUT17), .A3(new_n530), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(KEYINPUT18), .A2(G131), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n538), .B1(new_n527), .B2(new_n528), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT90), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n327), .A2(G146), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n349), .A2(new_n193), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n327), .A2(G146), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n544), .A2(new_n350), .A3(KEYINPUT90), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n539), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n527), .A2(new_n538), .A3(new_n528), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT91), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n527), .A2(KEYINPUT91), .A3(new_n538), .A4(new_n528), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n546), .A2(new_n551), .ZN(new_n552));
  XNOR2_X1  g366(.A(G113), .B(G122), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n553), .B(new_n381), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT92), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n554), .B(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n537), .A2(new_n552), .A3(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n554), .B1(new_n537), .B2(new_n552), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n318), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(G475), .ZN(new_n561));
  INV_X1    g375(.A(new_n330), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n349), .B(KEYINPUT19), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n562), .B1(new_n193), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n531), .A2(new_n533), .ZN(new_n565));
  AOI22_X1  g379(.A1(new_n551), .A2(new_n546), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n557), .B1(new_n566), .B2(new_n554), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT20), .ZN(new_n568));
  NOR2_X1   g382(.A1(G475), .A2(G902), .ZN(new_n569));
  AND3_X1   g383(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n568), .B1(new_n567), .B2(new_n569), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n561), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NOR3_X1   g386(.A1(new_n518), .A2(new_n525), .A3(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(G221), .B1(new_n459), .B2(G902), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  AND2_X1   g389(.A1(new_n204), .A2(new_n205), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n232), .B1(new_n196), .B2(KEYINPUT1), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n240), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n391), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT10), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n230), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n237), .A2(new_n391), .A3(KEYINPUT10), .A4(new_n246), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n211), .A2(new_n405), .A3(new_n404), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n581), .A2(new_n582), .A3(new_n583), .A4(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n417), .A2(new_n422), .A3(new_n240), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n579), .A2(new_n586), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n587), .A2(KEYINPUT12), .A3(new_n230), .ZN(new_n588));
  AOI21_X1  g402(.A(KEYINPUT12), .B1(new_n587), .B2(new_n230), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n585), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(G110), .B(G140), .ZN(new_n591));
  INV_X1    g405(.A(G227), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n592), .A2(G953), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n591), .B(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  AND2_X1   g409(.A1(new_n585), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n581), .A2(new_n583), .A3(new_n584), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n230), .ZN(new_n598));
  AOI22_X1  g412(.A1(new_n590), .A2(new_n594), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(G469), .B1(new_n599), .B2(G902), .ZN(new_n600));
  INV_X1    g414(.A(G469), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n588), .A2(new_n589), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n585), .A2(new_n595), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n595), .B1(new_n598), .B2(new_n585), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n601), .B(new_n318), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n575), .B1(new_n600), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n573), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n458), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n316), .A2(new_n371), .A3(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(KEYINPUT98), .B(G101), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(G3));
  OAI21_X1  g426(.A(new_n318), .B1(new_n294), .B2(new_n295), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(G472), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n187), .B1(new_n294), .B2(new_n295), .ZN(new_n615));
  INV_X1    g429(.A(new_n607), .ZN(new_n616));
  INV_X1    g430(.A(new_n371), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n614), .A2(new_n615), .A3(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT101), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n515), .A2(G902), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT33), .ZN(new_n622));
  AND3_X1   g436(.A1(new_n507), .A2(new_n622), .A3(new_n513), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n622), .B1(new_n507), .B2(new_n513), .ZN(new_n624));
  OAI211_X1 g438(.A(KEYINPUT99), .B(new_n621), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n621), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n507), .A2(new_n513), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(KEYINPUT33), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n507), .A2(new_n513), .A3(new_n622), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n626), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT99), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n631), .B1(new_n514), .B2(G478), .ZN(new_n632));
  OAI211_X1 g446(.A(new_n625), .B(new_n572), .C1(new_n630), .C2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(KEYINPUT100), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n627), .A2(new_n318), .ZN(new_n635));
  AOI21_X1  g449(.A(KEYINPUT99), .B1(new_n635), .B2(new_n515), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n621), .B1(new_n623), .B2(new_n624), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT100), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n638), .A2(new_n639), .A3(new_n572), .A4(new_n625), .ZN(new_n640));
  AND2_X1   g454(.A1(new_n634), .A2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n525), .ZN(new_n642));
  OAI211_X1 g456(.A(new_n374), .B(new_n642), .C1(new_n456), .C2(new_n457), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n620), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n634), .A2(new_n640), .ZN(new_n645));
  INV_X1    g459(.A(new_n455), .ZN(new_n646));
  INV_X1    g460(.A(new_n453), .ZN(new_n647));
  AND3_X1   g461(.A1(new_n448), .A2(new_n449), .A3(new_n437), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n449), .B1(new_n448), .B2(new_n437), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n647), .B1(new_n650), .B2(new_n447), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n445), .A2(new_n446), .ZN(new_n652));
  OR2_X1    g466(.A1(new_n425), .A2(new_n421), .ZN(new_n653));
  OAI211_X1 g467(.A(new_n652), .B(new_n653), .C1(new_n419), .C2(new_n420), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n318), .B1(new_n654), .B2(new_n431), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n646), .B1(new_n651), .B2(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n433), .A2(new_n454), .A3(new_n455), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n373), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n645), .A2(new_n658), .A3(KEYINPUT101), .A4(new_n642), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n619), .B1(new_n644), .B2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT34), .B(G104), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G6));
  INV_X1    g476(.A(KEYINPUT103), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n567), .A2(new_n569), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(KEYINPUT20), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n561), .A2(KEYINPUT102), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT102), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n560), .A2(new_n669), .A3(G475), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n667), .A2(new_n668), .A3(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n514), .A2(new_n517), .ZN(new_n672));
  AOI211_X1 g486(.A(G902), .B(new_n516), .C1(new_n507), .C2(new_n513), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n663), .B1(new_n643), .B2(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n658), .A2(KEYINPUT103), .A3(new_n642), .A4(new_n675), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n619), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(KEYINPUT35), .B(G107), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G9));
  NAND2_X1  g495(.A1(new_n361), .A2(new_n362), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n319), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT104), .ZN(new_n684));
  OR2_X1    g498(.A1(new_n356), .A2(KEYINPUT36), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n352), .B(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n686), .A2(new_n369), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n683), .A2(new_n684), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g503(.A(KEYINPUT104), .B1(new_n363), .B2(new_n687), .ZN(new_n690));
  AND2_X1   g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n609), .A2(new_n614), .A3(new_n615), .A4(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(KEYINPUT37), .B(G110), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(KEYINPUT105), .ZN(new_n694));
  XOR2_X1   g508(.A(new_n694), .B(KEYINPUT106), .Z(new_n695));
  XNOR2_X1  g509(.A(new_n692), .B(new_n695), .ZN(G12));
  NAND2_X1  g510(.A1(new_n600), .A2(new_n606), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n697), .A2(new_n689), .A3(new_n574), .A4(new_n690), .ZN(new_n698));
  INV_X1    g512(.A(G900), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n522), .A2(new_n699), .ZN(new_n700));
  AND2_X1   g514(.A1(new_n521), .A2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n675), .A2(new_n702), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n458), .A2(new_n698), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n316), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G128), .ZN(G30));
  NAND2_X1  g520(.A1(new_n313), .A2(new_n314), .ZN(new_n707));
  AND2_X1   g521(.A1(new_n278), .A2(new_n283), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n298), .A2(new_n290), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n318), .ZN(new_n711));
  AOI22_X1  g525(.A1(new_n707), .A2(new_n190), .B1(G472), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n615), .A2(new_n189), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n656), .A2(new_n657), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(KEYINPUT38), .ZN(new_n716));
  XOR2_X1   g530(.A(new_n701), .B(KEYINPUT39), .Z(new_n717));
  NAND2_X1  g531(.A1(new_n607), .A2(new_n717), .ZN(new_n718));
  OR2_X1    g532(.A1(new_n718), .A2(KEYINPUT40), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n363), .A2(new_n687), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n720), .A2(new_n374), .A3(new_n518), .A4(new_n572), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n721), .B1(new_n718), .B2(KEYINPUT40), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n714), .A2(new_n716), .A3(new_n719), .A4(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n242), .B(KEYINPUT107), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n723), .B(new_n724), .ZN(G45));
  NAND4_X1  g539(.A1(new_n638), .A2(new_n572), .A3(new_n625), .A4(new_n702), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n458), .A2(new_n698), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n316), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(KEYINPUT108), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT108), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n316), .A2(new_n730), .A3(new_n727), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G146), .ZN(G48));
  NAND2_X1  g547(.A1(new_n644), .A2(new_n659), .ZN(new_n734));
  AND2_X1   g548(.A1(new_n296), .A2(new_n310), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n617), .B1(new_n735), .B2(new_n713), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n318), .B1(new_n604), .B2(new_n605), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(G469), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n738), .A2(new_n574), .A3(new_n606), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT109), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n738), .A2(KEYINPUT109), .A3(new_n574), .A4(new_n606), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n734), .A2(new_n736), .A3(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(KEYINPUT41), .B(G113), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(KEYINPUT110), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n745), .B(new_n747), .ZN(G15));
  NAND2_X1  g562(.A1(new_n677), .A2(new_n678), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n736), .A2(new_n749), .A3(new_n744), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G116), .ZN(G18));
  NAND2_X1  g565(.A1(new_n691), .A2(new_n573), .ZN(new_n752));
  NOR3_X1   g566(.A1(new_n743), .A2(new_n752), .A3(new_n458), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n316), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G119), .ZN(G21));
  NAND3_X1  g569(.A1(new_n741), .A2(new_n642), .A3(new_n742), .ZN(new_n756));
  INV_X1    g570(.A(new_n572), .ZN(new_n757));
  OAI21_X1  g571(.A(KEYINPUT111), .B1(new_n757), .B2(new_n674), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT111), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n572), .B(new_n759), .C1(new_n672), .C2(new_n673), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g575(.A(KEYINPUT112), .B1(new_n458), .B2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(new_n760), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n759), .B1(new_n518), .B2(new_n572), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT112), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n658), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n756), .B1(new_n762), .B2(new_n767), .ZN(new_n768));
  AOI22_X1  g582(.A1(new_n300), .A2(new_n290), .B1(new_n292), .B2(new_n291), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n188), .B1(new_n769), .B2(new_n284), .ZN(new_n770));
  AOI211_X1 g584(.A(new_n617), .B(new_n770), .C1(new_n613), .C2(G472), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n768), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G122), .ZN(G24));
  AOI211_X1 g587(.A(new_n720), .B(new_n770), .C1(new_n613), .C2(G472), .ZN(new_n774));
  INV_X1    g588(.A(new_n726), .ZN(new_n775));
  AND4_X1   g589(.A1(new_n658), .A2(new_n775), .A3(new_n741), .A4(new_n742), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G125), .ZN(G27));
  NAND4_X1  g592(.A1(new_n607), .A2(new_n656), .A3(new_n374), .A4(new_n657), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n779), .A2(new_n726), .ZN(new_n780));
  AOI21_X1  g594(.A(KEYINPUT32), .B1(new_n707), .B2(new_n187), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n296), .A2(new_n310), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n780), .B(new_n371), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT42), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n316), .A2(KEYINPUT42), .A3(new_n371), .A4(new_n780), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G131), .ZN(G33));
  NOR2_X1   g602(.A1(new_n779), .A2(new_n703), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n316), .A2(new_n371), .A3(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G134), .ZN(G36));
  NAND3_X1  g605(.A1(new_n638), .A2(new_n757), .A3(new_n625), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(KEYINPUT43), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(new_n720), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n614), .A2(new_n615), .ZN(new_n795));
  AOI21_X1  g609(.A(KEYINPUT44), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(G469), .A2(G902), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n599), .A2(KEYINPUT45), .ZN(new_n798));
  OAI21_X1  g612(.A(G469), .B1(new_n599), .B2(KEYINPUT45), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n797), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT46), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(new_n606), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n800), .A2(new_n801), .ZN(new_n804));
  OR2_X1    g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n805), .A2(new_n574), .A3(new_n717), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n656), .A2(new_n374), .A3(new_n657), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n796), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n794), .A2(KEYINPUT44), .A3(new_n795), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n809), .A2(KEYINPUT113), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n809), .A2(KEYINPUT113), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n808), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(G137), .ZN(G39));
  NAND3_X1  g627(.A1(new_n805), .A2(KEYINPUT47), .A3(new_n574), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n574), .B1(new_n803), .B2(new_n804), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT47), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  NOR4_X1   g632(.A1(new_n316), .A2(new_n371), .A3(new_n726), .A4(new_n807), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(new_n322), .ZN(G42));
  AND2_X1   g635(.A1(new_n712), .A2(new_n713), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT38), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n715), .B(new_n823), .ZN(new_n824));
  NOR4_X1   g638(.A1(new_n617), .A2(new_n792), .A3(new_n373), .A4(new_n575), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n738), .A2(new_n606), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(KEYINPUT49), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n822), .A2(new_n824), .A3(new_n825), .A4(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT116), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n829), .A2(KEYINPUT50), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n793), .A2(new_n521), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(new_n771), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n824), .A2(new_n373), .A3(new_n744), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n829), .B(KEYINPUT50), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n831), .A2(new_n771), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n829), .A2(KEYINPUT50), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n716), .A2(new_n374), .A3(new_n743), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n830), .B1(new_n834), .B2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  NOR4_X1   g654(.A1(new_n743), .A2(new_n807), .A3(new_n617), .A4(new_n521), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n572), .B1(new_n638), .B2(new_n625), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n822), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT117), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n843), .B(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n807), .ZN(new_n846));
  AND4_X1   g660(.A1(new_n744), .A2(new_n831), .A3(new_n774), .A4(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n826), .A2(new_n575), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n814), .A2(new_n817), .A3(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n832), .A2(new_n807), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n847), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n840), .A2(KEYINPUT51), .A3(new_n845), .A4(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n736), .A2(new_n744), .A3(new_n846), .A4(new_n831), .ZN(new_n853));
  XOR2_X1   g667(.A(new_n853), .B(KEYINPUT48), .Z(new_n854));
  NOR3_X1   g668(.A1(new_n832), .A2(new_n458), .A3(new_n743), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n822), .A2(new_n841), .A3(new_n645), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n272), .A2(G952), .ZN(new_n857));
  XOR2_X1   g671(.A(new_n857), .B(KEYINPUT119), .Z(new_n858));
  NOR4_X1   g672(.A1(new_n854), .A2(new_n855), .A3(new_n856), .A4(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT118), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n840), .A2(new_n845), .A3(new_n851), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT51), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n845), .A2(new_n851), .ZN(new_n864));
  OAI211_X1 g678(.A(new_n860), .B(new_n862), .C1(new_n864), .C2(new_n839), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n852), .B(new_n859), .C1(new_n863), .C2(new_n866), .ZN(new_n867));
  AOI22_X1  g681(.A1(new_n774), .A2(new_n776), .B1(new_n316), .B2(new_n704), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n762), .A2(new_n767), .ZN(new_n869));
  INV_X1    g683(.A(new_n720), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n616), .A2(new_n870), .A3(new_n701), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n869), .A2(new_n714), .A3(new_n871), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n316), .A2(new_n730), .A3(new_n727), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n730), .B1(new_n316), .B2(new_n727), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n868), .B(new_n872), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(KEYINPUT52), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT52), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n732), .A2(new_n877), .A3(new_n868), .A4(new_n872), .ZN(new_n878));
  AND2_X1   g692(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n643), .A2(new_n633), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n880), .A2(new_n615), .A3(new_n614), .A4(new_n618), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n610), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(KEYINPUT114), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT114), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n610), .A2(new_n884), .A3(new_n881), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n757), .A2(new_n518), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n643), .A2(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n887), .A2(new_n615), .A3(new_n614), .A4(new_n618), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(new_n692), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n883), .A2(new_n885), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n770), .B1(new_n613), .B2(G472), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n892), .A2(new_n780), .A3(new_n870), .ZN(new_n893));
  OR3_X1    g707(.A1(new_n671), .A2(new_n518), .A3(new_n701), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n807), .A2(new_n698), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n316), .A2(new_n895), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n790), .A2(new_n893), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n787), .A2(new_n897), .ZN(new_n898));
  AOI22_X1  g712(.A1(new_n768), .A2(new_n771), .B1(new_n753), .B2(new_n316), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n899), .A2(new_n745), .A3(new_n750), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n891), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(KEYINPUT53), .B1(new_n879), .B2(new_n901), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n899), .A2(new_n745), .A3(new_n750), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n790), .A2(new_n893), .A3(new_n896), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n904), .B1(new_n785), .B2(new_n786), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n889), .B1(new_n882), .B2(KEYINPUT114), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n903), .A2(new_n905), .A3(new_n885), .A4(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n876), .A2(new_n878), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n777), .A2(new_n705), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(KEYINPUT52), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n911), .A2(KEYINPUT53), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n907), .A2(new_n908), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g727(.A(KEYINPUT54), .B1(new_n902), .B2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT53), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n911), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n879), .A2(new_n901), .A3(new_n916), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n915), .B1(new_n907), .B2(new_n908), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT54), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n914), .A2(KEYINPUT115), .A3(new_n920), .ZN(new_n921));
  AND3_X1   g735(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT115), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n867), .B1(new_n921), .B2(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(G952), .A2(G953), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n828), .B1(new_n925), .B2(new_n926), .ZN(G75));
  AOI21_X1  g741(.A(new_n318), .B1(new_n917), .B2(new_n918), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(G210), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT56), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n451), .B(new_n647), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT55), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n929), .A2(new_n930), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n932), .B1(new_n929), .B2(new_n930), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n272), .A2(G952), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(G51));
  XOR2_X1   g750(.A(new_n797), .B(KEYINPUT57), .Z(new_n937));
  AOI21_X1  g751(.A(new_n919), .B1(new_n917), .B2(new_n918), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n937), .B1(new_n922), .B2(new_n938), .ZN(new_n939));
  OR2_X1    g753(.A1(new_n604), .A2(new_n605), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n798), .A2(new_n799), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n928), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n935), .B1(new_n941), .B2(new_n943), .ZN(G54));
  INV_X1    g758(.A(KEYINPUT120), .ZN(new_n945));
  AND2_X1   g759(.A1(KEYINPUT58), .A2(G475), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n928), .A2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n567), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n945), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n935), .B1(new_n947), .B2(new_n948), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n928), .A2(KEYINPUT120), .A3(new_n567), .A4(new_n946), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(G60));
  NOR2_X1   g766(.A1(new_n623), .A2(new_n624), .ZN(new_n953));
  NAND2_X1  g767(.A1(G478), .A2(G902), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT59), .Z(new_n955));
  NOR2_X1   g769(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n956), .B1(new_n922), .B2(new_n938), .ZN(new_n957));
  INV_X1    g771(.A(new_n935), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(new_n955), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n921), .A2(new_n924), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n959), .B1(new_n953), .B2(new_n961), .ZN(G63));
  INV_X1    g776(.A(KEYINPUT61), .ZN(new_n963));
  NAND2_X1  g777(.A1(G217), .A2(G902), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT60), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n965), .B1(new_n917), .B2(new_n918), .ZN(new_n966));
  INV_X1    g780(.A(new_n686), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n958), .B1(new_n966), .B2(new_n367), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n963), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n917), .A2(new_n918), .ZN(new_n972));
  INV_X1    g786(.A(new_n965), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(new_n367), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n935), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n976), .A2(KEYINPUT61), .A3(new_n968), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n971), .A2(new_n977), .ZN(G66));
  NAND3_X1  g792(.A1(new_n903), .A2(new_n885), .A3(new_n906), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(new_n272), .ZN(new_n980));
  OAI21_X1  g794(.A(G953), .B1(new_n424), .B2(new_n523), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n980), .A2(KEYINPUT121), .A3(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n982), .B1(KEYINPUT121), .B2(new_n980), .ZN(new_n983));
  OAI211_X1 g797(.A(new_n650), .B(new_n447), .C1(G898), .C2(new_n272), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT122), .Z(new_n985));
  XNOR2_X1  g799(.A(new_n983), .B(new_n985), .ZN(G69));
  OAI21_X1  g800(.A(G953), .B1(new_n592), .B2(new_n699), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(KEYINPUT126), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n279), .A2(new_n248), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n563), .B(KEYINPUT123), .Z(new_n990));
  XOR2_X1   g804(.A(new_n989), .B(new_n990), .Z(new_n991));
  NAND2_X1  g805(.A1(new_n633), .A2(new_n886), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n992), .B(KEYINPUT124), .ZN(new_n993));
  NOR3_X1   g807(.A1(new_n993), .A2(new_n718), .A3(new_n807), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(new_n736), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n812), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n820), .B1(new_n996), .B2(KEYINPUT125), .ZN(new_n997));
  INV_X1    g811(.A(new_n995), .ZN(new_n998));
  OR2_X1    g812(.A1(new_n810), .A2(new_n811), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n998), .B1(new_n999), .B2(new_n808), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT125), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n909), .B1(new_n731), .B2(new_n729), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1003), .A2(new_n723), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT62), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n1003), .A2(KEYINPUT62), .A3(new_n723), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n997), .A2(new_n1002), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n991), .B1(new_n1009), .B2(new_n272), .ZN(new_n1010));
  INV_X1    g824(.A(new_n869), .ZN(new_n1011));
  OAI22_X1  g825(.A1(new_n806), .A2(new_n1011), .B1(new_n703), .B2(new_n779), .ZN(new_n1012));
  AOI22_X1  g826(.A1(new_n1012), .A2(new_n736), .B1(new_n818), .B2(new_n819), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n812), .A2(new_n1013), .A3(new_n787), .A4(new_n1003), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1014), .A2(new_n272), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n699), .A2(G953), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  AND2_X1   g831(.A1(new_n1017), .A2(new_n991), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n988), .B1(new_n1010), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g833(.A(new_n988), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1017), .A2(new_n991), .ZN(new_n1021));
  AOI22_X1  g835(.A1(new_n1000), .A2(new_n1001), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1022));
  AOI21_X1  g836(.A(G953), .B1(new_n1022), .B2(new_n997), .ZN(new_n1023));
  OAI211_X1 g837(.A(new_n1020), .B(new_n1021), .C1(new_n1023), .C2(new_n991), .ZN(new_n1024));
  AND2_X1   g838(.A1(new_n1019), .A2(new_n1024), .ZN(G72));
  NAND2_X1  g839(.A1(G472), .A2(G902), .ZN(new_n1026));
  XOR2_X1   g840(.A(new_n1026), .B(KEYINPUT63), .Z(new_n1027));
  OAI21_X1  g841(.A(new_n1027), .B1(new_n1014), .B2(new_n979), .ZN(new_n1028));
  NOR2_X1   g842(.A1(new_n306), .A2(new_n276), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n935), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n708), .A2(new_n307), .ZN(new_n1031));
  OAI211_X1 g845(.A(new_n1027), .B(new_n1031), .C1(new_n902), .C2(new_n913), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n306), .A2(new_n276), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n1027), .B1(new_n1009), .B2(new_n979), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1034), .B1(new_n1035), .B2(KEYINPUT127), .ZN(new_n1036));
  INV_X1    g850(.A(KEYINPUT127), .ZN(new_n1037));
  OAI211_X1 g851(.A(new_n1037), .B(new_n1027), .C1(new_n1009), .C2(new_n979), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n1033), .B1(new_n1036), .B2(new_n1038), .ZN(G57));
endmodule


