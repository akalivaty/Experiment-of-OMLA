//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 0 1 1 0 0 0 0 0 1 1 1 1 1 1 1 1 1 0 1 1 0 0 1 0 0 0 0 0 1 0 0 0 0 1 1 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:25 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT25), .ZN(new_n191));
  INV_X1    g005(.A(G110), .ZN(new_n192));
  INV_X1    g006(.A(G128), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n193), .A2(KEYINPUT23), .A3(G119), .ZN(new_n194));
  AND2_X1   g008(.A1(KEYINPUT68), .A2(G119), .ZN(new_n195));
  NOR2_X1   g009(.A1(KEYINPUT68), .A2(G119), .ZN(new_n196));
  OAI211_X1 g010(.A(KEYINPUT71), .B(new_n193), .C1(new_n195), .C2(new_n196), .ZN(new_n197));
  NOR3_X1   g011(.A1(new_n195), .A2(new_n196), .A3(new_n193), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT23), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n197), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT68), .ZN(new_n201));
  INV_X1    g015(.A(G119), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(KEYINPUT68), .A2(G119), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  AOI21_X1  g019(.A(KEYINPUT71), .B1(new_n205), .B2(new_n193), .ZN(new_n206));
  OAI211_X1 g020(.A(new_n192), .B(new_n194), .C1(new_n200), .C2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n193), .A2(G119), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n208), .B1(new_n205), .B2(new_n193), .ZN(new_n209));
  XNOR2_X1  g023(.A(KEYINPUT24), .B(G110), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n207), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT73), .ZN(new_n213));
  INV_X1    g027(.A(G140), .ZN(new_n214));
  AOI21_X1  g028(.A(KEYINPUT16), .B1(new_n214), .B2(G125), .ZN(new_n215));
  INV_X1    g029(.A(G125), .ZN(new_n216));
  NOR3_X1   g030(.A1(new_n216), .A2(KEYINPUT72), .A3(G140), .ZN(new_n217));
  XNOR2_X1  g031(.A(G125), .B(G140), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n217), .B1(new_n218), .B2(KEYINPUT72), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n215), .B1(new_n219), .B2(KEYINPUT16), .ZN(new_n220));
  INV_X1    g034(.A(G146), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n213), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n214), .A2(G125), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n216), .A2(G140), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n223), .A2(new_n224), .A3(KEYINPUT72), .ZN(new_n225));
  OR3_X1    g039(.A1(new_n216), .A2(KEYINPUT72), .A3(G140), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n225), .A2(new_n226), .A3(KEYINPUT16), .ZN(new_n227));
  INV_X1    g041(.A(new_n215), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n221), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(KEYINPUT73), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n218), .A2(new_n221), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n212), .A2(new_n222), .A3(new_n230), .A4(new_n231), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n194), .B1(new_n200), .B2(new_n206), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G110), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n227), .A2(new_n228), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G146), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n227), .A2(new_n221), .A3(new_n228), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n234), .B(new_n238), .C1(new_n209), .C2(new_n210), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n232), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G953), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n241), .A2(G221), .A3(G234), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n242), .B(KEYINPUT75), .ZN(new_n243));
  XNOR2_X1  g057(.A(KEYINPUT22), .B(G137), .ZN(new_n244));
  XNOR2_X1  g058(.A(new_n243), .B(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n240), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT74), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n240), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n232), .A2(new_n239), .A3(KEYINPUT74), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n245), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n247), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n191), .B1(new_n253), .B2(G902), .ZN(new_n254));
  AND3_X1   g068(.A1(new_n232), .A2(new_n239), .A3(KEYINPUT74), .ZN(new_n255));
  AOI21_X1  g069(.A(KEYINPUT74), .B1(new_n232), .B2(new_n239), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n252), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(new_n246), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n258), .A2(KEYINPUT25), .A3(new_n188), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n190), .B1(new_n254), .B2(new_n259), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n189), .A2(G902), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n253), .A2(new_n262), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(G137), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(KEYINPUT64), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT64), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(G137), .ZN(new_n269));
  AND2_X1   g083(.A1(KEYINPUT11), .A2(G134), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n267), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(KEYINPUT65), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT65), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n267), .A2(new_n269), .A3(new_n270), .A4(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n266), .A2(G134), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT11), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(G134), .ZN(new_n278));
  AOI21_X1  g092(.A(G131), .B1(new_n278), .B2(G137), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n272), .A2(new_n274), .A3(new_n277), .A4(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(KEYINPUT66), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n271), .A2(KEYINPUT65), .B1(new_n276), .B2(new_n275), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT66), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n282), .A2(new_n283), .A3(new_n274), .A4(new_n279), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g099(.A(G143), .B(G146), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n221), .A2(G143), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT1), .ZN(new_n288));
  AND3_X1   g102(.A1(new_n286), .A2(new_n288), .A3(G128), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n193), .B1(new_n287), .B2(KEYINPUT1), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n290), .A2(new_n286), .ZN(new_n291));
  INV_X1    g105(.A(new_n275), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n267), .A2(new_n269), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n292), .B1(new_n293), .B2(new_n278), .ZN(new_n294));
  INV_X1    g108(.A(G131), .ZN(new_n295));
  OAI22_X1  g109(.A1(new_n289), .A2(new_n291), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n285), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n278), .A2(G137), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n282), .A2(new_n274), .A3(new_n299), .ZN(new_n300));
  AOI22_X1  g114(.A1(new_n281), .A2(new_n284), .B1(G131), .B2(new_n300), .ZN(new_n301));
  NOR2_X1   g115(.A1(KEYINPUT0), .A2(G128), .ZN(new_n302));
  NAND2_X1  g116(.A1(KEYINPUT0), .A2(G128), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n302), .B1(new_n286), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G143), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G146), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n287), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n307), .A2(KEYINPUT0), .A3(G128), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n298), .B(KEYINPUT30), .C1(new_n301), .C2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT69), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n202), .A2(G116), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n195), .A2(new_n196), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n313), .B1(new_n314), .B2(G116), .ZN(new_n315));
  INV_X1    g129(.A(G113), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(KEYINPUT2), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT2), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G113), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n312), .B1(new_n315), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n203), .A2(G116), .A3(new_n204), .ZN(new_n322));
  INV_X1    g136(.A(new_n313), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n322), .A2(new_n320), .A3(new_n312), .A4(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  OAI22_X1  g139(.A1(new_n321), .A2(new_n325), .B1(new_n315), .B2(new_n320), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n311), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT67), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n300), .A2(G131), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n285), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n328), .B1(new_n330), .B2(new_n309), .ZN(new_n331));
  NOR3_X1   g145(.A1(new_n301), .A2(KEYINPUT67), .A3(new_n310), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n298), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT30), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n327), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n296), .B1(new_n281), .B2(new_n284), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n336), .B1(new_n330), .B2(new_n309), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n315), .A2(new_n320), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n322), .A2(new_n323), .A3(new_n320), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(KEYINPUT69), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n338), .B1(new_n324), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n337), .A2(new_n341), .ZN(new_n342));
  NOR2_X1   g156(.A1(G237), .A2(G953), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G210), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n344), .B(KEYINPUT27), .ZN(new_n345));
  XNOR2_X1  g159(.A(KEYINPUT26), .B(G101), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n345), .B(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n342), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(KEYINPUT31), .B1(new_n335), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n298), .B1(new_n301), .B2(new_n310), .ZN(new_n350));
  NOR3_X1   g164(.A1(new_n350), .A2(KEYINPUT28), .A3(new_n326), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT28), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n352), .B1(new_n337), .B2(new_n341), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n330), .A2(new_n328), .A3(new_n309), .ZN(new_n354));
  OAI21_X1  g168(.A(KEYINPUT67), .B1(new_n301), .B2(new_n310), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n336), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  OAI22_X1  g170(.A1(new_n351), .A2(new_n353), .B1(new_n356), .B2(new_n341), .ZN(new_n357));
  INV_X1    g171(.A(new_n347), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT31), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n350), .A2(new_n326), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n361), .A2(new_n358), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n356), .A2(KEYINPUT30), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n360), .B(new_n362), .C1(new_n363), .C2(new_n327), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n349), .A2(new_n359), .A3(new_n364), .ZN(new_n365));
  NOR2_X1   g179(.A1(G472), .A2(G902), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(KEYINPUT32), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT32), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n365), .A2(new_n369), .A3(new_n366), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n353), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n361), .A2(new_n352), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT70), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n350), .A2(new_n326), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT29), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n358), .A2(new_n377), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n374), .A2(new_n375), .A3(new_n376), .A4(new_n378), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n376), .B(new_n378), .C1(new_n351), .C2(new_n353), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT70), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n379), .A2(new_n188), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n357), .A2(new_n347), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n361), .A2(new_n347), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n384), .B1(new_n363), .B2(new_n327), .ZN(new_n385));
  AOI21_X1  g199(.A(KEYINPUT29), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(G472), .B1(new_n382), .B2(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n265), .B1(new_n371), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(G214), .B1(G237), .B2(G902), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT6), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT5), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n203), .A2(new_n391), .A3(G116), .A4(new_n204), .ZN(new_n392));
  AND2_X1   g206(.A1(new_n392), .A2(G113), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n322), .A2(KEYINPUT5), .A3(new_n323), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(G104), .ZN(new_n396));
  OAI21_X1  g210(.A(KEYINPUT3), .B1(new_n396), .B2(G107), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT3), .ZN(new_n398));
  INV_X1    g212(.A(G107), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n398), .A2(new_n399), .A3(G104), .ZN(new_n400));
  INV_X1    g214(.A(G101), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n396), .A2(G107), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n397), .A2(new_n400), .A3(new_n401), .A4(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n396), .A2(G107), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n399), .A2(G104), .ZN(new_n405));
  OAI21_X1  g219(.A(G101), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n395), .B(new_n408), .C1(new_n321), .C2(new_n325), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n397), .A2(new_n400), .A3(new_n402), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(G101), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n411), .A2(KEYINPUT4), .A3(new_n403), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT4), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n410), .A2(new_n413), .A3(G101), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n409), .B1(new_n341), .B2(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(G110), .B(G122), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n390), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  AND2_X1   g233(.A1(new_n412), .A2(new_n414), .ZN(new_n420));
  AOI22_X1  g234(.A1(new_n340), .A2(new_n324), .B1(new_n393), .B2(new_n394), .ZN(new_n421));
  AOI22_X1  g235(.A1(new_n326), .A2(new_n420), .B1(new_n421), .B2(new_n408), .ZN(new_n422));
  AOI21_X1  g236(.A(KEYINPUT80), .B1(new_n422), .B2(new_n417), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n409), .B(new_n417), .C1(new_n341), .C2(new_n415), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT80), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n419), .B1(new_n423), .B2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n416), .A2(new_n390), .A3(new_n418), .ZN(new_n428));
  OR2_X1    g242(.A1(new_n428), .A2(KEYINPUT81), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(KEYINPUT81), .ZN(new_n430));
  OR2_X1    g244(.A1(new_n290), .A2(new_n286), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n290), .A2(new_n286), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n431), .A2(new_n216), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n304), .A2(new_n308), .A3(G125), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n433), .A2(new_n434), .A3(KEYINPUT82), .ZN(new_n435));
  OR2_X1    g249(.A1(new_n434), .A2(KEYINPUT82), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n241), .A2(G224), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n438), .B(KEYINPUT83), .ZN(new_n439));
  XOR2_X1   g253(.A(new_n437), .B(new_n439), .Z(new_n440));
  NAND4_X1  g254(.A1(new_n427), .A2(new_n429), .A3(new_n430), .A4(new_n440), .ZN(new_n441));
  XOR2_X1   g255(.A(new_n417), .B(KEYINPUT8), .Z(new_n442));
  OR2_X1    g256(.A1(new_n421), .A2(new_n408), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n442), .B1(new_n443), .B2(new_n409), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT7), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n439), .A2(new_n445), .ZN(new_n446));
  AND2_X1   g260(.A1(new_n437), .A2(new_n446), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n437), .A2(new_n446), .ZN(new_n448));
  NOR3_X1   g262(.A1(new_n444), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n424), .B(new_n425), .ZN(new_n450));
  AOI21_X1  g264(.A(G902), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(G210), .B1(G237), .B2(G902), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n441), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  XOR2_X1   g267(.A(new_n452), .B(KEYINPUT84), .Z(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n455), .B1(new_n441), .B2(new_n451), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n453), .B1(new_n456), .B2(KEYINPUT85), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT85), .ZN(new_n458));
  AOI211_X1 g272(.A(new_n458), .B(new_n455), .C1(new_n441), .C2(new_n451), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n389), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(KEYINPUT9), .B(G234), .ZN(new_n461));
  OAI21_X1  g275(.A(G221), .B1(new_n461), .B2(G902), .ZN(new_n462));
  XNOR2_X1  g276(.A(G110), .B(G140), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n463), .A2(KEYINPUT76), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n463), .A2(KEYINPUT76), .ZN(new_n465));
  OR3_X1    g279(.A1(new_n464), .A2(new_n465), .A3(KEYINPUT77), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n241), .A2(G227), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n463), .B(KEYINPUT76), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(KEYINPUT77), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n466), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n467), .B1(new_n466), .B2(new_n469), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n412), .A2(new_n309), .A3(new_n414), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT78), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n412), .A2(new_n309), .A3(KEYINPUT78), .A4(new_n414), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n403), .B(new_n406), .C1(new_n289), .C2(new_n291), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(KEYINPUT10), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT10), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n408), .B(new_n480), .C1(new_n289), .C2(new_n291), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n483), .A2(new_n330), .ZN(new_n484));
  AOI22_X1  g298(.A1(new_n475), .A2(new_n476), .B1(new_n479), .B2(new_n481), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n485), .A2(new_n301), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n472), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n472), .B1(new_n485), .B2(new_n301), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n431), .A2(new_n407), .A3(new_n432), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n478), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n330), .A2(KEYINPUT12), .A3(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT12), .ZN(new_n492));
  AND2_X1   g306(.A1(new_n478), .A2(new_n489), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n492), .B1(new_n301), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n488), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(G902), .B1(new_n487), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(G469), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI22_X1  g313(.A1(new_n491), .A2(new_n494), .B1(new_n485), .B2(new_n301), .ZN(new_n500));
  INV_X1    g314(.A(new_n472), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n485), .A2(new_n301), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n501), .ZN(new_n503));
  OAI22_X1  g317(.A1(new_n500), .A2(new_n501), .B1(new_n503), .B2(new_n486), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n498), .B1(new_n504), .B2(new_n188), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n499), .B1(new_n505), .B2(KEYINPUT79), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n495), .A2(new_n502), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n483), .A2(new_n330), .ZN(new_n508));
  AOI22_X1  g322(.A1(new_n507), .A2(new_n472), .B1(new_n488), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(G469), .B1(new_n509), .B2(G902), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT79), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n462), .B1(new_n506), .B2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT20), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n343), .A2(G143), .A3(G214), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(G143), .B1(new_n343), .B2(G214), .ZN(new_n517));
  OAI21_X1  g331(.A(G131), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n343), .A2(G214), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(new_n305), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n520), .A2(new_n295), .A3(new_n515), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT17), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n518), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n520), .A2(new_n515), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n524), .A2(KEYINPUT17), .A3(G131), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n236), .A2(new_n523), .A3(new_n237), .A4(new_n525), .ZN(new_n526));
  XNOR2_X1  g340(.A(G113), .B(G122), .ZN(new_n527));
  XNOR2_X1  g341(.A(KEYINPUT87), .B(G104), .ZN(new_n528));
  OR2_X1    g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n527), .A2(new_n528), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(KEYINPUT89), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT89), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n529), .A2(new_n533), .A3(new_n530), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n219), .A2(G146), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n231), .ZN(new_n537));
  AND2_X1   g351(.A1(KEYINPUT18), .A2(G131), .ZN(new_n538));
  OR2_X1    g352(.A1(new_n524), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n524), .A2(new_n538), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n537), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n526), .A2(new_n535), .A3(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  AND3_X1   g357(.A1(new_n537), .A2(new_n539), .A3(new_n540), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n229), .B(new_n213), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT86), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT19), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n218), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  AOI22_X1  g362(.A1(new_n225), .A2(new_n226), .B1(new_n218), .B2(KEYINPUT86), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n548), .B(new_n221), .C1(new_n549), .C2(new_n547), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n518), .A2(new_n521), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n544), .B1(new_n545), .B2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n531), .ZN(new_n554));
  OAI21_X1  g368(.A(KEYINPUT88), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n222), .A2(new_n230), .A3(new_n551), .A4(new_n550), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n554), .B1(new_n556), .B2(new_n541), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT88), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n543), .B1(new_n555), .B2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT90), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n514), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n557), .A2(new_n558), .ZN(new_n563));
  AOI211_X1 g377(.A(KEYINPUT88), .B(new_n554), .C1(new_n556), .C2(new_n541), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n542), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NOR2_X1   g379(.A1(G475), .A2(G902), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n562), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n565), .A2(new_n561), .A3(new_n514), .A4(new_n566), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT91), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n554), .B1(new_n526), .B2(new_n541), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n570), .B(new_n188), .C1(new_n543), .C2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(G475), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n188), .B1(new_n543), .B2(new_n571), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n573), .B1(new_n574), .B2(KEYINPUT91), .ZN(new_n575));
  AOI22_X1  g389(.A1(new_n568), .A2(new_n569), .B1(new_n572), .B2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(G478), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n577), .A2(KEYINPUT15), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(G122), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(G116), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT14), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT92), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n583), .B1(new_n580), .B2(G116), .ZN(new_n584));
  INV_X1    g398(.A(G116), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n585), .A2(KEYINPUT92), .A3(G122), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n582), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT93), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n581), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  AOI211_X1 g403(.A(KEYINPUT93), .B(new_n582), .C1(new_n584), .C2(new_n586), .ZN(new_n590));
  OAI21_X1  g404(.A(KEYINPUT94), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AND3_X1   g405(.A1(new_n585), .A2(KEYINPUT92), .A3(G122), .ZN(new_n592));
  AOI21_X1  g406(.A(KEYINPUT92), .B1(new_n585), .B2(G122), .ZN(new_n593));
  OAI21_X1  g407(.A(KEYINPUT14), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(KEYINPUT93), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT94), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n587), .A2(new_n588), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n595), .A2(new_n596), .A3(new_n597), .A4(new_n581), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n584), .A2(new_n582), .A3(new_n586), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n591), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(G107), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n305), .A2(G128), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n193), .A2(G143), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(G134), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n584), .A2(new_n586), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n606), .A2(new_n399), .A3(new_n581), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n601), .A2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT13), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n603), .A2(new_n611), .A3(G134), .ZN(new_n612));
  OR2_X1    g426(.A1(new_n605), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n607), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n399), .B1(new_n606), .B2(new_n581), .ZN(new_n615));
  OR2_X1    g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n605), .A2(new_n612), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n613), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n461), .A2(new_n187), .A3(G953), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n610), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n619), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n608), .B1(new_n600), .B2(G107), .ZN(new_n622));
  INV_X1    g436(.A(new_n618), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n579), .B1(new_n625), .B2(new_n188), .ZN(new_n626));
  AOI211_X1 g440(.A(G902), .B(new_n578), .C1(new_n620), .C2(new_n624), .ZN(new_n627));
  AOI211_X1 g441(.A(new_n188), .B(new_n241), .C1(G234), .C2(G237), .ZN(new_n628));
  XNOR2_X1  g442(.A(KEYINPUT21), .B(G898), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  OR2_X1    g444(.A1(KEYINPUT95), .A2(G952), .ZN(new_n631));
  NAND2_X1  g445(.A1(KEYINPUT95), .A2(G952), .ZN(new_n632));
  AOI21_X1  g446(.A(G953), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(G234), .ZN(new_n634));
  INV_X1    g448(.A(G237), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n633), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n630), .A2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NOR3_X1   g452(.A1(new_n626), .A2(new_n627), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n576), .A2(new_n639), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n460), .A2(new_n513), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n388), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(G101), .ZN(G3));
  NAND2_X1  g457(.A1(new_n365), .A2(new_n188), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(G472), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n264), .A2(new_n645), .A3(new_n367), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n462), .ZN(new_n648));
  AOI22_X1  g462(.A1(new_n510), .A2(new_n511), .B1(new_n498), .B2(new_n497), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n505), .A2(KEYINPUT79), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g465(.A(KEYINPUT33), .B1(new_n619), .B2(KEYINPUT96), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n625), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n625), .A2(new_n652), .ZN(new_n654));
  OAI21_X1  g468(.A(G478), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n577), .A2(new_n188), .ZN(new_n656));
  AOI21_X1  g470(.A(G902), .B1(new_n620), .B2(new_n624), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n656), .B1(new_n657), .B2(new_n577), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n576), .A2(new_n638), .A3(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n389), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n441), .A2(new_n451), .ZN(new_n662));
  INV_X1    g476(.A(new_n452), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n661), .B1(new_n664), .B2(new_n453), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n647), .A2(new_n651), .A3(new_n660), .A4(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT34), .B(G104), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G6));
  XNOR2_X1  g482(.A(new_n637), .B(KEYINPUT97), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n651), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n646), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n626), .A2(new_n627), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n575), .A2(new_n572), .ZN(new_n674));
  INV_X1    g488(.A(new_n566), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n514), .B1(new_n560), .B2(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n565), .A2(KEYINPUT20), .A3(new_n566), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n673), .A2(new_n674), .A3(new_n676), .A4(new_n677), .ZN(new_n678));
  AND3_X1   g492(.A1(new_n441), .A2(new_n451), .A3(new_n452), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n452), .B1(new_n441), .B2(new_n451), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n389), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n671), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT35), .B(G107), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G9));
  AOI21_X1  g499(.A(KEYINPUT25), .B1(new_n258), .B2(new_n188), .ZN(new_n686));
  AOI211_X1 g500(.A(new_n191), .B(G902), .C1(new_n257), .C2(new_n246), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n189), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT36), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n245), .A2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT98), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n693), .B1(new_n255), .B2(new_n256), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n249), .A2(new_n250), .A3(new_n692), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g510(.A(KEYINPUT99), .B1(new_n696), .B2(new_n261), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT99), .ZN(new_n698));
  AOI211_X1 g512(.A(new_n698), .B(new_n262), .C1(new_n694), .C2(new_n695), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n688), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n645), .A2(new_n701), .A3(new_n367), .ZN(new_n702));
  OR2_X1    g516(.A1(new_n702), .A2(KEYINPUT100), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(KEYINPUT100), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n703), .A2(new_n641), .A3(new_n704), .ZN(new_n705));
  XOR2_X1   g519(.A(KEYINPUT37), .B(G110), .Z(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G12));
  AOI21_X1  g521(.A(new_n262), .B1(new_n694), .B2(new_n695), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(KEYINPUT99), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n709), .A2(new_n260), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n710), .A2(new_n513), .ZN(new_n711));
  AND3_X1   g525(.A1(new_n365), .A2(new_n369), .A3(new_n366), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n369), .B1(new_n365), .B2(new_n366), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n387), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(G900), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n628), .A2(new_n715), .ZN(new_n716));
  AND2_X1   g530(.A1(new_n716), .A2(new_n636), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n717), .B1(new_n575), .B2(new_n572), .ZN(new_n718));
  AND3_X1   g532(.A1(new_n676), .A2(new_n718), .A3(new_n677), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n673), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n720), .A2(new_n681), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n711), .A2(new_n714), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G128), .ZN(G30));
  NOR2_X1   g537(.A1(new_n457), .A2(new_n459), .ZN(new_n724));
  XNOR2_X1  g538(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n725));
  OR2_X1    g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n724), .A2(new_n725), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT102), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n347), .B1(new_n335), .B2(new_n361), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(new_n384), .ZN(new_n732));
  INV_X1    g546(.A(new_n376), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n188), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g548(.A(G472), .B1(new_n731), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n735), .B1(new_n712), .B2(new_n713), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n565), .A2(KEYINPUT90), .ZN(new_n737));
  AOI22_X1  g551(.A1(new_n737), .A2(new_n514), .B1(new_n565), .B2(new_n566), .ZN(new_n738));
  INV_X1    g552(.A(new_n569), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n674), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n673), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n741), .A2(new_n701), .A3(new_n661), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n728), .A2(new_n729), .A3(new_n736), .A4(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n742), .A2(new_n726), .A3(new_n727), .ZN(new_n744));
  INV_X1    g558(.A(new_n736), .ZN(new_n745));
  OAI21_X1  g559(.A(KEYINPUT102), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  XOR2_X1   g560(.A(new_n717), .B(KEYINPUT39), .Z(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n513), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(KEYINPUT40), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n743), .A2(new_n746), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(KEYINPUT103), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT103), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n743), .A2(new_n746), .A3(new_n753), .A4(new_n750), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(new_n305), .ZN(G45));
  INV_X1    g570(.A(new_n659), .ZN(new_n757));
  INV_X1    g571(.A(new_n717), .ZN(new_n758));
  AND4_X1   g572(.A1(new_n740), .A2(new_n665), .A3(new_n757), .A4(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n711), .A2(new_n759), .A3(new_n714), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G146), .ZN(G48));
  NAND2_X1  g575(.A1(new_n508), .A2(new_n502), .ZN(new_n762));
  AOI22_X1  g576(.A1(new_n762), .A2(new_n472), .B1(new_n495), .B2(new_n488), .ZN(new_n763));
  OAI21_X1  g577(.A(G469), .B1(new_n763), .B2(G902), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n499), .A2(new_n764), .A3(new_n462), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n681), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n714), .A2(new_n660), .A3(new_n264), .A4(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(KEYINPUT41), .B(G113), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n767), .B(new_n768), .ZN(G15));
  INV_X1    g583(.A(new_n765), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n770), .A2(new_n669), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n714), .A2(new_n264), .A3(new_n771), .A4(new_n682), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G116), .ZN(G18));
  INV_X1    g587(.A(new_n714), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n766), .A2(new_n576), .A3(new_n639), .A4(new_n701), .ZN(new_n775));
  OAI21_X1  g589(.A(KEYINPUT104), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n710), .A2(new_n640), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT104), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n777), .A2(new_n714), .A3(new_n778), .A4(new_n766), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n776), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G119), .ZN(G21));
  NOR3_X1   g595(.A1(new_n576), .A2(new_n681), .A3(new_n672), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n733), .B1(new_n372), .B2(new_n373), .ZN(new_n783));
  OAI211_X1 g597(.A(new_n349), .B(new_n364), .C1(new_n347), .C2(new_n783), .ZN(new_n784));
  AOI22_X1  g598(.A1(new_n644), .A2(G472), .B1(new_n784), .B2(new_n366), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n782), .A2(new_n771), .A3(new_n264), .A4(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G122), .ZN(G24));
  NOR3_X1   g601(.A1(new_n576), .A2(new_n659), .A3(new_n717), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(new_n766), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n784), .A2(new_n366), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n645), .A2(new_n701), .A3(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT105), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n785), .A2(KEYINPUT105), .A3(new_n701), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n789), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(new_n216), .ZN(G27));
  NAND2_X1  g610(.A1(new_n714), .A2(new_n264), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n457), .A2(new_n459), .A3(new_n661), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n648), .B1(new_n499), .B2(new_n510), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n788), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  AND2_X1   g614(.A1(KEYINPUT106), .A2(KEYINPUT42), .ZN(new_n801));
  NOR2_X1   g615(.A1(KEYINPUT106), .A2(KEYINPUT42), .ZN(new_n802));
  OAI22_X1  g616(.A1(new_n797), .A2(new_n800), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n740), .A2(new_n757), .A3(new_n758), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n662), .A2(new_n454), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(new_n458), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n456), .A2(KEYINPUT85), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n806), .A2(new_n389), .A3(new_n807), .A4(new_n453), .ZN(new_n808));
  INV_X1    g622(.A(new_n799), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n804), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n802), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n388), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n803), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(G131), .ZN(G33));
  INV_X1    g628(.A(KEYINPUT107), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n798), .A2(new_n673), .A3(new_n719), .A4(new_n799), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n815), .B1(new_n797), .B2(new_n816), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n808), .A2(new_n809), .A3(new_n720), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n818), .A2(KEYINPUT107), .A3(new_n714), .A4(new_n264), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(G134), .ZN(G36));
  NAND2_X1  g635(.A1(new_n576), .A2(new_n757), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT43), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n822), .B(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n710), .B1(new_n367), .B2(new_n645), .ZN(new_n825));
  AOI21_X1  g639(.A(KEYINPUT44), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT45), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n498), .B1(new_n504), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n828), .B1(new_n827), .B2(new_n504), .ZN(new_n829));
  NAND2_X1  g643(.A1(G469), .A2(G902), .ZN(new_n830));
  AOI21_X1  g644(.A(KEYINPUT46), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n499), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n829), .A2(KEYINPUT46), .A3(new_n830), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(new_n462), .ZN(new_n836));
  NOR4_X1   g650(.A1(new_n826), .A2(new_n748), .A3(new_n808), .A4(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n824), .A2(KEYINPUT44), .A3(new_n825), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g653(.A(KEYINPUT108), .B(G137), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n839), .B(new_n840), .ZN(G39));
  INV_X1    g655(.A(KEYINPUT47), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n836), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n835), .A2(KEYINPUT47), .A3(new_n462), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NOR4_X1   g659(.A1(new_n714), .A2(new_n804), .A3(new_n264), .A4(new_n808), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(G140), .ZN(G42));
  OAI211_X1 g662(.A(new_n711), .B(new_n714), .C1(new_n759), .C2(new_n721), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n710), .A2(KEYINPUT111), .A3(new_n758), .ZN(new_n850));
  AND4_X1   g664(.A1(new_n740), .A2(new_n665), .A3(new_n673), .A4(new_n799), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT111), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n852), .B1(new_n701), .B2(new_n717), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n850), .A2(new_n851), .A3(new_n736), .A4(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n849), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(KEYINPUT112), .B1(new_n855), .B2(new_n795), .ZN(new_n856));
  INV_X1    g670(.A(new_n789), .ZN(new_n857));
  INV_X1    g671(.A(new_n794), .ZN(new_n858));
  AOI21_X1  g672(.A(KEYINPUT105), .B1(new_n785), .B2(new_n701), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n857), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT112), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n860), .A2(new_n861), .A3(new_n849), .A4(new_n854), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n856), .A2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT52), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n793), .A2(new_n794), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n651), .A2(new_n724), .A3(new_n389), .A4(new_n701), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT109), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n868), .B1(new_n626), .B2(new_n627), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n619), .B1(new_n610), .B2(new_n618), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n622), .A2(new_n623), .A3(new_n621), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n188), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(new_n578), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n657), .A2(new_n579), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n873), .A2(KEYINPUT109), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n869), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n676), .A2(new_n718), .A3(new_n677), .ZN(new_n877));
  OAI21_X1  g691(.A(KEYINPUT110), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT110), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n719), .A2(new_n879), .A3(new_n875), .A4(new_n869), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n867), .A2(new_n881), .ZN(new_n882));
  AOI22_X1  g696(.A1(new_n866), .A2(new_n810), .B1(new_n882), .B2(new_n714), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n740), .A2(new_n757), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n576), .A2(new_n876), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n460), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AOI22_X1  g700(.A1(new_n671), .A2(new_n886), .B1(new_n388), .B2(new_n641), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n883), .A2(new_n820), .A3(new_n705), .A4(new_n887), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n767), .A2(new_n772), .A3(new_n786), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n813), .A2(new_n889), .A3(new_n780), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n856), .A2(new_n862), .A3(KEYINPUT52), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n865), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT53), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT54), .ZN(new_n896));
  INV_X1    g710(.A(new_n855), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n864), .B1(new_n897), .B2(new_n860), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n898), .B1(new_n863), .B2(new_n864), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT113), .ZN(new_n900));
  OR2_X1    g714(.A1(new_n888), .A2(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n813), .A2(new_n889), .A3(KEYINPUT53), .A4(new_n780), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n902), .B1(new_n900), .B2(new_n888), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n899), .A2(new_n901), .A3(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n895), .A2(new_n896), .A3(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n899), .A2(new_n894), .A3(new_n891), .ZN(new_n906));
  INV_X1    g720(.A(new_n893), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n906), .B1(new_n907), .B2(new_n894), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n905), .B1(new_n908), .B2(new_n896), .ZN(new_n909));
  INV_X1    g723(.A(new_n636), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n808), .A2(new_n765), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n745), .A2(new_n264), .A3(new_n910), .A4(new_n911), .ZN(new_n912));
  OR3_X1    g726(.A1(new_n912), .A2(new_n740), .A3(new_n757), .ZN(new_n913));
  INV_X1    g727(.A(new_n866), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n824), .A2(new_n910), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n911), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n785), .A2(new_n264), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT115), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n770), .B(new_n661), .C1(new_n919), .C2(KEYINPUT50), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n918), .A2(new_n728), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n919), .A2(KEYINPUT50), .ZN(new_n922));
  OAI221_X1 g736(.A(new_n913), .B1(new_n914), .B2(new_n916), .C1(new_n921), .C2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT51), .ZN(new_n924));
  INV_X1    g738(.A(new_n764), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n832), .A2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT114), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n462), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n928), .B1(new_n927), .B2(new_n926), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n843), .A2(new_n844), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(new_n798), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n728), .A2(new_n920), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(new_n922), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n918), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  OR3_X1    g748(.A1(new_n923), .A2(new_n924), .A3(new_n934), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n924), .B1(new_n923), .B2(new_n934), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n916), .A2(new_n797), .ZN(new_n937));
  XOR2_X1   g751(.A(KEYINPUT116), .B(KEYINPUT48), .Z(new_n938));
  XNOR2_X1  g752(.A(new_n937), .B(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(new_n766), .ZN(new_n940));
  OAI221_X1 g754(.A(new_n633), .B1(new_n884), .B2(new_n912), .C1(new_n918), .C2(new_n940), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n935), .A2(new_n936), .A3(new_n942), .ZN(new_n943));
  OAI22_X1  g757(.A1(new_n909), .A2(new_n943), .B1(G952), .B2(G953), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n926), .B(KEYINPUT49), .Z(new_n945));
  NAND3_X1  g759(.A1(new_n264), .A2(new_n462), .A3(new_n389), .ZN(new_n946));
  OR4_X1    g760(.A1(new_n728), .A2(new_n945), .A3(new_n822), .A4(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n944), .B1(new_n736), .B2(new_n947), .ZN(G75));
  OR2_X1    g762(.A1(new_n241), .A2(G952), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT118), .Z(new_n950));
  AOI211_X1 g764(.A(new_n188), .B(new_n455), .C1(new_n895), .C2(new_n904), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n427), .A2(new_n430), .A3(new_n429), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(new_n440), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n953), .B(KEYINPUT55), .Z(new_n954));
  OR2_X1    g768(.A1(new_n954), .A2(KEYINPUT56), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n950), .B1(new_n951), .B2(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT117), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n188), .B1(new_n895), .B2(new_n904), .ZN(new_n958));
  AOI21_X1  g772(.A(KEYINPUT56), .B1(new_n958), .B2(G210), .ZN(new_n959));
  INV_X1    g773(.A(new_n954), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n957), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(G210), .ZN(new_n962));
  AOI211_X1 g776(.A(new_n962), .B(new_n188), .C1(new_n895), .C2(new_n904), .ZN(new_n963));
  OAI211_X1 g777(.A(KEYINPUT117), .B(new_n954), .C1(new_n963), .C2(KEYINPUT56), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n956), .B1(new_n961), .B2(new_n964), .ZN(G51));
  INV_X1    g779(.A(new_n950), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n830), .B(KEYINPUT57), .Z(new_n967));
  INV_X1    g781(.A(new_n905), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n896), .B1(new_n895), .B2(new_n904), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n967), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n763), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n829), .B(KEYINPUT119), .Z(new_n973));
  NAND2_X1  g787(.A1(new_n958), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n966), .B1(new_n972), .B2(new_n974), .ZN(G54));
  NAND3_X1  g789(.A1(new_n958), .A2(KEYINPUT58), .A3(G475), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n565), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n958), .A2(KEYINPUT58), .A3(G475), .A4(new_n560), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n966), .B1(new_n977), .B2(new_n978), .ZN(G60));
  NOR2_X1   g793(.A1(new_n653), .A2(new_n654), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(KEYINPUT120), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n656), .B(KEYINPUT59), .Z(new_n982));
  OAI211_X1 g796(.A(new_n981), .B(new_n982), .C1(new_n968), .C2(new_n969), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(new_n950), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n981), .B1(new_n909), .B2(new_n982), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n984), .A2(new_n985), .ZN(G63));
  XNOR2_X1  g800(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n187), .A2(new_n188), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n987), .B(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(KEYINPUT52), .B1(new_n856), .B2(new_n862), .ZN(new_n990));
  NOR3_X1   g804(.A1(new_n990), .A2(new_n890), .A3(new_n888), .ZN(new_n991));
  AOI21_X1  g805(.A(KEYINPUT53), .B1(new_n991), .B2(new_n892), .ZN(new_n992));
  AND3_X1   g806(.A1(new_n899), .A2(new_n901), .A3(new_n903), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n989), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n966), .B1(new_n994), .B2(new_n253), .ZN(new_n995));
  INV_X1    g809(.A(new_n989), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n996), .B1(new_n895), .B2(new_n904), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(new_n696), .ZN(new_n998));
  OAI211_X1 g812(.A(new_n995), .B(new_n998), .C1(KEYINPUT122), .C2(KEYINPUT61), .ZN(new_n999));
  OAI211_X1 g813(.A(KEYINPUT122), .B(new_n950), .C1(new_n997), .C2(new_n258), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT61), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n950), .B1(new_n997), .B2(new_n258), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n895), .A2(new_n904), .ZN(new_n1003));
  AND3_X1   g817(.A1(new_n1003), .A2(new_n696), .A3(new_n989), .ZN(new_n1004));
  OAI211_X1 g818(.A(new_n1000), .B(new_n1001), .C1(new_n1002), .C2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n999), .A2(new_n1005), .ZN(G66));
  AND2_X1   g820(.A1(new_n889), .A2(new_n780), .ZN(new_n1007));
  AND2_X1   g821(.A1(new_n887), .A2(new_n705), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(G224), .A2(G953), .ZN(new_n1010));
  OAI22_X1  g824(.A1(new_n1009), .A2(G953), .B1(new_n629), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n952), .B1(G898), .B2(new_n241), .ZN(new_n1012));
  XOR2_X1   g826(.A(new_n1011), .B(new_n1012), .Z(G69));
  OAI21_X1  g827(.A(new_n311), .B1(new_n356), .B2(KEYINPUT30), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n548), .B1(new_n549), .B2(new_n547), .ZN(new_n1015));
  XOR2_X1   g829(.A(new_n1015), .B(KEYINPUT123), .Z(new_n1016));
  XNOR2_X1  g830(.A(new_n1014), .B(new_n1016), .ZN(new_n1017));
  XOR2_X1   g831(.A(new_n1017), .B(KEYINPUT124), .Z(new_n1018));
  AOI21_X1  g832(.A(new_n808), .B1(new_n884), .B2(new_n885), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n388), .A2(new_n749), .A3(new_n1019), .ZN(new_n1020));
  XOR2_X1   g834(.A(new_n1020), .B(KEYINPUT125), .Z(new_n1021));
  NAND3_X1  g835(.A1(new_n839), .A2(new_n847), .A3(new_n1021), .ZN(new_n1022));
  AND2_X1   g836(.A1(new_n860), .A2(new_n849), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n752), .A2(new_n754), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g838(.A(KEYINPUT62), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND4_X1  g840(.A1(new_n752), .A2(KEYINPUT62), .A3(new_n754), .A4(new_n1023), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n1022), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n1018), .B1(new_n1028), .B2(G953), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n1017), .B1(G900), .B2(G953), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n836), .A2(new_n748), .ZN(new_n1031));
  NOR3_X1   g845(.A1(new_n797), .A2(new_n681), .A3(new_n741), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  AND3_X1   g847(.A1(new_n847), .A2(new_n813), .A3(new_n1033), .ZN(new_n1034));
  NAND4_X1  g848(.A1(new_n1034), .A2(new_n820), .A3(new_n839), .A4(new_n1023), .ZN(new_n1035));
  OAI21_X1  g849(.A(new_n1030), .B1(new_n1035), .B2(G953), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1029), .A2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g851(.A(new_n241), .B1(G227), .B2(G900), .ZN(new_n1038));
  XNOR2_X1  g852(.A(new_n1037), .B(new_n1038), .ZN(G72));
  NAND2_X1  g853(.A1(G472), .A2(G902), .ZN(new_n1040));
  XOR2_X1   g854(.A(new_n1040), .B(KEYINPUT63), .Z(new_n1041));
  XOR2_X1   g855(.A(new_n1041), .B(KEYINPUT126), .Z(new_n1042));
  OAI21_X1  g856(.A(new_n1042), .B1(new_n1035), .B2(new_n1009), .ZN(new_n1043));
  INV_X1    g857(.A(new_n385), .ZN(new_n1044));
  AOI21_X1  g858(.A(new_n966), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g859(.A1(new_n730), .A2(new_n385), .A3(new_n1041), .ZN(new_n1046));
  OAI21_X1  g860(.A(new_n1045), .B1(new_n908), .B2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g861(.A1(new_n1028), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1048));
  NAND2_X1  g862(.A1(new_n1048), .A2(new_n1042), .ZN(new_n1049));
  AOI21_X1  g863(.A(new_n730), .B1(new_n1049), .B2(KEYINPUT127), .ZN(new_n1050));
  INV_X1    g864(.A(KEYINPUT127), .ZN(new_n1051));
  NAND3_X1  g865(.A1(new_n1048), .A2(new_n1051), .A3(new_n1042), .ZN(new_n1052));
  AOI21_X1  g866(.A(new_n1047), .B1(new_n1050), .B2(new_n1052), .ZN(G57));
endmodule


