//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 0 1 0 0 0 1 0 0 0 1 0 1 0 0 1 0 1 0 0 1 1 1 0 0 0 1 1 1 0 1 1 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:33 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n768, new_n769, new_n770, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061;
  INV_X1    g000(.A(G237), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(new_n188), .A3(G210), .ZN(new_n189));
  XOR2_X1   g003(.A(new_n189), .B(KEYINPUT27), .Z(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT26), .B(G101), .ZN(new_n191));
  XOR2_X1   g005(.A(new_n190), .B(new_n191), .Z(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(G116), .B(G119), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT2), .B(G113), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  XOR2_X1   g011(.A(KEYINPUT2), .B(G113), .Z(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(new_n194), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  XNOR2_X1  g014(.A(G143), .B(G146), .ZN(new_n201));
  XNOR2_X1  g015(.A(KEYINPUT0), .B(G128), .ZN(new_n202));
  OAI21_X1  g016(.A(KEYINPUT64), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  AND2_X1   g017(.A1(KEYINPUT0), .A2(G128), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n201), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G146), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G143), .ZN(new_n207));
  INV_X1    g021(.A(G143), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  NOR2_X1   g024(.A1(KEYINPUT0), .A2(G128), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n204), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT64), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n210), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n203), .A2(new_n205), .A3(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G137), .ZN(new_n216));
  AND2_X1   g030(.A1(KEYINPUT66), .A2(G134), .ZN(new_n217));
  NOR2_X1   g031(.A1(KEYINPUT66), .A2(G134), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT67), .ZN(new_n220));
  XNOR2_X1  g034(.A(KEYINPUT65), .B(KEYINPUT11), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  AND3_X1   g036(.A1(new_n216), .A2(KEYINPUT11), .A3(G134), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n217), .A2(new_n218), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n223), .B1(new_n224), .B2(G137), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n220), .B1(new_n219), .B2(new_n221), .ZN(new_n227));
  OAI21_X1  g041(.A(G131), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  OR2_X1    g042(.A1(KEYINPUT66), .A2(G134), .ZN(new_n229));
  NAND2_X1  g043(.A1(KEYINPUT66), .A2(G134), .ZN(new_n230));
  AOI21_X1  g044(.A(G137), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  XOR2_X1   g045(.A(KEYINPUT65), .B(KEYINPUT11), .Z(new_n232));
  OAI21_X1  g046(.A(KEYINPUT67), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G131), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n233), .A2(new_n234), .A3(new_n222), .A4(new_n225), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n215), .B1(new_n228), .B2(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(KEYINPUT1), .B1(new_n208), .B2(G146), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n210), .A2(G128), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G128), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n207), .B(new_n209), .C1(KEYINPUT1), .C2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  OR2_X1    g055(.A1(new_n216), .A2(G134), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n234), .B1(new_n219), .B2(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  AND2_X1   g058(.A1(new_n235), .A2(new_n244), .ZN(new_n245));
  OAI211_X1 g059(.A(KEYINPUT68), .B(new_n200), .C1(new_n236), .C2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(KEYINPUT28), .ZN(new_n247));
  NOR3_X1   g061(.A1(new_n236), .A2(new_n245), .A3(new_n200), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n248), .A2(KEYINPUT68), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n200), .B1(new_n236), .B2(new_n245), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n247), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n248), .A2(KEYINPUT28), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n193), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT30), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n228), .A2(new_n235), .ZN(new_n255));
  INV_X1    g069(.A(new_n215), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n245), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n254), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NOR3_X1   g073(.A1(new_n236), .A2(new_n245), .A3(KEYINPUT30), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n200), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n200), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n257), .A2(new_n258), .A3(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n261), .A2(new_n192), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(KEYINPUT31), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT31), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n261), .A2(new_n266), .A3(new_n192), .A4(new_n263), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n253), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  NOR2_X1   g082(.A1(G472), .A2(G902), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT32), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n257), .A2(new_n258), .A3(new_n254), .ZN(new_n273));
  OAI21_X1  g087(.A(KEYINPUT30), .B1(new_n236), .B2(new_n245), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n262), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NOR3_X1   g089(.A1(new_n275), .A2(new_n192), .A3(new_n248), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT29), .ZN(new_n277));
  AOI21_X1  g091(.A(G902), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT68), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n263), .A2(new_n279), .A3(new_n250), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n280), .A2(KEYINPUT28), .A3(new_n246), .ZN(new_n281));
  INV_X1    g095(.A(new_n252), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n281), .A2(new_n277), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(new_n192), .ZN(new_n284));
  NOR3_X1   g098(.A1(new_n248), .A2(KEYINPUT70), .A3(KEYINPUT28), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT70), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT28), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n286), .B1(new_n263), .B2(new_n287), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT69), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n263), .A2(new_n290), .A3(new_n250), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n257), .A2(new_n258), .A3(KEYINPUT69), .A4(new_n262), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n291), .A2(KEYINPUT28), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n277), .B1(new_n289), .B2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n278), .B1(new_n284), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(G472), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n268), .A2(KEYINPUT32), .A3(new_n269), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n272), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  XOR2_X1   g112(.A(G119), .B(G128), .Z(new_n299));
  XNOR2_X1  g113(.A(KEYINPUT24), .B(G110), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(KEYINPUT72), .B1(new_n239), .B2(G119), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT23), .ZN(new_n303));
  OR2_X1    g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n303), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n304), .B(new_n305), .C1(G119), .C2(new_n239), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n301), .B1(new_n306), .B2(G110), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(KEYINPUT73), .B(G125), .ZN(new_n309));
  NOR3_X1   g123(.A1(new_n309), .A2(KEYINPUT16), .A3(G140), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G140), .ZN(new_n312));
  INV_X1    g126(.A(G125), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(KEYINPUT73), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT73), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G125), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n312), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  NOR2_X1   g131(.A1(G125), .A2(G140), .ZN(new_n318));
  OAI211_X1 g132(.A(KEYINPUT74), .B(KEYINPUT16), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n318), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n321), .B1(new_n309), .B2(new_n312), .ZN(new_n322));
  AOI21_X1  g136(.A(KEYINPUT74), .B1(new_n322), .B2(KEYINPUT16), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n311), .B1(new_n320), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(new_n206), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT74), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n314), .A2(new_n316), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n318), .B1(new_n327), .B2(G140), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT16), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n326), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(new_n319), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(G146), .A3(new_n311), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n308), .B1(new_n325), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n299), .A2(new_n300), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n334), .B1(new_n306), .B2(G110), .ZN(new_n335));
  XNOR2_X1  g149(.A(G125), .B(G140), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n336), .B(KEYINPUT75), .ZN(new_n337));
  OR2_X1    g151(.A1(new_n337), .A2(G146), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  AOI211_X1 g153(.A(new_n206), .B(new_n310), .C1(new_n330), .C2(new_n319), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(KEYINPUT76), .B1(new_n333), .B2(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(G146), .B1(new_n331), .B2(new_n311), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n307), .B1(new_n343), .B2(new_n340), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT76), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n332), .A2(new_n338), .A3(new_n335), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  XNOR2_X1  g161(.A(KEYINPUT22), .B(G137), .ZN(new_n348));
  INV_X1    g162(.A(G221), .ZN(new_n349));
  INV_X1    g163(.A(G234), .ZN(new_n350));
  NOR3_X1   g164(.A1(new_n349), .A2(new_n350), .A3(G953), .ZN(new_n351));
  XOR2_X1   g165(.A(new_n348), .B(new_n351), .Z(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n342), .A2(new_n347), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n344), .A2(new_n346), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n355), .A2(KEYINPUT76), .A3(new_n352), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(G217), .B1(new_n350), .B2(G902), .ZN(new_n359));
  INV_X1    g173(.A(G902), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n357), .A2(new_n360), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT77), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT25), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(G902), .B1(new_n354), .B2(new_n356), .ZN(new_n367));
  OAI21_X1  g181(.A(KEYINPUT25), .B1(new_n367), .B2(KEYINPUT77), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  XOR2_X1   g183(.A(new_n359), .B(KEYINPUT71), .Z(new_n370));
  AOI21_X1  g184(.A(new_n362), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n298), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT78), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n298), .A2(KEYINPUT78), .A3(new_n371), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n215), .A2(new_n327), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT85), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n215), .A2(KEYINPUT85), .A3(new_n327), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n237), .A2(G128), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n381), .A2(new_n201), .ZN(new_n382));
  INV_X1    g196(.A(new_n240), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n309), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n379), .A2(new_n380), .A3(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(G224), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n386), .A2(G953), .ZN(new_n387));
  XOR2_X1   g201(.A(new_n385), .B(new_n387), .Z(new_n388));
  INV_X1    g202(.A(KEYINPUT83), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT80), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT79), .ZN(new_n391));
  INV_X1    g205(.A(G107), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(new_n392), .A3(G104), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(KEYINPUT3), .ZN(new_n394));
  INV_X1    g208(.A(G101), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT3), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n391), .A2(new_n396), .A3(new_n392), .A4(G104), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n392), .A2(G104), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n394), .A2(new_n395), .A3(new_n397), .A4(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(KEYINPUT4), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n398), .B1(new_n393), .B2(KEYINPUT3), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n395), .B1(new_n402), .B2(new_n397), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n390), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n394), .A2(new_n397), .A3(new_n399), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(G101), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n406), .A2(KEYINPUT80), .A3(KEYINPUT4), .A4(new_n400), .ZN(new_n407));
  AND2_X1   g221(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT4), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n405), .A2(new_n409), .A3(G101), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n200), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n389), .B1(new_n408), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(G119), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(G116), .ZN(new_n414));
  INV_X1    g228(.A(G116), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(G119), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n414), .A2(new_n416), .A3(KEYINPUT5), .ZN(new_n417));
  OR3_X1    g231(.A1(new_n415), .A2(KEYINPUT5), .A3(G119), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n417), .A2(new_n418), .A3(G113), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(new_n199), .ZN(new_n420));
  INV_X1    g234(.A(G104), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n421), .A2(G107), .ZN(new_n422));
  OAI21_X1  g236(.A(G101), .B1(new_n422), .B2(new_n398), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n400), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT81), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT81), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n400), .A2(new_n426), .A3(new_n423), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n420), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n411), .B1(new_n404), .B2(new_n407), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n428), .B1(new_n429), .B2(KEYINPUT83), .ZN(new_n430));
  XNOR2_X1  g244(.A(G110), .B(G122), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n412), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(KEYINPUT6), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n412), .A2(new_n430), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n431), .B(KEYINPUT84), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n434), .A2(KEYINPUT6), .A3(new_n435), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n388), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(KEYINPUT7), .B1(new_n386), .B2(G953), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n379), .A2(new_n380), .A3(new_n384), .A4(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n384), .A2(KEYINPUT87), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT87), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n241), .A2(new_n444), .A3(new_n309), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n443), .A2(new_n377), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n440), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n424), .A2(new_n420), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n400), .A2(new_n419), .A3(new_n199), .A4(new_n423), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  XOR2_X1   g264(.A(new_n431), .B(KEYINPUT8), .Z(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(KEYINPUT86), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT86), .ZN(new_n454));
  AOI211_X1 g268(.A(new_n454), .B(new_n451), .C1(new_n448), .C2(new_n449), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n442), .B(new_n447), .C1(new_n453), .C2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(KEYINPUT88), .ZN(new_n457));
  AND4_X1   g271(.A1(new_n400), .A2(new_n419), .A3(new_n199), .A4(new_n423), .ZN(new_n458));
  AOI22_X1  g272(.A1(new_n400), .A2(new_n423), .B1(new_n419), .B2(new_n199), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n452), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n454), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n450), .A2(KEYINPUT86), .A3(new_n452), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT88), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n463), .A2(new_n464), .A3(new_n442), .A4(new_n447), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n457), .A2(new_n432), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n360), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(KEYINPUT89), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT89), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n466), .A2(new_n469), .A3(new_n360), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n439), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(G210), .B1(G237), .B2(G902), .ZN(new_n472));
  XOR2_X1   g286(.A(new_n472), .B(KEYINPUT90), .Z(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(KEYINPUT91), .B1(new_n471), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n388), .ZN(new_n476));
  AOI22_X1  g290(.A1(new_n432), .A2(KEYINPUT6), .B1(new_n434), .B2(new_n435), .ZN(new_n477));
  INV_X1    g291(.A(new_n438), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  AND3_X1   g293(.A1(new_n466), .A2(new_n469), .A3(new_n360), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n469), .B1(new_n466), .B2(new_n360), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n474), .B(new_n479), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT91), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n483), .A2(new_n484), .A3(new_n473), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n475), .A2(new_n482), .A3(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(G214), .B1(G237), .B2(G902), .ZN(new_n487));
  XNOR2_X1  g301(.A(KEYINPUT93), .B(G475), .ZN(new_n488));
  MUX2_X1   g302(.A(new_n322), .B(new_n337), .S(new_n206), .Z(new_n489));
  NAND3_X1  g303(.A1(new_n187), .A2(new_n188), .A3(G214), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(new_n208), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n187), .A2(new_n188), .A3(G143), .A4(G214), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(KEYINPUT18), .A2(G131), .ZN(new_n494));
  XOR2_X1   g308(.A(new_n493), .B(new_n494), .Z(new_n495));
  NOR2_X1   g309(.A1(new_n489), .A2(new_n495), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n343), .A2(new_n340), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n493), .A2(G131), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT17), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n493), .B(new_n234), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n500), .B1(new_n501), .B2(new_n499), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n496), .B1(new_n497), .B2(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(G113), .B(G122), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n504), .B(G104), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(KEYINPUT94), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  OR2_X1    g321(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(G902), .B1(new_n503), .B2(new_n507), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n488), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT19), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n337), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n322), .A2(KEYINPUT19), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n501), .B1(new_n515), .B2(new_n206), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n332), .ZN(new_n517));
  OR2_X1    g331(.A1(new_n489), .A2(new_n495), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n517), .A2(new_n505), .A3(new_n518), .ZN(new_n519));
  OAI211_X1 g333(.A(KEYINPUT92), .B(new_n519), .C1(new_n503), .C2(new_n505), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT92), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n325), .A2(new_n332), .A3(new_n502), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n505), .B1(new_n522), .B2(new_n518), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n505), .B1(new_n489), .B2(new_n495), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n524), .B1(new_n516), .B2(new_n332), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n521), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g340(.A1(G475), .A2(G902), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n520), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  AND2_X1   g342(.A1(new_n528), .A2(KEYINPUT20), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n519), .B1(new_n503), .B2(new_n505), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT20), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n527), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n511), .B1(new_n529), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(G469), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n400), .A2(new_n423), .A3(new_n240), .A4(new_n238), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n424), .A2(new_n241), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(KEYINPUT82), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT82), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n424), .A2(new_n540), .A3(new_n241), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n537), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n255), .ZN(new_n543));
  OAI21_X1  g357(.A(KEYINPUT12), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n425), .A2(new_n427), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT10), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n241), .A2(new_n546), .ZN(new_n547));
  AOI22_X1  g361(.A1(new_n545), .A2(new_n547), .B1(new_n546), .B2(new_n536), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n404), .A2(new_n407), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n215), .B1(new_n409), .B2(new_n403), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n548), .A2(new_n551), .A3(new_n543), .ZN(new_n552));
  INV_X1    g366(.A(new_n541), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n540), .B1(new_n424), .B2(new_n241), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n536), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT12), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n555), .A2(new_n556), .A3(new_n255), .ZN(new_n557));
  XNOR2_X1  g371(.A(G110), .B(G140), .ZN(new_n558));
  AND2_X1   g372(.A1(new_n188), .A2(G227), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n558), .B(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n544), .A2(new_n552), .A3(new_n557), .A4(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n545), .A2(new_n547), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n536), .A2(new_n546), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n256), .A2(new_n410), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n567), .B1(new_n404), .B2(new_n407), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n255), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n561), .B1(new_n569), .B2(new_n552), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n535), .B(new_n360), .C1(new_n563), .C2(new_n570), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n535), .A2(new_n360), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n544), .A2(new_n552), .A3(new_n557), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n560), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n569), .A2(new_n552), .A3(new_n561), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n575), .A2(G469), .A3(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n571), .A2(new_n573), .A3(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(KEYINPUT9), .B(G234), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n349), .B1(new_n580), .B2(new_n360), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  XOR2_X1   g397(.A(G116), .B(G122), .Z(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(G107), .ZN(new_n585));
  XNOR2_X1  g399(.A(G116), .B(G122), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n392), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n208), .A2(G128), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT13), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n239), .A2(G143), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n589), .A2(new_n590), .ZN(new_n594));
  OAI21_X1  g408(.A(G134), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n224), .A2(new_n589), .A3(new_n592), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n588), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n589), .A2(new_n592), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n598), .B1(new_n218), .B2(new_n217), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n596), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n415), .A2(KEYINPUT14), .A3(G122), .ZN(new_n601));
  OAI211_X1 g415(.A(G107), .B(new_n601), .C1(new_n584), .C2(KEYINPUT14), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n600), .A2(new_n602), .A3(new_n587), .ZN(new_n603));
  INV_X1    g417(.A(G217), .ZN(new_n604));
  NOR3_X1   g418(.A1(new_n579), .A2(new_n604), .A3(G953), .ZN(new_n605));
  AND3_X1   g419(.A1(new_n597), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n605), .B1(new_n597), .B2(new_n603), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n608), .A2(G902), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT15), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(G478), .ZN(new_n611));
  AOI21_X1  g425(.A(KEYINPUT96), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  OR3_X1    g426(.A1(new_n608), .A2(KEYINPUT95), .A3(G902), .ZN(new_n613));
  OAI21_X1  g427(.A(KEYINPUT95), .B1(new_n608), .B2(G902), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n612), .B1(new_n615), .B2(new_n611), .ZN(new_n616));
  INV_X1    g430(.A(new_n611), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n613), .A2(KEYINPUT96), .A3(new_n617), .A4(new_n614), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n188), .A2(G952), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n620), .B1(G234), .B2(G237), .ZN(new_n621));
  AOI211_X1 g435(.A(new_n360), .B(new_n188), .C1(G234), .C2(G237), .ZN(new_n622));
  XNOR2_X1  g436(.A(KEYINPUT21), .B(G898), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n619), .A2(new_n625), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n534), .A2(new_n583), .A3(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n486), .A2(new_n487), .A3(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n376), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(G101), .ZN(G3));
  INV_X1    g445(.A(KEYINPUT97), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(G472), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n268), .A2(new_n360), .A3(new_n633), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n633), .B1(new_n268), .B2(new_n360), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n583), .ZN(new_n637));
  XOR2_X1   g451(.A(new_n608), .B(KEYINPUT33), .Z(new_n638));
  NAND3_X1  g452(.A1(new_n638), .A2(G478), .A3(new_n360), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n639), .B1(new_n615), .B2(G478), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n533), .B1(new_n528), .B2(KEYINPUT20), .ZN(new_n641));
  OAI211_X1 g455(.A(new_n640), .B(new_n625), .C1(new_n641), .C2(new_n510), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n636), .A2(new_n371), .A3(new_n637), .A4(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n487), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n483), .A2(new_n473), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n645), .B1(new_n646), .B2(new_n482), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(KEYINPUT34), .B(G104), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G6));
  NAND2_X1  g465(.A1(new_n528), .A2(KEYINPUT20), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n520), .A2(new_n526), .A3(new_n531), .A4(new_n527), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n510), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n619), .ZN(new_n655));
  AND3_X1   g469(.A1(new_n654), .A2(new_n655), .A3(new_n625), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n647), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n636), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n365), .B1(new_n363), .B2(new_n364), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n367), .A2(KEYINPUT77), .A3(KEYINPUT25), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n370), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n661), .B1(new_n358), .B2(new_n361), .ZN(new_n662));
  NOR4_X1   g476(.A1(new_n657), .A2(new_n658), .A3(new_n662), .A4(new_n583), .ZN(new_n663));
  XNOR2_X1  g477(.A(KEYINPUT35), .B(G107), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G9));
  INV_X1    g479(.A(KEYINPUT98), .ZN(new_n666));
  INV_X1    g480(.A(new_n370), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n667), .B1(new_n366), .B2(new_n368), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n353), .A2(KEYINPUT36), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n355), .B(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n361), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n666), .B1(new_n668), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n661), .A2(KEYINPUT98), .A3(new_n672), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n674), .A2(new_n675), .A3(new_n636), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n628), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(KEYINPUT37), .B(G110), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G12));
  NAND3_X1  g493(.A1(new_n674), .A2(new_n675), .A3(new_n298), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n647), .A2(new_n637), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n652), .A2(new_n653), .ZN(new_n682));
  INV_X1    g496(.A(G900), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n621), .B1(new_n622), .B2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n682), .A2(new_n655), .A3(new_n511), .A4(new_n685), .ZN(new_n686));
  NOR3_X1   g500(.A1(new_n680), .A2(new_n681), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(new_n239), .ZN(G30));
  NOR2_X1   g502(.A1(new_n668), .A2(new_n673), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n641), .A2(new_n510), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n690), .A2(new_n619), .ZN(new_n691));
  AND3_X1   g505(.A1(new_n689), .A2(new_n487), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n261), .A2(new_n263), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n192), .ZN(new_n694));
  AND2_X1   g508(.A1(new_n291), .A2(new_n292), .ZN(new_n695));
  OAI211_X1 g509(.A(new_n694), .B(new_n360), .C1(new_n192), .C2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(G472), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n272), .A2(new_n297), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n692), .A2(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT40), .ZN(new_n700));
  XNOR2_X1  g514(.A(KEYINPUT99), .B(KEYINPUT39), .ZN(new_n701));
  XOR2_X1   g515(.A(new_n684), .B(new_n701), .Z(new_n702));
  NOR2_X1   g516(.A1(new_n583), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n699), .B1(new_n700), .B2(new_n703), .ZN(new_n704));
  OR2_X1    g518(.A1(new_n486), .A2(KEYINPUT38), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n486), .A2(KEYINPUT38), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  OAI211_X1 g521(.A(new_n704), .B(new_n707), .C1(new_n700), .C2(new_n703), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G143), .ZN(G45));
  INV_X1    g523(.A(KEYINPUT101), .ZN(new_n710));
  AOI211_X1 g524(.A(new_n645), .B(new_n583), .C1(new_n646), .C2(new_n482), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n711), .A2(new_n298), .A3(new_n674), .A4(new_n675), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT100), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n534), .A2(new_n713), .A3(new_n640), .A4(new_n685), .ZN(new_n714));
  OAI211_X1 g528(.A(new_n640), .B(new_n685), .C1(new_n641), .C2(new_n510), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(KEYINPUT100), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n710), .B1(new_n712), .B2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(new_n680), .ZN(new_n719));
  INV_X1    g533(.A(new_n717), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n719), .A2(KEYINPUT101), .A3(new_n711), .A4(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G146), .ZN(G48));
  AND3_X1   g537(.A1(new_n548), .A2(new_n551), .A3(new_n543), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n543), .B1(new_n548), .B2(new_n551), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n560), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n562), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n535), .B1(new_n727), .B2(new_n360), .ZN(new_n728));
  AOI211_X1 g542(.A(G469), .B(G902), .C1(new_n726), .C2(new_n562), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(KEYINPUT102), .B1(new_n730), .B2(new_n582), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT102), .ZN(new_n732));
  NOR4_X1   g546(.A1(new_n728), .A2(new_n729), .A3(new_n732), .A4(new_n581), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(new_n647), .ZN(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  AND2_X1   g550(.A1(new_n298), .A2(new_n371), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT103), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n736), .A2(new_n737), .A3(new_n738), .A4(new_n643), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n298), .A2(new_n371), .A3(new_n643), .ZN(new_n740));
  OAI21_X1  g554(.A(KEYINPUT103), .B1(new_n740), .B2(new_n735), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(KEYINPUT41), .B(G113), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n742), .B(new_n743), .ZN(G15));
  NAND3_X1  g558(.A1(new_n734), .A2(new_n298), .A3(new_n371), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n745), .A2(new_n657), .ZN(new_n746));
  XNOR2_X1  g560(.A(KEYINPUT104), .B(G116), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(G18));
  NOR2_X1   g562(.A1(new_n534), .A2(new_n626), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n734), .A2(new_n647), .A3(new_n749), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n750), .A2(new_n680), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(new_n413), .ZN(G21));
  NAND2_X1  g566(.A1(new_n647), .A2(new_n691), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n265), .A2(new_n267), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n192), .B1(new_n289), .B2(new_n293), .ZN(new_n755));
  OAI211_X1 g569(.A(KEYINPUT105), .B(new_n269), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n268), .A2(new_n360), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(G472), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n269), .B1(new_n754), .B2(new_n755), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT105), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n371), .A2(new_n756), .A3(new_n758), .A4(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(new_n731), .ZN(new_n763));
  INV_X1    g577(.A(new_n733), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n763), .A2(new_n625), .A3(new_n764), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n753), .A2(new_n762), .A3(new_n765), .ZN(new_n766));
  XOR2_X1   g580(.A(new_n766), .B(G122), .Z(G24));
  NAND2_X1  g581(.A1(new_n661), .A2(new_n672), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n768), .A2(new_n756), .A3(new_n758), .A4(new_n761), .ZN(new_n769));
  NOR3_X1   g583(.A1(new_n769), .A2(new_n735), .A3(new_n717), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(new_n313), .ZN(G27));
  AND3_X1   g585(.A1(new_n714), .A2(new_n716), .A3(KEYINPUT42), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n645), .B1(new_n471), .B2(new_n474), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n729), .A2(new_n572), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n576), .A2(KEYINPUT106), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n576), .A2(KEYINPUT106), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n775), .A2(G469), .A3(new_n575), .A4(new_n776), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n581), .B1(new_n774), .B2(new_n777), .ZN(new_n778));
  AND4_X1   g592(.A1(new_n475), .A2(new_n773), .A3(new_n485), .A4(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT107), .ZN(new_n780));
  AND3_X1   g594(.A1(new_n268), .A2(KEYINPUT32), .A3(new_n269), .ZN(new_n781));
  AOI21_X1  g595(.A(KEYINPUT32), .B1(new_n268), .B2(new_n269), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n780), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n272), .A2(KEYINPUT107), .A3(new_n297), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n783), .A2(new_n784), .A3(new_n296), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n772), .A2(new_n779), .A3(new_n785), .A4(new_n371), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n475), .A2(new_n773), .A3(new_n485), .A4(new_n778), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n372), .A2(new_n787), .A3(new_n717), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n786), .B1(new_n788), .B2(KEYINPUT42), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT108), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n786), .B(KEYINPUT108), .C1(new_n788), .C2(KEYINPUT42), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(new_n234), .ZN(G33));
  INV_X1    g608(.A(KEYINPUT109), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n686), .B(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n737), .A2(new_n779), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(KEYINPUT110), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT110), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n737), .A2(new_n779), .A3(new_n796), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G134), .ZN(G36));
  NAND4_X1  g616(.A1(new_n775), .A2(KEYINPUT45), .A3(new_n575), .A4(new_n776), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n575), .A2(new_n576), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT45), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n535), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n572), .B1(new_n803), .B2(new_n806), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n807), .A2(KEYINPUT46), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n571), .B1(new_n807), .B2(KEYINPUT46), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n582), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  OR2_X1    g624(.A1(new_n810), .A2(new_n702), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n690), .A2(new_n640), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT111), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT43), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n812), .A2(new_n813), .A3(KEYINPUT43), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n816), .A2(new_n658), .A3(new_n768), .A4(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT44), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n811), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n475), .A2(new_n773), .A3(new_n485), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n820), .B(new_n821), .C1(new_n819), .C2(new_n818), .ZN(new_n822));
  XOR2_X1   g636(.A(KEYINPUT112), .B(G137), .Z(new_n823));
  XNOR2_X1  g637(.A(new_n822), .B(new_n823), .ZN(G39));
  INV_X1    g638(.A(KEYINPUT47), .ZN(new_n825));
  OR2_X1    g639(.A1(new_n810), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n810), .A2(new_n825), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n717), .A2(new_n298), .A3(new_n371), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n828), .A2(new_n821), .A3(new_n829), .ZN(new_n830));
  XOR2_X1   g644(.A(KEYINPUT113), .B(G140), .Z(new_n831));
  XNOR2_X1  g645(.A(new_n830), .B(new_n831), .ZN(G42));
  NAND2_X1  g646(.A1(new_n785), .A2(new_n371), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n821), .A2(new_n734), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n816), .A2(new_n621), .A3(new_n817), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  OR2_X1    g650(.A1(new_n836), .A2(KEYINPUT48), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(KEYINPUT48), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n662), .A2(new_n698), .ZN(new_n839));
  AND4_X1   g653(.A1(new_n621), .A2(new_n839), .A3(new_n734), .A4(new_n821), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n534), .A2(new_n640), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n620), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n835), .A2(new_n762), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(new_n736), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n837), .B(new_n838), .C1(new_n845), .C2(KEYINPUT124), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n846), .B1(KEYINPUT124), .B2(new_n845), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n734), .A2(new_n645), .ZN(new_n848));
  XOR2_X1   g662(.A(new_n848), .B(KEYINPUT120), .Z(new_n849));
  INV_X1    g663(.A(new_n707), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n849), .A2(new_n850), .A3(new_n843), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT121), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT50), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n730), .B(KEYINPUT114), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT119), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n582), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n858), .B1(new_n857), .B2(new_n856), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n826), .A2(new_n827), .A3(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n860), .A2(new_n821), .A3(new_n843), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n834), .A2(new_n835), .ZN(new_n862));
  AND4_X1   g676(.A1(new_n768), .A2(new_n756), .A3(new_n758), .A4(new_n761), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n534), .A2(new_n640), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n840), .A2(new_n865), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n861), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n851), .A2(new_n852), .A3(KEYINPUT50), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n855), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n847), .B1(new_n869), .B2(KEYINPUT51), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n855), .A2(new_n868), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n866), .A2(new_n864), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT122), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n872), .B(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(KEYINPUT123), .B1(new_n871), .B2(new_n874), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n872), .B(KEYINPUT122), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT123), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n876), .A2(new_n877), .A3(new_n868), .A4(new_n855), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n861), .A2(KEYINPUT51), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n870), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT118), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n698), .A2(new_n689), .A3(new_n685), .A4(new_n778), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n882), .B1(new_n883), .B2(new_n753), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n646), .A2(new_n482), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n885), .A2(new_n487), .A3(new_n691), .ZN(new_n886));
  AND4_X1   g700(.A1(new_n661), .A2(new_n778), .A3(new_n672), .A4(new_n685), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n886), .A2(KEYINPUT118), .A3(new_n698), .A4(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n889), .B1(new_n718), .B2(new_n721), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n770), .A2(new_n687), .ZN(new_n891));
  AOI21_X1  g705(.A(KEYINPUT52), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n889), .ZN(new_n893));
  AND4_X1   g707(.A1(KEYINPUT52), .A2(new_n722), .A3(new_n891), .A4(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n792), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n737), .A2(new_n779), .A3(new_n720), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT42), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(KEYINPUT108), .B1(new_n899), .B2(new_n786), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n896), .A2(new_n900), .ZN(new_n901));
  OAI22_X1  g715(.A1(new_n750), .A2(new_n680), .B1(new_n745), .B2(new_n657), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n902), .A2(new_n766), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n903), .A2(new_n742), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n769), .A2(new_n787), .A3(new_n717), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n684), .B1(new_n616), .B2(new_n618), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n654), .A2(new_n582), .A3(new_n578), .A4(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n674), .A2(new_n675), .A3(new_n298), .A4(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n475), .A2(new_n773), .A3(new_n485), .ZN(new_n910));
  OAI21_X1  g724(.A(KEYINPUT116), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(KEYINPUT98), .B1(new_n661), .B2(new_n672), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n668), .A2(new_n666), .A3(new_n673), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT116), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n781), .A2(new_n782), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n907), .B1(new_n916), .B2(new_n296), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n914), .A2(new_n915), .A3(new_n917), .A4(new_n821), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n905), .B1(new_n911), .B2(new_n918), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n801), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n486), .A2(new_n487), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n921), .A2(new_n644), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n922), .B1(new_n376), .B2(new_n629), .ZN(new_n923));
  NOR4_X1   g737(.A1(new_n641), .A2(new_n619), .A3(new_n510), .A4(new_n624), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n636), .A2(new_n371), .A3(new_n637), .A4(new_n924), .ZN(new_n925));
  OAI22_X1  g739(.A1(new_n628), .A2(new_n676), .B1(new_n921), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(KEYINPUT115), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT115), .ZN(new_n928));
  OAI221_X1 g742(.A(new_n928), .B1(new_n921), .B2(new_n925), .C1(new_n628), .C2(new_n676), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n923), .A2(new_n927), .A3(new_n929), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n901), .A2(new_n904), .A3(new_n920), .A4(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(KEYINPUT53), .B1(new_n895), .B2(new_n931), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n801), .A2(new_n919), .A3(new_n742), .A4(new_n903), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n923), .A2(new_n927), .A3(new_n929), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n793), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n736), .A2(new_n863), .A3(new_n720), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT117), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n936), .B(new_n937), .C1(new_n686), .C2(new_n712), .ZN(new_n938));
  OAI21_X1  g752(.A(KEYINPUT117), .B1(new_n770), .B2(new_n687), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n940), .A2(new_n890), .A3(KEYINPUT52), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n722), .A2(new_n893), .A3(new_n891), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT52), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT53), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n935), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n932), .A2(KEYINPUT54), .A3(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n946), .B1(new_n895), .B2(new_n931), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n789), .A2(KEYINPUT53), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n933), .A2(new_n934), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(KEYINPUT54), .B1(new_n945), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n881), .A2(new_n948), .A3(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n954), .B1(G952), .B2(G953), .ZN(new_n955));
  INV_X1    g769(.A(new_n856), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n956), .A2(KEYINPUT49), .ZN(new_n957));
  NOR4_X1   g771(.A1(new_n957), .A2(new_n645), .A3(new_n581), .A4(new_n812), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n956), .A2(KEYINPUT49), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n958), .A2(new_n850), .A3(new_n839), .A4(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n955), .A2(new_n960), .ZN(G75));
  NAND3_X1  g775(.A1(new_n890), .A2(KEYINPUT52), .A3(new_n891), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n944), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(KEYINPUT53), .B1(new_n935), .B2(new_n963), .ZN(new_n964));
  AND3_X1   g778(.A1(new_n722), .A2(KEYINPUT52), .A3(new_n893), .ZN(new_n965));
  AOI22_X1  g779(.A1(new_n965), .A2(new_n940), .B1(new_n942), .B2(new_n943), .ZN(new_n966));
  INV_X1    g780(.A(new_n950), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n920), .A2(new_n930), .A3(new_n967), .A4(new_n904), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  OAI211_X1 g783(.A(G902), .B(new_n473), .C1(new_n964), .C2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT56), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n477), .A2(new_n478), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(new_n476), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT55), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n970), .A2(new_n971), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n974), .B1(new_n970), .B2(new_n971), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n188), .A2(G952), .ZN(new_n977));
  NOR3_X1   g791(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(G51));
  INV_X1    g792(.A(KEYINPUT54), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n979), .B1(new_n966), .B2(new_n968), .ZN(new_n980));
  OAI21_X1  g794(.A(KEYINPUT125), .B1(new_n964), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(KEYINPUT54), .B1(new_n964), .B2(new_n969), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT125), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n949), .A2(new_n983), .A3(new_n952), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n981), .A2(new_n982), .A3(new_n984), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n572), .B(KEYINPUT57), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n987), .A2(new_n727), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n964), .A2(new_n969), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n989), .A2(new_n360), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n990), .A2(new_n803), .A3(new_n806), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n977), .B1(new_n988), .B2(new_n991), .ZN(G54));
  NAND2_X1  g806(.A1(KEYINPUT58), .A2(G475), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n993), .B(KEYINPUT126), .Z(new_n994));
  NAND2_X1  g808(.A1(new_n990), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n520), .A2(new_n526), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g811(.A(new_n977), .ZN(new_n998));
  NAND4_X1  g812(.A1(new_n990), .A2(new_n526), .A3(new_n520), .A4(new_n994), .ZN(new_n999));
  AND3_X1   g813(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(G60));
  NAND2_X1  g814(.A1(G478), .A2(G902), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n1001), .B(KEYINPUT59), .Z(new_n1002));
  AOI21_X1  g816(.A(new_n1002), .B1(new_n948), .B2(new_n953), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n998), .B1(new_n1003), .B2(new_n638), .ZN(new_n1004));
  INV_X1    g818(.A(new_n1002), .ZN(new_n1005));
  AND2_X1   g819(.A1(new_n638), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n1004), .B1(new_n985), .B2(new_n1006), .ZN(G63));
  NAND2_X1  g821(.A1(G217), .A2(G902), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n1008), .B(KEYINPUT60), .Z(new_n1009));
  INV_X1    g823(.A(new_n1009), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n358), .B1(new_n989), .B2(new_n1010), .ZN(new_n1011));
  OAI211_X1 g825(.A(new_n670), .B(new_n1009), .C1(new_n964), .C2(new_n969), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1011), .A2(new_n998), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT61), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n1011), .A2(KEYINPUT61), .A3(new_n998), .A4(new_n1012), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1015), .A2(new_n1016), .ZN(G66));
  OAI21_X1  g831(.A(G953), .B1(new_n623), .B2(new_n386), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n930), .A2(new_n904), .ZN(new_n1019));
  INV_X1    g833(.A(new_n1019), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1018), .B1(new_n1020), .B2(G953), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n972), .B1(G898), .B2(new_n188), .ZN(new_n1022));
  XNOR2_X1  g836(.A(new_n1021), .B(new_n1022), .ZN(G69));
  AOI21_X1  g837(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n1024));
  INV_X1    g838(.A(new_n1024), .ZN(new_n1025));
  NOR2_X1   g839(.A1(new_n259), .A2(new_n260), .ZN(new_n1026));
  XOR2_X1   g840(.A(new_n515), .B(KEYINPUT127), .Z(new_n1027));
  XOR2_X1   g841(.A(new_n1026), .B(new_n1027), .Z(new_n1028));
  INV_X1    g842(.A(new_n1028), .ZN(new_n1029));
  NOR2_X1   g843(.A1(new_n683), .A2(new_n188), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n822), .A2(new_n830), .ZN(new_n1032));
  INV_X1    g846(.A(new_n801), .ZN(new_n1033));
  NOR3_X1   g847(.A1(new_n811), .A2(new_n753), .A3(new_n833), .ZN(new_n1034));
  NOR3_X1   g848(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  AND2_X1   g849(.A1(new_n940), .A2(new_n722), .ZN(new_n1036));
  NAND3_X1  g850(.A1(new_n1035), .A2(new_n901), .A3(new_n1036), .ZN(new_n1037));
  OAI21_X1  g851(.A(new_n1031), .B1(new_n1037), .B2(G953), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1036), .A2(new_n708), .ZN(new_n1039));
  OR2_X1    g853(.A1(new_n1039), .A2(KEYINPUT62), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n1039), .A2(KEYINPUT62), .ZN(new_n1041));
  NOR2_X1   g855(.A1(new_n534), .A2(new_n619), .ZN(new_n1042));
  OAI21_X1  g856(.A(new_n703), .B1(new_n841), .B2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g857(.A1(new_n1043), .A2(new_n910), .ZN(new_n1044));
  AOI21_X1  g858(.A(new_n1032), .B1(new_n376), .B2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g859(.A1(new_n1040), .A2(new_n1041), .A3(new_n1045), .ZN(new_n1046));
  AND2_X1   g860(.A1(new_n1046), .A2(new_n188), .ZN(new_n1047));
  OAI211_X1 g861(.A(new_n1025), .B(new_n1038), .C1(new_n1047), .C2(new_n1028), .ZN(new_n1048));
  AOI21_X1  g862(.A(new_n1028), .B1(new_n1046), .B2(new_n188), .ZN(new_n1049));
  INV_X1    g863(.A(new_n1038), .ZN(new_n1050));
  OAI21_X1  g864(.A(new_n1024), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n1048), .A2(new_n1051), .ZN(G72));
  NAND2_X1  g866(.A1(G472), .A2(G902), .ZN(new_n1053));
  XOR2_X1   g867(.A(new_n1053), .B(KEYINPUT63), .Z(new_n1054));
  OAI21_X1  g868(.A(new_n1054), .B1(new_n1046), .B2(new_n1019), .ZN(new_n1055));
  NAND3_X1  g869(.A1(new_n1055), .A2(new_n192), .A3(new_n693), .ZN(new_n1056));
  INV_X1    g870(.A(new_n276), .ZN(new_n1057));
  AND3_X1   g871(.A1(new_n1057), .A2(new_n694), .A3(new_n1054), .ZN(new_n1058));
  NAND3_X1  g872(.A1(new_n932), .A2(new_n947), .A3(new_n1058), .ZN(new_n1059));
  OAI21_X1  g873(.A(new_n1054), .B1(new_n1037), .B2(new_n1019), .ZN(new_n1060));
  AOI21_X1  g874(.A(new_n977), .B1(new_n1060), .B2(new_n276), .ZN(new_n1061));
  AND3_X1   g875(.A1(new_n1056), .A2(new_n1059), .A3(new_n1061), .ZN(G57));
endmodule


