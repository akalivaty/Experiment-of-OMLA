//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 1 1 1 1 0 0 1 0 0 1 0 0 1 0 1 0 0 0 0 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 0 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n657, new_n658, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n827,
    new_n828, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n872, new_n873, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945;
  XNOR2_X1  g000(.A(KEYINPUT31), .B(G50gat), .ZN(new_n202));
  INV_X1    g001(.A(G106gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G228gat), .ZN(new_n206));
  INV_X1    g005(.A(G233gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  OR2_X1    g008(.A1(G197gat), .A2(G204gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(G197gat), .A2(G204gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT22), .ZN(new_n212));
  NAND2_X1  g011(.A1(G211gat), .A2(G218gat), .ZN(new_n213));
  AOI22_X1  g012(.A1(new_n210), .A2(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n213), .ZN(new_n216));
  NOR2_X1   g015(.A1(G211gat), .A2(G218gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n215), .A2(KEYINPUT70), .A3(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT70), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n218), .B1(new_n214), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT29), .ZN(new_n225));
  XOR2_X1   g024(.A(G141gat), .B(G148gat), .Z(new_n226));
  INV_X1    g025(.A(G155gat), .ZN(new_n227));
  INV_X1    g026(.A(G162gat), .ZN(new_n228));
  OAI21_X1  g027(.A(KEYINPUT2), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(G141gat), .ZN(new_n231));
  INV_X1    g030(.A(G148gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT73), .ZN(new_n234));
  NAND2_X1  g033(.A1(G141gat), .A2(G148gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(G155gat), .B(G162gat), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n230), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n240));
  OAI211_X1 g039(.A(new_n226), .B(new_n229), .C1(new_n234), .C2(new_n237), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n239), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n224), .B1(new_n225), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n239), .A2(new_n241), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT29), .B1(new_n215), .B2(new_n219), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n246), .B1(new_n219), .B2(new_n215), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n245), .B1(new_n240), .B2(new_n247), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n209), .B1(new_n243), .B2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n220), .A2(new_n225), .A3(new_n222), .ZN(new_n250));
  OR2_X1    g049(.A1(new_n250), .A2(KEYINPUT78), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT3), .B1(new_n250), .B2(KEYINPUT78), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n245), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT71), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n223), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n220), .A2(KEYINPUT71), .A3(new_n222), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  AND2_X1   g056(.A1(new_n242), .A2(new_n225), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n208), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n249), .B1(new_n253), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(G22gat), .ZN(new_n261));
  INV_X1    g060(.A(G78gat), .ZN(new_n262));
  INV_X1    g061(.A(G22gat), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n249), .B(new_n263), .C1(new_n253), .C2(new_n259), .ZN(new_n264));
  AND3_X1   g063(.A1(new_n261), .A2(new_n262), .A3(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n262), .B1(new_n261), .B2(new_n264), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n205), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n261), .A2(new_n264), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(G78gat), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n261), .A2(new_n262), .A3(new_n264), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n269), .A2(new_n270), .A3(new_n204), .ZN(new_n271));
  AND2_X1   g070(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G8gat), .B(G36gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n273), .B(KEYINPUT72), .ZN(new_n274));
  XNOR2_X1  g073(.A(G64gat), .B(G92gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n274), .B(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(KEYINPUT27), .B(G183gat), .ZN(new_n278));
  INV_X1    g077(.A(G190gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT28), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n278), .A2(KEYINPUT28), .A3(new_n279), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(G183gat), .A2(G190gat), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(G169gat), .A2(G176gat), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(G169gat), .ZN(new_n289));
  INV_X1    g088(.A(G176gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n288), .B1(KEYINPUT26), .B2(new_n291), .ZN(new_n292));
  OR2_X1    g091(.A1(new_n291), .A2(KEYINPUT26), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n286), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n284), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT23), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n296), .B1(G169gat), .B2(G176gat), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT25), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n297), .A2(new_n298), .A3(new_n287), .ZN(new_n299));
  XNOR2_X1  g098(.A(KEYINPUT65), .B(G176gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n296), .A2(G169gat), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n299), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(G183gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(new_n279), .ZN(new_n304));
  NAND3_X1  g103(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n305));
  OAI211_X1 g104(.A(new_n304), .B(new_n305), .C1(new_n286), .C2(KEYINPUT24), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n302), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n295), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n287), .B1(new_n291), .B2(new_n296), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT66), .ZN(new_n310));
  NOR2_X1   g109(.A1(G169gat), .A2(G176gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(KEYINPUT23), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT66), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n312), .A2(new_n313), .A3(new_n287), .ZN(new_n314));
  AOI22_X1  g113(.A1(new_n310), .A2(new_n314), .B1(new_n296), .B2(new_n291), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n286), .A2(KEYINPUT67), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT67), .ZN(new_n317));
  AOI21_X1  g116(.A(KEYINPUT24), .B1(new_n285), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n319), .A2(new_n304), .A3(new_n305), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n298), .B1(new_n315), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(G226gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n322), .A2(new_n207), .ZN(new_n323));
  OAI22_X1  g122(.A1(new_n308), .A2(new_n321), .B1(KEYINPUT29), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n314), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n313), .B1(new_n312), .B2(new_n287), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n297), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  AND3_X1   g126(.A1(new_n319), .A2(new_n304), .A3(new_n305), .ZN(new_n328));
  OAI21_X1  g127(.A(KEYINPUT25), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  AOI22_X1  g128(.A1(new_n284), .A2(new_n294), .B1(new_n306), .B2(new_n302), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n329), .B(new_n330), .C1(new_n322), .C2(new_n207), .ZN(new_n331));
  AND3_X1   g130(.A1(new_n324), .A2(new_n223), .A3(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n257), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n333), .B1(new_n324), .B2(new_n331), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n277), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n324), .A2(new_n331), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(new_n257), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n324), .A2(new_n223), .A3(new_n331), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(new_n338), .A3(new_n276), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n335), .A2(new_n339), .A3(KEYINPUT30), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n337), .A2(new_n338), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT30), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n341), .A2(new_n342), .A3(new_n277), .ZN(new_n343));
  AND2_X1   g142(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT68), .ZN(new_n345));
  INV_X1    g144(.A(G127gat), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n346), .A2(G134gat), .ZN(new_n347));
  INV_X1    g146(.A(G134gat), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n348), .A2(G127gat), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n345), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n348), .A2(G127gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n346), .A2(G134gat), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n351), .A2(new_n352), .A3(KEYINPUT68), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT1), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n354), .B1(G113gat), .B2(G120gat), .ZN(new_n355));
  AND2_X1   g154(.A1(G113gat), .A2(G120gat), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n350), .A2(new_n353), .A3(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(G127gat), .B(G134gat), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n359), .B(KEYINPUT68), .C1(new_n356), .C2(new_n355), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n361), .A2(new_n241), .A3(new_n239), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(KEYINPUT4), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT4), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n361), .A2(new_n364), .A3(new_n241), .A4(new_n239), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT77), .ZN(new_n366));
  AND3_X1   g165(.A1(new_n365), .A2(KEYINPUT76), .A3(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n366), .B1(new_n365), .B2(KEYINPUT76), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n363), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n365), .A2(KEYINPUT76), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT77), .ZN(new_n371));
  INV_X1    g170(.A(new_n363), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n365), .A2(KEYINPUT76), .A3(new_n366), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n244), .A2(KEYINPUT3), .ZN(new_n375));
  INV_X1    g174(.A(new_n361), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n375), .A2(new_n376), .A3(new_n242), .ZN(new_n377));
  NAND2_X1  g176(.A1(G225gat), .A2(G233gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(KEYINPUT75), .B(KEYINPUT5), .ZN(new_n379));
  AND3_X1   g178(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n369), .A2(new_n374), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n363), .A2(new_n365), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n382), .A2(new_n378), .A3(new_n377), .ZN(new_n383));
  INV_X1    g182(.A(new_n379), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n376), .A2(new_n244), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT74), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n385), .A2(new_n386), .A3(new_n362), .ZN(new_n387));
  INV_X1    g186(.A(new_n378), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n376), .A2(new_n244), .A3(KEYINPUT74), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n387), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n383), .A2(new_n384), .A3(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(G1gat), .B(G29gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n392), .B(KEYINPUT0), .ZN(new_n393));
  XNOR2_X1  g192(.A(G57gat), .B(G85gat), .ZN(new_n394));
  XOR2_X1   g193(.A(new_n393), .B(new_n394), .Z(new_n395));
  NAND3_X1  g194(.A1(new_n381), .A2(new_n391), .A3(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT6), .ZN(new_n397));
  AND2_X1   g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n381), .A2(new_n391), .ZN(new_n399));
  INV_X1    g198(.A(new_n395), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n395), .B1(new_n381), .B2(new_n391), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT6), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n344), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n361), .B1(new_n308), .B2(new_n321), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n329), .A2(new_n330), .A3(new_n376), .ZN(new_n407));
  NAND2_X1  g206(.A1(G227gat), .A2(G233gat), .ZN(new_n408));
  XOR2_X1   g207(.A(new_n408), .B(KEYINPUT64), .Z(new_n409));
  NAND3_X1  g208(.A1(new_n406), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(KEYINPUT32), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT33), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  XOR2_X1   g212(.A(G15gat), .B(G43gat), .Z(new_n414));
  XNOR2_X1  g213(.A(G71gat), .B(G99gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n411), .A2(new_n413), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n406), .A2(new_n407), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(new_n408), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n409), .A2(KEYINPUT34), .ZN(new_n420));
  AOI22_X1  g219(.A1(new_n419), .A2(KEYINPUT34), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n416), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n410), .B(KEYINPUT32), .C1(new_n412), .C2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n417), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n421), .B1(new_n423), .B2(new_n417), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n272), .A2(new_n405), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n340), .A2(new_n343), .ZN(new_n429));
  AND4_X1   g228(.A1(new_n271), .A2(new_n267), .A3(new_n429), .A4(new_n427), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT79), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n401), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n403), .A2(KEYINPUT79), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n432), .A2(new_n398), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(KEYINPUT35), .B1(new_n434), .B2(new_n404), .ZN(new_n435));
  AOI22_X1  g234(.A1(new_n428), .A2(KEYINPUT35), .B1(new_n430), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n267), .A2(new_n271), .ZN(new_n437));
  AOI21_X1  g236(.A(KEYINPUT79), .B1(new_n399), .B2(new_n400), .ZN(new_n438));
  AOI211_X1 g237(.A(new_n431), .B(new_n395), .C1(new_n381), .C2(new_n391), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT40), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n369), .A2(new_n374), .A3(new_n377), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT39), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n442), .A2(new_n443), .A3(new_n388), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n395), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n387), .A2(new_n389), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n443), .B1(new_n446), .B2(new_n378), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n448), .B1(new_n442), .B2(new_n388), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n441), .B1(new_n445), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n442), .A2(new_n388), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(new_n447), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n452), .A2(KEYINPUT40), .A3(new_n395), .A4(new_n444), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n440), .A2(new_n450), .A3(new_n453), .A4(new_n344), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT80), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NOR3_X1   g255(.A1(new_n429), .A2(new_n438), .A3(new_n439), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n457), .A2(KEYINPUT80), .A3(new_n450), .A4(new_n453), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n437), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  XOR2_X1   g258(.A(KEYINPUT82), .B(KEYINPUT37), .Z(new_n460));
  AOI21_X1  g259(.A(new_n277), .B1(new_n341), .B2(new_n460), .ZN(new_n461));
  XOR2_X1   g260(.A(KEYINPUT81), .B(KEYINPUT38), .Z(new_n462));
  INV_X1    g261(.A(KEYINPUT37), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n463), .B1(new_n336), .B2(new_n224), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n324), .A2(new_n333), .A3(new_n331), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n462), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AOI22_X1  g265(.A1(new_n461), .A2(new_n466), .B1(new_n341), .B2(new_n277), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n434), .A2(new_n404), .A3(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT83), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n434), .A2(KEYINPUT83), .A3(new_n404), .A4(new_n467), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n461), .B1(new_n463), .B2(new_n341), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(new_n462), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n470), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n426), .ZN(new_n476));
  AND2_X1   g275(.A1(KEYINPUT69), .A2(KEYINPUT36), .ZN(new_n477));
  NOR2_X1   g276(.A1(KEYINPUT69), .A2(KEYINPUT36), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n476), .A2(new_n424), .A3(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n481), .B1(new_n427), .B2(new_n477), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n482), .B1(new_n272), .B2(new_n405), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n436), .B1(new_n475), .B2(new_n484), .ZN(new_n485));
  XOR2_X1   g284(.A(G43gat), .B(G50gat), .Z(new_n486));
  INV_X1    g285(.A(G36gat), .ZN(new_n487));
  AND2_X1   g286(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n488));
  NOR2_X1   g287(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(G29gat), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n491), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n486), .B1(new_n493), .B2(KEYINPUT15), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT15), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n490), .A2(new_n495), .A3(new_n492), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n493), .A2(KEYINPUT15), .A3(new_n486), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(G15gat), .B(G22gat), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT16), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n500), .B1(new_n501), .B2(G1gat), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n502), .B1(G1gat), .B2(new_n500), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(G8gat), .ZN(new_n504));
  INV_X1    g303(.A(G8gat), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n502), .B(new_n505), .C1(G1gat), .C2(new_n500), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n499), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT84), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT84), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n499), .A2(new_n507), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(G229gat), .A2(G233gat), .ZN(new_n513));
  INV_X1    g312(.A(new_n507), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n499), .A2(KEYINPUT17), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT17), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n516), .B1(new_n497), .B2(new_n498), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n514), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n512), .A2(new_n513), .A3(new_n518), .ZN(new_n519));
  NOR2_X1   g318(.A1(KEYINPUT85), .A2(KEYINPUT18), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(G113gat), .B(G141gat), .ZN(new_n522));
  INV_X1    g321(.A(G197gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n522), .B(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(KEYINPUT11), .B(G169gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n524), .B(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n526), .B(KEYINPUT12), .ZN(new_n527));
  AND3_X1   g326(.A1(new_n499), .A2(new_n510), .A3(new_n507), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n510), .B1(new_n499), .B2(new_n507), .ZN(new_n529));
  OAI22_X1  g328(.A1(new_n528), .A2(new_n529), .B1(new_n507), .B2(new_n499), .ZN(new_n530));
  XOR2_X1   g329(.A(new_n513), .B(KEYINPUT13), .Z(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n520), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n512), .A2(new_n518), .A3(new_n513), .A4(new_n533), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n521), .A2(new_n527), .A3(new_n532), .A4(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT86), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AND2_X1   g336(.A1(new_n534), .A2(new_n532), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n538), .A2(KEYINPUT86), .A3(new_n527), .A4(new_n521), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n521), .ZN(new_n541));
  INV_X1    g340(.A(new_n527), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n485), .A2(new_n545), .ZN(new_n546));
  XOR2_X1   g345(.A(G183gat), .B(G211gat), .Z(new_n547));
  INV_X1    g346(.A(G71gat), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n548), .A2(new_n262), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n549), .A2(KEYINPUT9), .ZN(new_n550));
  XNOR2_X1  g349(.A(G57gat), .B(G64gat), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT87), .ZN(new_n553));
  NOR2_X1   g352(.A1(G71gat), .A2(G78gat), .ZN(new_n554));
  OAI22_X1  g353(.A1(new_n551), .A2(new_n553), .B1(new_n549), .B2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n552), .B(new_n555), .ZN(new_n556));
  OR2_X1    g355(.A1(new_n556), .A2(KEYINPUT21), .ZN(new_n557));
  NAND2_X1  g356(.A1(G231gat), .A2(G233gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n557), .B(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(G127gat), .B(G155gat), .ZN(new_n560));
  XOR2_X1   g359(.A(new_n560), .B(KEYINPUT20), .Z(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n558), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n557), .B(new_n564), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n565), .A2(new_n561), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n547), .B1(new_n563), .B2(new_n566), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n507), .B1(new_n556), .B2(KEYINPUT21), .ZN(new_n568));
  XNOR2_X1  g367(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n565), .A2(new_n561), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n559), .A2(new_n562), .ZN(new_n572));
  INV_X1    g371(.A(new_n547), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  AND3_X1   g373(.A1(new_n567), .A2(new_n570), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n570), .B1(new_n567), .B2(new_n574), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AND2_X1   g376(.A1(G232gat), .A2(G233gat), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n578), .A2(KEYINPUT41), .ZN(new_n579));
  XNOR2_X1  g378(.A(G134gat), .B(G162gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT90), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT7), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(KEYINPUT90), .A2(KEYINPUT7), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n584), .A2(G85gat), .A3(G92gat), .A4(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(G85gat), .ZN(new_n587));
  INV_X1    g386(.A(G92gat), .ZN(new_n588));
  OAI211_X1 g387(.A(new_n582), .B(new_n583), .C1(new_n587), .C2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(G99gat), .A2(G106gat), .ZN(new_n590));
  AOI22_X1  g389(.A1(KEYINPUT8), .A2(new_n590), .B1(new_n587), .B2(new_n588), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n586), .A2(new_n589), .A3(new_n591), .ZN(new_n592));
  XOR2_X1   g391(.A(G99gat), .B(G106gat), .Z(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n592), .B(new_n594), .ZN(new_n595));
  AOI22_X1  g394(.A1(new_n499), .A2(new_n595), .B1(KEYINPUT41), .B2(new_n578), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT91), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n592), .B(new_n593), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n599), .B1(new_n515), .B2(new_n517), .ZN(new_n600));
  XNOR2_X1  g399(.A(G190gat), .B(G218gat), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n598), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n601), .B1(new_n598), .B2(new_n600), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n581), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n598), .A2(new_n600), .ZN(new_n606));
  INV_X1    g405(.A(new_n601), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT92), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n581), .B(KEYINPUT89), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n608), .A2(new_n609), .A3(new_n602), .A4(new_n610), .ZN(new_n611));
  AND2_X1   g410(.A1(new_n605), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n608), .A2(new_n602), .A3(new_n610), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(KEYINPUT92), .ZN(new_n614));
  INV_X1    g413(.A(new_n551), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n615), .B1(KEYINPUT9), .B2(new_n549), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(new_n555), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(new_n599), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n556), .A2(new_n595), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT10), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n556), .A2(new_n595), .A3(KEYINPUT10), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(G230gat), .A2(G233gat), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g424(.A(G120gat), .B(G148gat), .Z(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT93), .ZN(new_n627));
  XNOR2_X1  g426(.A(G176gat), .B(G204gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  AND2_X1   g428(.A1(new_n618), .A2(new_n619), .ZN(new_n630));
  OAI211_X1 g429(.A(new_n625), .B(new_n629), .C1(new_n630), .C2(new_n624), .ZN(new_n631));
  INV_X1    g430(.A(new_n629), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n630), .A2(new_n624), .ZN(new_n633));
  INV_X1    g432(.A(new_n624), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n634), .B1(new_n621), .B2(new_n622), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n632), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT94), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n631), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  OAI211_X1 g437(.A(KEYINPUT94), .B(new_n632), .C1(new_n633), .C2(new_n635), .ZN(new_n639));
  AND2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n577), .A2(new_n612), .A3(new_n614), .A4(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n546), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n402), .A2(new_n404), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g445(.A(new_n646), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g446(.A1(new_n644), .A2(new_n429), .ZN(new_n648));
  XOR2_X1   g447(.A(KEYINPUT16), .B(G8gat), .Z(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n650), .B1(new_n505), .B2(new_n648), .ZN(new_n651));
  MUX2_X1   g450(.A(new_n650), .B(new_n651), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g451(.A(G15gat), .B1(new_n644), .B2(new_n482), .ZN(new_n653));
  INV_X1    g452(.A(new_n427), .ZN(new_n654));
  OR2_X1    g453(.A1(new_n654), .A2(G15gat), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n653), .B1(new_n644), .B2(new_n655), .ZN(G1326gat));
  NOR2_X1   g455(.A1(new_n644), .A2(new_n272), .ZN(new_n657));
  XOR2_X1   g456(.A(KEYINPUT43), .B(G22gat), .Z(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(G1327gat));
  INV_X1    g458(.A(new_n577), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(new_n641), .ZN(new_n661));
  AND2_X1   g460(.A1(new_n612), .A2(new_n614), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(KEYINPUT95), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n546), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n645), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n666), .A2(new_n491), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT45), .ZN(new_n669));
  NOR2_X1   g468(.A1(KEYINPUT97), .A2(KEYINPUT44), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n670), .B1(new_n485), .B2(new_n662), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n612), .A2(new_n614), .ZN(new_n672));
  XOR2_X1   g471(.A(KEYINPUT97), .B(KEYINPUT44), .Z(new_n673));
  AOI21_X1  g472(.A(new_n483), .B1(new_n459), .B2(new_n474), .ZN(new_n674));
  OAI211_X1 g473(.A(new_n672), .B(new_n673), .C1(new_n674), .C2(new_n436), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n661), .A2(new_n545), .ZN(new_n676));
  XOR2_X1   g475(.A(new_n676), .B(KEYINPUT96), .Z(new_n677));
  NAND3_X1  g476(.A1(new_n671), .A2(new_n675), .A3(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(G29gat), .B1(new_n678), .B2(new_n645), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n669), .A2(new_n679), .ZN(G1328gat));
  NOR3_X1   g479(.A1(new_n665), .A2(G36gat), .A3(new_n429), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(KEYINPUT46), .ZN(new_n682));
  OAI21_X1  g481(.A(G36gat), .B1(new_n678), .B2(new_n429), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(G1329gat));
  NOR2_X1   g483(.A1(new_n654), .A2(G43gat), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT47), .ZN(new_n686));
  AOI22_X1  g485(.A1(new_n666), .A2(new_n685), .B1(KEYINPUT98), .B2(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(G43gat), .B1(new_n678), .B2(new_n482), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n686), .A2(KEYINPUT98), .ZN(new_n690));
  XOR2_X1   g489(.A(new_n689), .B(new_n690), .Z(G1330gat));
  OAI21_X1  g490(.A(G50gat), .B1(new_n678), .B2(new_n272), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT99), .ZN(new_n693));
  AOI21_X1  g492(.A(KEYINPUT48), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  OR2_X1    g493(.A1(new_n272), .A2(G50gat), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n692), .B1(new_n665), .B2(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n694), .B(new_n696), .ZN(G1331gat));
  NAND4_X1  g496(.A1(new_n662), .A2(new_n545), .A3(new_n577), .A4(new_n640), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n485), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(new_n667), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g500(.A(new_n429), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT100), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n699), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n705));
  XOR2_X1   g504(.A(new_n704), .B(new_n705), .Z(G1333gat));
  XOR2_X1   g505(.A(new_n427), .B(KEYINPUT102), .Z(new_n707));
  NAND2_X1  g506(.A1(new_n699), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(new_n548), .ZN(new_n709));
  INV_X1    g508(.A(new_n482), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n699), .A2(G71gat), .A3(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT101), .ZN(new_n712));
  AND2_X1   g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n711), .A2(new_n712), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n709), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g515(.A1(new_n699), .A2(new_n437), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g517(.A1(new_n577), .A2(new_n544), .A3(new_n641), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n671), .A2(new_n675), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(G85gat), .B1(new_n720), .B2(new_n645), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n475), .A2(new_n484), .ZN(new_n722));
  INV_X1    g521(.A(new_n436), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n662), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n577), .A2(new_n544), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n724), .A2(KEYINPUT103), .A3(KEYINPUT51), .A4(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT103), .ZN(new_n727));
  OAI211_X1 g526(.A(new_n672), .B(new_n725), .C1(new_n674), .C2(new_n436), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT51), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n728), .A2(new_n729), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT104), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n728), .A2(KEYINPUT104), .A3(new_n729), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  AND2_X1   g535(.A1(new_n731), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n667), .A2(new_n587), .A3(new_n640), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n721), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(KEYINPUT105), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT105), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n741), .B(new_n721), .C1(new_n737), .C2(new_n738), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n742), .ZN(G1336gat));
  NAND2_X1  g542(.A1(new_n640), .A2(new_n344), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n744), .A2(G92gat), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n746), .B1(new_n731), .B2(new_n736), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n671), .A2(new_n344), .A3(new_n675), .A4(new_n719), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(G92gat), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT52), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n728), .B(new_n729), .ZN(new_n752));
  AOI22_X1  g551(.A1(new_n752), .A2(new_n745), .B1(new_n748), .B2(G92gat), .ZN(new_n753));
  OAI22_X1  g552(.A1(new_n747), .A2(new_n751), .B1(new_n753), .B2(new_n750), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT106), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  OAI221_X1 g555(.A(KEYINPUT106), .B1(new_n753), .B2(new_n750), .C1(new_n747), .C2(new_n751), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(G1337gat));
  INV_X1    g557(.A(G99gat), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n427), .A2(new_n640), .A3(new_n759), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(KEYINPUT107), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n761), .B1(new_n731), .B2(new_n736), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n720), .A2(new_n482), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n763), .A2(new_n759), .ZN(new_n764));
  OR3_X1    g563(.A1(new_n762), .A2(new_n764), .A3(KEYINPUT108), .ZN(new_n765));
  OAI21_X1  g564(.A(KEYINPUT108), .B1(new_n762), .B2(new_n764), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(G1338gat));
  NAND4_X1  g566(.A1(new_n671), .A2(new_n437), .A3(new_n675), .A4(new_n719), .ZN(new_n768));
  AOI21_X1  g567(.A(KEYINPUT53), .B1(new_n768), .B2(G106gat), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n272), .A2(G106gat), .A3(new_n641), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n769), .B1(new_n737), .B2(new_n771), .ZN(new_n772));
  AND3_X1   g571(.A1(new_n768), .A2(KEYINPUT109), .A3(G106gat), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n752), .A2(new_n770), .ZN(new_n774));
  AOI21_X1  g573(.A(KEYINPUT109), .B1(new_n768), .B2(G106gat), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n773), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT53), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n772), .B1(new_n776), .B2(new_n777), .ZN(G1339gat));
  NOR2_X1   g577(.A1(new_n642), .A2(new_n544), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n621), .A2(new_n622), .A3(new_n634), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(KEYINPUT110), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT110), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n621), .A2(new_n782), .A3(new_n622), .A4(new_n634), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n781), .A2(new_n625), .A3(KEYINPUT54), .A4(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT54), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n629), .B1(new_n635), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT55), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n784), .A2(KEYINPUT55), .A3(new_n786), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n789), .A2(new_n631), .A3(new_n790), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n512), .A2(new_n518), .ZN(new_n792));
  OAI22_X1  g591(.A1(new_n792), .A2(new_n513), .B1(new_n530), .B2(new_n531), .ZN(new_n793));
  AOI22_X1  g592(.A1(new_n537), .A2(new_n539), .B1(new_n526), .B2(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n672), .A2(new_n791), .A3(new_n794), .ZN(new_n795));
  AOI22_X1  g594(.A1(new_n544), .A2(new_n791), .B1(new_n794), .B2(new_n640), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n795), .B1(new_n796), .B2(new_n672), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n779), .B1(new_n797), .B2(new_n660), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n272), .A2(new_n427), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n667), .A2(new_n429), .ZN(new_n800));
  OR3_X1    g599(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n801), .B(KEYINPUT113), .ZN(new_n802));
  INV_X1    g601(.A(G113gat), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n802), .A2(new_n803), .A3(new_n544), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT112), .ZN(new_n805));
  OAI21_X1  g604(.A(KEYINPUT111), .B1(new_n798), .B2(new_n437), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT111), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n789), .A2(new_n631), .A3(new_n790), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n808), .B1(new_n543), .B2(new_n540), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n526), .ZN(new_n810));
  AND3_X1   g609(.A1(new_n540), .A2(new_n640), .A3(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n662), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n577), .B1(new_n812), .B2(new_n795), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n807), .B(new_n272), .C1(new_n813), .C2(new_n779), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n806), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n800), .A2(new_n654), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n805), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(new_n816), .ZN(new_n818));
  AOI211_X1 g617(.A(KEYINPUT112), .B(new_n818), .C1(new_n806), .C2(new_n814), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n817), .A2(new_n819), .A3(new_n545), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n804), .B1(new_n820), .B2(new_n803), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(KEYINPUT114), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT114), .ZN(new_n823));
  OAI211_X1 g622(.A(new_n804), .B(new_n823), .C1(new_n820), .C2(new_n803), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(new_n824), .ZN(G1340gat));
  INV_X1    g624(.A(G120gat), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n802), .A2(new_n826), .A3(new_n640), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n817), .A2(new_n819), .A3(new_n641), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n827), .B1(new_n828), .B2(new_n826), .ZN(G1341gat));
  NOR2_X1   g628(.A1(new_n817), .A2(new_n819), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n660), .A2(new_n346), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT115), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n830), .A2(KEYINPUT115), .A3(new_n831), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n346), .B1(new_n801), .B2(new_n660), .ZN(new_n836));
  AND3_X1   g635(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(G1342gat));
  AOI21_X1  g636(.A(G134gat), .B1(KEYINPUT116), .B2(KEYINPUT56), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n430), .A2(new_n667), .A3(new_n672), .A4(new_n838), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n798), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g639(.A1(KEYINPUT116), .A2(KEYINPUT56), .ZN(new_n841));
  XOR2_X1   g640(.A(new_n840), .B(new_n841), .Z(new_n842));
  NOR3_X1   g641(.A1(new_n817), .A2(new_n819), .A3(new_n662), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n842), .B1(new_n843), .B2(new_n348), .ZN(G1343gat));
  INV_X1    g643(.A(KEYINPUT57), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n845), .B1(new_n798), .B2(new_n272), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT117), .ZN(new_n847));
  OAI211_X1 g646(.A(KEYINPUT57), .B(new_n437), .C1(new_n813), .C2(new_n779), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n798), .A2(new_n272), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n850), .A2(KEYINPUT117), .A3(KEYINPUT57), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n710), .A2(new_n800), .ZN(new_n852));
  AND3_X1   g651(.A1(new_n849), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n231), .B1(new_n853), .B2(new_n544), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n850), .A2(new_n852), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n855), .A2(G141gat), .A3(new_n545), .ZN(new_n856));
  OR3_X1    g655(.A1(new_n854), .A2(KEYINPUT58), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(KEYINPUT58), .B1(new_n854), .B2(new_n856), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(G1344gat));
  INV_X1    g658(.A(KEYINPUT119), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n846), .A2(new_n860), .A3(new_n848), .ZN(new_n861));
  OAI211_X1 g660(.A(KEYINPUT119), .B(new_n845), .C1(new_n798), .C2(new_n272), .ZN(new_n862));
  AND4_X1   g661(.A1(new_n640), .A2(new_n861), .A3(new_n852), .A4(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(KEYINPUT59), .B1(new_n863), .B2(new_n232), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n849), .A2(new_n851), .A3(new_n640), .A4(new_n852), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n232), .A2(KEYINPUT59), .ZN(new_n866));
  AND3_X1   g665(.A1(new_n865), .A2(KEYINPUT118), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(KEYINPUT118), .B1(new_n865), .B2(new_n866), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n864), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n640), .A2(new_n232), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n869), .B1(new_n855), .B2(new_n870), .ZN(G1345gat));
  AOI21_X1  g670(.A(new_n227), .B1(new_n853), .B2(new_n577), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n855), .A2(G155gat), .A3(new_n660), .ZN(new_n873));
  OR2_X1    g672(.A1(new_n872), .A2(new_n873), .ZN(G1346gat));
  NOR2_X1   g673(.A1(new_n662), .A2(new_n228), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n850), .A2(new_n672), .A3(new_n852), .ZN(new_n876));
  AOI22_X1  g675(.A1(new_n853), .A2(new_n875), .B1(new_n228), .B2(new_n876), .ZN(G1347gat));
  INV_X1    g676(.A(new_n798), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n799), .A2(new_n667), .A3(new_n429), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(G169gat), .B1(new_n881), .B2(new_n544), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n707), .A2(new_n645), .A3(new_n344), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n883), .B1(new_n806), .B2(new_n814), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n545), .A2(new_n289), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n882), .B1(new_n884), .B2(new_n885), .ZN(G1348gat));
  OAI21_X1  g685(.A(new_n290), .B1(new_n880), .B2(new_n641), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n887), .B(KEYINPUT120), .ZN(new_n888));
  INV_X1    g687(.A(new_n884), .ZN(new_n889));
  OR2_X1    g688(.A1(new_n641), .A2(new_n300), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(KEYINPUT121), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT121), .ZN(new_n893));
  OAI211_X1 g692(.A(new_n888), .B(new_n893), .C1(new_n889), .C2(new_n890), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n892), .A2(new_n894), .ZN(G1349gat));
  NAND3_X1  g694(.A1(new_n881), .A2(new_n278), .A3(new_n577), .ZN(new_n896));
  XOR2_X1   g695(.A(new_n896), .B(KEYINPUT122), .Z(new_n897));
  NOR2_X1   g696(.A1(new_n889), .A2(new_n660), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n898), .A2(new_n303), .ZN(new_n899));
  OAI21_X1  g698(.A(KEYINPUT60), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n896), .B(KEYINPUT122), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT60), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n901), .B(new_n902), .C1(new_n303), .C2(new_n898), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n900), .A2(new_n903), .ZN(G1350gat));
  INV_X1    g703(.A(KEYINPUT61), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n884), .A2(new_n672), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT123), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n906), .A2(new_n907), .A3(G190gat), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n907), .B1(new_n906), .B2(G190gat), .ZN(new_n910));
  OAI211_X1 g709(.A(KEYINPUT124), .B(new_n905), .C1(new_n909), .C2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(new_n910), .ZN(new_n912));
  XNOR2_X1  g711(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n912), .A2(new_n908), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n881), .A2(new_n279), .A3(new_n672), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n911), .A2(new_n914), .A3(new_n915), .ZN(G1351gat));
  NOR3_X1   g715(.A1(new_n710), .A2(new_n667), .A3(new_n429), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n850), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n918), .B(KEYINPUT125), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n919), .A2(new_n523), .A3(new_n544), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n861), .A2(new_n862), .A3(new_n917), .ZN(new_n921));
  OAI21_X1  g720(.A(G197gat), .B1(new_n921), .B2(new_n545), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(KEYINPUT126), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT126), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n920), .A2(new_n925), .A3(new_n922), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n926), .ZN(G1352gat));
  OAI21_X1  g726(.A(G204gat), .B1(new_n921), .B2(new_n641), .ZN(new_n928));
  NOR4_X1   g727(.A1(new_n710), .A2(G204gat), .A3(new_n667), .A4(new_n744), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n850), .A2(new_n929), .ZN(new_n930));
  XOR2_X1   g729(.A(new_n930), .B(KEYINPUT62), .Z(new_n931));
  NAND2_X1  g730(.A1(new_n928), .A2(new_n931), .ZN(G1353gat));
  INV_X1    g731(.A(G211gat), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n919), .A2(new_n933), .A3(new_n577), .ZN(new_n934));
  NAND4_X1  g733(.A1(new_n861), .A2(new_n577), .A3(new_n862), .A4(new_n917), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n935), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n936));
  AOI21_X1  g735(.A(KEYINPUT63), .B1(new_n935), .B2(G211gat), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n934), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT127), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  OAI211_X1 g739(.A(KEYINPUT127), .B(new_n934), .C1(new_n936), .C2(new_n937), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(G1354gat));
  INV_X1    g741(.A(G218gat), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n919), .A2(new_n943), .A3(new_n672), .ZN(new_n944));
  OAI21_X1  g743(.A(G218gat), .B1(new_n921), .B2(new_n662), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(G1355gat));
endmodule


