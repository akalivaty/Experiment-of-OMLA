//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 1 1 1 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 1 1 0 1 1 0 0 0 0 1 1 1 0 0 0 0 0 0 1 1 0 0 0 0 0 0 0 1 1 1 1 1 1 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:22 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1245, new_n1246, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  OAI21_X1  g0002(.A(G50), .B1(G58), .B2(G68), .ZN(new_n203));
  INV_X1    g0003(.A(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(G1), .A2(G13), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n204), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(new_n206), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT65), .ZN(new_n216));
  INV_X1    g0016(.A(G58), .ZN(new_n217));
  INV_X1    g0017(.A(G232), .ZN(new_n218));
  INV_X1    g0018(.A(G107), .ZN(new_n219));
  INV_X1    g0019(.A(G264), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n222));
  INV_X1    g0022(.A(G50), .ZN(new_n223));
  INV_X1    g0023(.A(G226), .ZN(new_n224));
  INV_X1    g0024(.A(G116), .ZN(new_n225));
  INV_X1    g0025(.A(G270), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT64), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n211), .B1(new_n221), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n208), .B(new_n214), .C1(new_n229), .C2(KEYINPUT1), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G68), .B(G77), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT66), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G87), .B(G97), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  AOI21_X1  g0047(.A(new_n205), .B1(G33), .B2(G41), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT67), .ZN(new_n249));
  AND2_X1   g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  NOR2_X1   g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n249), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT3), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n255), .A2(KEYINPUT67), .A3(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n252), .A2(new_n257), .A3(G1698), .ZN(new_n258));
  XNOR2_X1  g0058(.A(new_n258), .B(KEYINPUT68), .ZN(new_n259));
  AND2_X1   g0059(.A1(new_n259), .A2(G223), .ZN(new_n260));
  NOR3_X1   g0060(.A1(new_n250), .A2(new_n251), .A3(new_n249), .ZN(new_n261));
  AOI21_X1  g0061(.A(KEYINPUT67), .B1(new_n255), .B2(new_n256), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G1698), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n263), .A2(G222), .A3(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G77), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n265), .B1(new_n266), .B2(new_n263), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n248), .B1(new_n260), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n248), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G274), .ZN(new_n272));
  INV_X1    g0072(.A(new_n205), .ZN(new_n273));
  NAND2_X1  g0073(.A1(G33), .A2(G41), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  AOI22_X1  g0075(.A1(new_n271), .A2(G226), .B1(new_n275), .B2(new_n270), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n268), .A2(new_n276), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n277), .A2(G179), .ZN(new_n278));
  INV_X1    g0078(.A(G13), .ZN(new_n279));
  NOR3_X1   g0079(.A1(new_n279), .A2(new_n206), .A3(G1), .ZN(new_n280));
  NAND3_X1  g0080(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n205), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n209), .A2(G20), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n283), .A2(G50), .A3(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n279), .A2(G1), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G20), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n285), .B1(G50), .B2(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(G50), .A2(G58), .ZN(new_n289));
  INV_X1    g0089(.A(G68), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n206), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  XNOR2_X1  g0091(.A(new_n291), .B(KEYINPUT69), .ZN(new_n292));
  XNOR2_X1  g0092(.A(KEYINPUT8), .B(G58), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n206), .A2(G33), .ZN(new_n294));
  INV_X1    g0094(.A(G150), .ZN(new_n295));
  NOR2_X1   g0095(.A1(G20), .A2(G33), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  OAI22_X1  g0097(.A1(new_n293), .A2(new_n294), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  OR2_X1    g0098(.A1(new_n292), .A2(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n288), .B1(new_n299), .B2(new_n282), .ZN(new_n300));
  AOI21_X1  g0100(.A(G169), .B1(new_n268), .B2(new_n276), .ZN(new_n301));
  OR3_X1    g0101(.A1(new_n278), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n302), .A2(KEYINPUT70), .ZN(new_n303));
  NOR3_X1   g0103(.A1(new_n278), .A2(new_n301), .A3(new_n300), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT70), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G179), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n273), .A2(new_n274), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n308), .A2(new_n270), .A3(G274), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n269), .ZN(new_n310));
  INV_X1    g0110(.A(G244), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n263), .A2(G232), .ZN(new_n314));
  OAI22_X1  g0114(.A1(new_n314), .A2(G1698), .B1(new_n219), .B2(new_n263), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n315), .B1(G238), .B2(new_n259), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n307), .B(new_n313), .C1(new_n316), .C2(new_n308), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT71), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n283), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(KEYINPUT71), .B1(new_n280), .B2(new_n282), .ZN(new_n320));
  AND2_X1   g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n321), .A2(G77), .A3(new_n284), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n280), .A2(new_n266), .ZN(new_n323));
  OAI22_X1  g0123(.A1(new_n293), .A2(new_n297), .B1(new_n206), .B2(new_n266), .ZN(new_n324));
  XNOR2_X1  g0124(.A(KEYINPUT15), .B(G87), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n325), .A2(new_n294), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n282), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n322), .A2(new_n323), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n259), .A2(G238), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n252), .A2(new_n257), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n330), .A2(new_n218), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n331), .A2(new_n264), .B1(G107), .B2(new_n330), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n329), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n312), .B1(new_n333), .B2(new_n248), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n317), .B(new_n328), .C1(new_n334), .C2(G169), .ZN(new_n335));
  OAI211_X1 g0135(.A(G190), .B(new_n313), .C1(new_n316), .C2(new_n308), .ZN(new_n336));
  INV_X1    g0136(.A(new_n328), .ZN(new_n337));
  INV_X1    g0137(.A(G200), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n336), .B(new_n337), .C1(new_n334), .C2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n335), .A2(new_n339), .ZN(new_n340));
  OAI22_X1  g0140(.A1(new_n303), .A2(new_n306), .B1(KEYINPUT72), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n277), .A2(G200), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n268), .A2(G190), .A3(new_n276), .ZN(new_n343));
  XOR2_X1   g0143(.A(new_n300), .B(KEYINPUT9), .Z(new_n344));
  NAND3_X1  g0144(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(KEYINPUT10), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT10), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n342), .A2(new_n347), .A3(new_n344), .A4(new_n343), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n224), .A2(G1698), .ZN(new_n350));
  OAI221_X1 g0150(.A(new_n350), .B1(G223), .B2(G1698), .C1(new_n250), .C2(new_n251), .ZN(new_n351));
  NAND2_X1  g0151(.A1(G33), .A2(G87), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n248), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n271), .A2(G232), .B1(new_n275), .B2(new_n270), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n354), .A2(new_n355), .A3(G179), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n309), .B1(new_n310), .B2(new_n218), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n308), .B1(new_n351), .B2(new_n352), .ZN(new_n358));
  OAI21_X1  g0158(.A(G169), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  AND2_X1   g0159(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n282), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n217), .A2(new_n290), .ZN(new_n362));
  NOR2_X1   g0162(.A1(G58), .A2(G68), .ZN(new_n363));
  OAI21_X1  g0163(.A(G20), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n296), .A2(G159), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n255), .A2(new_n206), .A3(new_n256), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT7), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n255), .A2(KEYINPUT7), .A3(new_n206), .A4(new_n256), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n366), .B1(new_n371), .B2(G68), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n361), .B1(new_n372), .B2(KEYINPUT16), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n370), .A2(KEYINPUT76), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n250), .A2(new_n251), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT76), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n375), .A2(new_n376), .A3(KEYINPUT7), .A4(new_n206), .ZN(new_n377));
  AOI21_X1  g0177(.A(G20), .B1(new_n252), .B2(new_n257), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n374), .B(new_n377), .C1(new_n378), .C2(KEYINPUT7), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n366), .B1(new_n379), .B2(G68), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n373), .B1(new_n380), .B2(KEYINPUT16), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n293), .B1(new_n209), .B2(G20), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n382), .A2(new_n283), .B1(new_n280), .B2(new_n293), .ZN(new_n383));
  AOI211_X1 g0183(.A(KEYINPUT18), .B(new_n360), .C1(new_n381), .C2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT18), .ZN(new_n385));
  AOI21_X1  g0185(.A(KEYINPUT7), .B1(new_n330), .B2(new_n206), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n374), .A2(new_n377), .ZN(new_n387));
  OAI21_X1  g0187(.A(G68), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n366), .ZN(new_n389));
  AOI21_X1  g0189(.A(KEYINPUT16), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT7), .B1(new_n375), .B2(new_n206), .ZN(new_n391));
  INV_X1    g0191(.A(new_n370), .ZN(new_n392));
  OAI21_X1  g0192(.A(G68), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n393), .A2(KEYINPUT16), .A3(new_n389), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(new_n282), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n383), .B1(new_n390), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n356), .A2(new_n359), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n385), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n384), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(G190), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n354), .A2(new_n355), .A3(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n338), .B1(new_n357), .B2(new_n358), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n383), .B(new_n403), .C1(new_n390), .C2(new_n395), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT17), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n381), .A2(KEYINPUT17), .A3(new_n383), .A4(new_n403), .ZN(new_n407));
  AND2_X1   g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n340), .A2(KEYINPUT72), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n349), .A2(new_n399), .A3(new_n408), .A4(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(G238), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n309), .B1(new_n310), .B2(new_n411), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n252), .A2(new_n257), .A3(G232), .A4(G1698), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n252), .A2(new_n257), .A3(G226), .A4(new_n264), .ZN(new_n414));
  INV_X1    g0214(.A(G97), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n413), .B(new_n414), .C1(new_n254), .C2(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n412), .B1(new_n416), .B2(new_n248), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT13), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AOI211_X1 g0219(.A(KEYINPUT13), .B(new_n412), .C1(new_n416), .C2(new_n248), .ZN(new_n420));
  OAI21_X1  g0220(.A(G169), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT14), .ZN(new_n422));
  INV_X1    g0222(.A(new_n417), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT73), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n423), .A2(new_n424), .A3(KEYINPUT13), .ZN(new_n425));
  OAI21_X1  g0225(.A(KEYINPUT73), .B1(new_n417), .B2(new_n418), .ZN(new_n426));
  INV_X1    g0226(.A(new_n420), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n425), .A2(new_n426), .A3(G179), .A4(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT14), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n429), .B(G169), .C1(new_n419), .C2(new_n420), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n422), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n290), .A2(G20), .ZN(new_n432));
  OAI221_X1 g0232(.A(new_n432), .B1(new_n294), .B2(new_n266), .C1(new_n297), .C2(new_n223), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n282), .ZN(new_n434));
  XNOR2_X1  g0234(.A(new_n434), .B(KEYINPUT74), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(KEYINPUT11), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT74), .ZN(new_n437));
  XNOR2_X1  g0237(.A(new_n434), .B(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT11), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n432), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT12), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n441), .B(new_n286), .C1(KEYINPUT75), .C2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(KEYINPUT75), .ZN(new_n444));
  XNOR2_X1  g0244(.A(new_n443), .B(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n321), .A2(G68), .A3(new_n284), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n436), .A2(new_n440), .A3(new_n445), .A4(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n431), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n447), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n425), .A2(new_n426), .A3(G190), .A4(new_n427), .ZN(new_n450));
  OAI21_X1  g0250(.A(G200), .B1(new_n419), .B2(new_n420), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n448), .A2(new_n452), .ZN(new_n453));
  NOR3_X1   g0253(.A1(new_n341), .A2(new_n410), .A3(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(G45), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n456), .A2(G1), .ZN(new_n457));
  XNOR2_X1  g0257(.A(KEYINPUT5), .B(G41), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n275), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n457), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(new_n308), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n459), .B1(new_n461), .B2(new_n226), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n255), .A2(new_n256), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n220), .A2(new_n264), .ZN(new_n464));
  AOI22_X1  g0264(.A1(new_n330), .A2(G303), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(G257), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n466), .A2(G1698), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n467), .B1(new_n250), .B2(new_n251), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(KEYINPUT81), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT81), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n463), .A2(new_n470), .A3(new_n467), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n465), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n462), .B1(new_n473), .B2(new_n248), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(G179), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n308), .B1(new_n465), .B2(new_n472), .ZN(new_n476));
  OAI211_X1 g0276(.A(KEYINPUT21), .B(G169), .C1(new_n476), .C2(new_n462), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(G20), .B1(G33), .B2(G283), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n479), .B1(G33), .B2(new_n415), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n225), .A2(G20), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n480), .A2(new_n282), .A3(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT20), .ZN(new_n483));
  AND2_X1   g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n482), .A2(new_n483), .ZN(new_n485));
  INV_X1    g0285(.A(new_n286), .ZN(new_n486));
  OAI22_X1  g0286(.A1(new_n484), .A2(new_n485), .B1(new_n486), .B2(new_n481), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n254), .A2(G1), .ZN(new_n488));
  XNOR2_X1  g0288(.A(new_n488), .B(KEYINPUT78), .ZN(new_n489));
  AND4_X1   g0289(.A1(G116), .A2(new_n319), .A3(new_n320), .A4(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n478), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(KEYINPUT82), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT82), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n478), .A2(new_n495), .A3(new_n492), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(G169), .ZN(new_n498));
  NOR3_X1   g0298(.A1(new_n491), .A2(new_n474), .A3(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n499), .A2(KEYINPUT21), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n474), .A2(G190), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n502), .B(new_n491), .C1(new_n338), .C2(new_n474), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n497), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n206), .B(G87), .C1(new_n250), .C2(new_n251), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(KEYINPUT22), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT83), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n505), .A2(KEYINPUT83), .A3(KEYINPUT22), .ZN(new_n509));
  INV_X1    g0309(.A(G87), .ZN(new_n510));
  NOR3_X1   g0310(.A1(new_n510), .A2(KEYINPUT22), .A3(G20), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n508), .A2(new_n509), .B1(new_n263), .B2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT23), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n513), .B1(new_n206), .B2(G107), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n219), .A2(KEYINPUT23), .A3(G20), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(G33), .A2(G116), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n516), .B1(G20), .B2(new_n517), .ZN(new_n518));
  NOR3_X1   g0318(.A1(new_n512), .A2(KEYINPUT24), .A3(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT24), .ZN(new_n520));
  INV_X1    g0320(.A(new_n509), .ZN(new_n521));
  AOI21_X1  g0321(.A(KEYINPUT83), .B1(new_n505), .B2(KEYINPUT22), .ZN(new_n522));
  INV_X1    g0322(.A(new_n511), .ZN(new_n523));
  OAI22_X1  g0323(.A1(new_n521), .A2(new_n522), .B1(new_n330), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n518), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n520), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n282), .B1(new_n519), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n460), .A2(G264), .A3(new_n308), .ZN(new_n528));
  NOR2_X1   g0328(.A1(G250), .A2(G1698), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n529), .B1(new_n466), .B2(G1698), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n530), .A2(new_n463), .B1(G33), .B2(G294), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n528), .B(new_n459), .C1(new_n531), .C2(new_n308), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n338), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(G190), .B2(new_n532), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n280), .A2(KEYINPUT25), .A3(new_n219), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT84), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT25), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n537), .B1(new_n287), .B2(G107), .ZN(new_n538));
  OR2_X1    g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n536), .A2(new_n538), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n489), .A2(new_n283), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n539), .A2(new_n540), .B1(new_n542), .B2(G107), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n527), .A2(new_n534), .A3(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n287), .A2(G97), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n545), .B1(new_n542), .B2(G97), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n296), .A2(G77), .ZN(new_n547));
  XNOR2_X1  g0347(.A(new_n547), .B(KEYINPUT77), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT6), .ZN(new_n549));
  NOR3_X1   g0349(.A1(new_n549), .A2(new_n415), .A3(G107), .ZN(new_n550));
  XNOR2_X1  g0350(.A(G97), .B(G107), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n550), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n548), .B1(new_n206), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n553), .B1(new_n379), .B2(G107), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n546), .B1(new_n554), .B2(new_n361), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n459), .B1(new_n461), .B2(new_n466), .ZN(new_n556));
  OAI211_X1 g0356(.A(G244), .B(new_n264), .C1(new_n250), .C2(new_n251), .ZN(new_n557));
  XNOR2_X1  g0357(.A(KEYINPUT79), .B(KEYINPUT4), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n557), .A2(new_n558), .B1(G33), .B2(G283), .ZN(new_n559));
  AND2_X1   g0359(.A1(KEYINPUT4), .A2(G244), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n252), .A2(new_n257), .A3(new_n264), .A4(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(G250), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n559), .B(new_n561), .C1(new_n562), .C2(new_n258), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n556), .B1(new_n563), .B2(new_n248), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n307), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n555), .B(new_n565), .C1(G169), .C2(new_n564), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n206), .B1(new_n261), .B2(new_n262), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n368), .ZN(new_n568));
  XNOR2_X1  g0368(.A(new_n370), .B(new_n376), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n219), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n282), .B1(new_n570), .B2(new_n553), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n564), .A2(G200), .ZN(new_n572));
  AOI211_X1 g0372(.A(G190), .B(new_n556), .C1(new_n563), .C2(new_n248), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n571), .B(new_n546), .C1(new_n572), .C2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n544), .A2(new_n566), .A3(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n532), .A2(G179), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n576), .B1(new_n498), .B2(new_n532), .ZN(new_n577));
  OAI21_X1  g0377(.A(KEYINPUT24), .B1(new_n512), .B2(new_n518), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n524), .A2(new_n520), .A3(new_n525), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n361), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n543), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n577), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n206), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n510), .A2(new_n415), .A3(new_n219), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n206), .B(G68), .C1(new_n250), .C2(new_n251), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT19), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n588), .B1(new_n294), .B2(new_n415), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n586), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n590), .A2(new_n282), .B1(new_n280), .B2(new_n325), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n591), .B1(new_n541), .B2(new_n325), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n457), .A2(new_n562), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n275), .A2(new_n457), .B1(new_n593), .B2(new_n308), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n411), .A2(new_n264), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n311), .A2(G1698), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n595), .B(new_n596), .C1(new_n250), .C2(new_n251), .ZN(new_n597));
  AND2_X1   g0397(.A1(new_n597), .A2(new_n517), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n594), .B1(new_n598), .B2(new_n308), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n498), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n593), .A2(new_n308), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n308), .A2(G274), .A3(new_n457), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n308), .B1(new_n597), .B2(new_n517), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n307), .ZN(new_n606));
  AND3_X1   g0406(.A1(new_n592), .A2(new_n600), .A3(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(G200), .B1(new_n603), .B2(new_n604), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n489), .A2(G87), .A3(new_n283), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n608), .A2(new_n591), .A3(KEYINPUT80), .A4(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n605), .A2(G190), .ZN(new_n611));
  AND2_X1   g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT80), .ZN(new_n613));
  INV_X1    g0413(.A(new_n608), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n591), .A2(new_n609), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n607), .B1(new_n612), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n582), .A2(new_n617), .ZN(new_n618));
  NOR4_X1   g0418(.A1(new_n455), .A2(new_n504), .A3(new_n575), .A4(new_n618), .ZN(G372));
  NOR2_X1   g0419(.A1(new_n303), .A2(new_n306), .ZN(new_n620));
  INV_X1    g0420(.A(new_n408), .ZN(new_n621));
  INV_X1    g0421(.A(new_n335), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n452), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n621), .B1(new_n623), .B2(new_n448), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT86), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n625), .B1(new_n384), .B2(new_n398), .ZN(new_n626));
  INV_X1    g0426(.A(new_n383), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT16), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n290), .B1(new_n568), .B2(new_n569), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n628), .B1(new_n629), .B2(new_n366), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n627), .B1(new_n630), .B2(new_n373), .ZN(new_n631));
  OAI21_X1  g0431(.A(KEYINPUT18), .B1(new_n631), .B2(new_n360), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n396), .A2(new_n385), .A3(new_n397), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n632), .A2(KEYINPUT86), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n626), .A2(new_n634), .ZN(new_n635));
  OR2_X1    g0435(.A1(new_n624), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n620), .B1(new_n636), .B2(new_n349), .ZN(new_n637));
  INV_X1    g0437(.A(new_n607), .ZN(new_n638));
  AOI22_X1  g0438(.A1(new_n608), .A2(KEYINPUT85), .B1(new_n605), .B2(G190), .ZN(new_n639));
  INV_X1    g0439(.A(new_n615), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n639), .B(new_n640), .C1(KEYINPUT85), .C2(new_n608), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n642), .A2(new_n566), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT26), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n607), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n566), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(new_n617), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(KEYINPUT26), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n501), .A2(new_n493), .ZN(new_n649));
  INV_X1    g0449(.A(new_n582), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n566), .A2(new_n574), .ZN(new_n652));
  INV_X1    g0452(.A(new_n642), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n652), .A2(new_n653), .A3(new_n544), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n645), .B(new_n648), .C1(new_n651), .C2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n637), .B1(new_n455), .B2(new_n656), .ZN(G369));
  OR3_X1    g0457(.A1(new_n486), .A2(KEYINPUT27), .A3(G20), .ZN(new_n658));
  OAI21_X1  g0458(.A(KEYINPUT27), .B1(new_n486), .B2(G20), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(G213), .A3(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(G343), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n492), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g0463(.A(new_n663), .B(KEYINPUT87), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n649), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n665), .B1(new_n504), .B2(new_n664), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n666), .A2(G330), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n662), .B1(new_n580), .B2(new_n581), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n650), .B1(new_n544), .B2(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n582), .A2(new_n662), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g0472(.A(new_n672), .B(KEYINPUT88), .ZN(new_n673));
  INV_X1    g0473(.A(new_n670), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n500), .B1(new_n494), .B2(new_n496), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n675), .A2(new_n662), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n671), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n673), .A2(new_n674), .A3(new_n677), .ZN(G399));
  INV_X1    g0478(.A(new_n212), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n679), .A2(G41), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n585), .A2(G116), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(G1), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n683), .B1(new_n203), .B2(new_n681), .ZN(new_n684));
  XOR2_X1   g0484(.A(new_n684), .B(KEYINPUT28), .Z(new_n685));
  NOR2_X1   g0485(.A1(new_n575), .A2(new_n618), .ZN(new_n686));
  INV_X1    g0486(.A(new_n662), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n686), .A2(new_n675), .A3(new_n503), .A4(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n528), .B1(new_n531), .B2(new_n308), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n599), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n474), .A2(new_n564), .A3(G179), .A4(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT30), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n532), .A2(new_n599), .A3(new_n307), .ZN(new_n694));
  OR3_X1    g0494(.A1(new_n474), .A2(new_n564), .A3(new_n694), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n476), .A2(new_n307), .A3(new_n462), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n696), .A2(KEYINPUT30), .A3(new_n564), .A4(new_n690), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n693), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(new_n662), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(KEYINPUT31), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT31), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n698), .A2(new_n701), .A3(new_n662), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n688), .A2(new_n703), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n704), .A2(G330), .ZN(new_n705));
  INV_X1    g0505(.A(new_n654), .ZN(new_n706));
  INV_X1    g0506(.A(new_n675), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n706), .B1(new_n707), .B2(new_n650), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n647), .A2(KEYINPUT26), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n638), .B1(new_n643), .B2(new_n644), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n662), .B1(new_n708), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(KEYINPUT29), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n655), .A2(new_n687), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT29), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n705), .B1(new_n713), .B2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n685), .B1(new_n718), .B2(new_n209), .ZN(new_n719));
  XOR2_X1   g0519(.A(new_n719), .B(KEYINPUT89), .Z(G364));
  NOR2_X1   g0520(.A1(new_n279), .A2(G20), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n209), .B1(new_n721), .B2(G45), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n680), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n667), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n725), .B1(G330), .B2(new_n666), .ZN(new_n726));
  NOR2_X1   g0526(.A1(G13), .A2(G33), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(new_n206), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n205), .B1(G20), .B2(new_n498), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n243), .A2(G45), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n679), .A2(new_n463), .ZN(new_n734));
  OAI211_X1 g0534(.A(new_n733), .B(new_n734), .C1(G45), .C2(new_n203), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n679), .A2(new_n330), .ZN(new_n736));
  AOI22_X1  g0536(.A1(new_n736), .A2(G355), .B1(new_n225), .B2(new_n679), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n732), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n730), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n400), .A2(new_n338), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n206), .A2(G179), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(G303), .ZN(new_n743));
  NAND2_X1  g0543(.A1(G20), .A2(G179), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(G190), .A2(G200), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(G311), .ZN(new_n748));
  OAI22_X1  g0548(.A1(new_n742), .A2(new_n743), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NOR3_X1   g0549(.A1(new_n400), .A2(G179), .A3(G200), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(new_n206), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  AOI211_X1 g0552(.A(new_n749), .B(new_n263), .C1(G294), .C2(new_n752), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n744), .A2(new_n400), .A3(G200), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(G322), .ZN(new_n756));
  XOR2_X1   g0556(.A(KEYINPUT33), .B(G317), .Z(new_n757));
  NOR2_X1   g0557(.A1(new_n338), .A2(G190), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(new_n745), .ZN(new_n759));
  OAI22_X1  g0559(.A1(new_n755), .A2(new_n756), .B1(new_n757), .B2(new_n759), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n760), .B(KEYINPUT90), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n741), .A2(new_n746), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(G329), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n740), .A2(new_n745), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n741), .A2(new_n758), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI22_X1  g0568(.A1(G326), .A2(new_n766), .B1(new_n768), .B2(G283), .ZN(new_n769));
  NAND4_X1  g0569(.A1(new_n753), .A2(new_n761), .A3(new_n764), .A4(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G159), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n762), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT32), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n752), .A2(G97), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n765), .A2(new_n223), .B1(new_n759), .B2(new_n290), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n767), .A2(new_n219), .B1(new_n747), .B2(new_n266), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n755), .A2(new_n217), .B1(new_n742), .B2(new_n510), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n330), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n773), .A2(new_n774), .A3(new_n777), .A4(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n739), .B1(new_n770), .B2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n724), .ZN(new_n782));
  NOR3_X1   g0582(.A1(new_n738), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n783), .B1(new_n666), .B2(new_n728), .ZN(new_n784));
  AND2_X1   g0584(.A1(new_n726), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(G396));
  NAND2_X1  g0586(.A1(new_n328), .A2(new_n662), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n335), .A2(new_n339), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(KEYINPUT94), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n622), .A2(new_n662), .ZN(new_n790));
  INV_X1    g0590(.A(KEYINPUT94), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n335), .A2(new_n339), .A3(new_n791), .A4(new_n787), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n789), .A2(new_n790), .A3(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(new_n727), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n730), .A2(new_n727), .ZN(new_n796));
  XOR2_X1   g0596(.A(new_n796), .B(KEYINPUT91), .Z(new_n797));
  OAI21_X1  g0597(.A(new_n724), .B1(new_n797), .B2(G77), .ZN(new_n798));
  INV_X1    g0598(.A(G294), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n755), .A2(new_n799), .B1(new_n747), .B2(new_n225), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n742), .A2(new_n219), .B1(new_n767), .B2(new_n510), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n765), .A2(new_n743), .B1(new_n762), .B2(new_n748), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(new_n263), .ZN(new_n804));
  INV_X1    g0604(.A(KEYINPUT92), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n759), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n758), .A2(new_n745), .A3(KEYINPUT92), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(G283), .ZN(new_n809));
  NAND4_X1  g0609(.A1(new_n802), .A2(new_n804), .A3(new_n809), .A4(new_n774), .ZN(new_n810));
  INV_X1    g0610(.A(G137), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n765), .A2(new_n811), .B1(new_n759), .B2(new_n295), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(KEYINPUT93), .ZN(new_n813));
  INV_X1    g0613(.A(G143), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n813), .B1(new_n814), .B2(new_n755), .C1(new_n771), .C2(new_n747), .ZN(new_n815));
  XOR2_X1   g0615(.A(new_n815), .B(KEYINPUT34), .Z(new_n816));
  AOI22_X1  g0616(.A1(G68), .A2(new_n768), .B1(new_n763), .B2(G132), .ZN(new_n817));
  INV_X1    g0617(.A(new_n742), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n375), .B1(new_n818), .B2(G50), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n817), .B(new_n819), .C1(new_n217), .C2(new_n751), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n810), .B1(new_n816), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n798), .B1(new_n821), .B2(new_n730), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n795), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n714), .A2(new_n794), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n789), .A2(new_n792), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n655), .A2(new_n687), .A3(new_n825), .ZN(new_n826));
  AND2_X1   g0626(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  OR2_X1    g0627(.A1(new_n827), .A2(new_n705), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n724), .B1(new_n828), .B2(KEYINPUT96), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(KEYINPUT96), .B2(new_n828), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n827), .A2(new_n705), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT95), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n823), .B1(new_n830), .B2(new_n832), .ZN(G384));
  INV_X1    g0633(.A(new_n552), .ZN(new_n834));
  OR2_X1    g0634(.A1(new_n834), .A2(KEYINPUT35), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(KEYINPUT35), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n835), .A2(G116), .A3(new_n207), .A4(new_n836), .ZN(new_n837));
  XOR2_X1   g0637(.A(new_n837), .B(KEYINPUT36), .Z(new_n838));
  OAI211_X1 g0638(.A(new_n204), .B(G77), .C1(new_n217), .C2(new_n290), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n223), .A2(G68), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n209), .B(G13), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n448), .A2(new_n662), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT38), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n290), .B1(new_n369), .B2(new_n370), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n628), .B1(new_n846), .B2(new_n366), .ZN(new_n847));
  AND3_X1   g0647(.A1(new_n847), .A2(new_n394), .A3(new_n282), .ZN(new_n848));
  OR2_X1    g0648(.A1(new_n848), .A2(new_n627), .ZN(new_n849));
  INV_X1    g0649(.A(new_n660), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n851), .B1(new_n399), .B2(new_n408), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n396), .A2(new_n397), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n396), .A2(new_n850), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT37), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n853), .A2(new_n854), .A3(new_n855), .A4(new_n404), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n848), .A2(new_n627), .B1(new_n397), .B2(new_n850), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n404), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(KEYINPUT37), .ZN(new_n859));
  AND2_X1   g0659(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n845), .B1(new_n852), .B2(new_n860), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n632), .A2(new_n633), .A3(new_n406), .A4(new_n407), .ZN(new_n862));
  INV_X1    g0662(.A(new_n851), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n856), .A2(new_n859), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n864), .A2(KEYINPUT38), .A3(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n861), .A2(KEYINPUT97), .A3(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT98), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT97), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n869), .B(new_n845), .C1(new_n852), .C2(new_n860), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n867), .A2(new_n868), .A3(KEYINPUT39), .A4(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n867), .A2(KEYINPUT39), .A3(new_n870), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(KEYINPUT98), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT99), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n866), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n864), .A2(KEYINPUT99), .A3(KEYINPUT38), .A4(new_n865), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n626), .A2(new_n634), .A3(new_n408), .ZN(new_n878));
  INV_X1    g0678(.A(new_n854), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n853), .A2(new_n854), .A3(new_n404), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(KEYINPUT37), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n856), .ZN(new_n883));
  AOI21_X1  g0683(.A(KEYINPUT38), .B1(new_n880), .B2(new_n883), .ZN(new_n884));
  NOR3_X1   g0684(.A1(new_n877), .A2(KEYINPUT39), .A3(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n871), .B1(new_n873), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(KEYINPUT100), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n878), .A2(new_n879), .B1(new_n856), .B2(new_n882), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n875), .B(new_n876), .C1(KEYINPUT38), .C2(new_n888), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n872), .B(KEYINPUT98), .C1(new_n889), .C2(KEYINPUT39), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT100), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n890), .A2(new_n891), .A3(new_n871), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n844), .B1(new_n887), .B2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n335), .A2(new_n662), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n826), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n447), .A2(new_n662), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n448), .A2(new_n452), .A3(new_n897), .ZN(new_n898));
  AND3_X1   g0698(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n447), .B(new_n662), .C1(new_n899), .C2(new_n431), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n896), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n903), .A2(new_n870), .A3(new_n867), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n635), .A2(new_n660), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n893), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n454), .A2(new_n713), .A3(new_n716), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n908), .A2(new_n637), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n907), .B(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT40), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n867), .A2(new_n870), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n704), .A2(new_n793), .A3(new_n901), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n911), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AND3_X1   g0714(.A1(new_n704), .A2(new_n793), .A3(new_n901), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n889), .A2(new_n915), .A3(KEYINPUT40), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n454), .A2(new_n704), .ZN(new_n918));
  OR2_X1    g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n917), .A2(new_n918), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n919), .A2(G330), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n910), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n209), .B2(new_n721), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n910), .A2(new_n921), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n842), .B1(new_n923), .B2(new_n924), .ZN(G367));
  NAND2_X1  g0725(.A1(new_n555), .A2(new_n662), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n565), .B1(G169), .B2(new_n564), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n928), .A2(KEYINPUT101), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n652), .A2(new_n926), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n928), .A2(KEYINPUT101), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n929), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n566), .B1(new_n933), .B2(new_n582), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n932), .A2(new_n671), .A3(new_n676), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n934), .A2(new_n687), .B1(KEYINPUT42), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(KEYINPUT42), .B2(new_n935), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n615), .A2(new_n662), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n653), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n638), .B2(new_n938), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(KEYINPUT43), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n937), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n940), .A2(KEYINPUT43), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n673), .A2(new_n933), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n942), .A2(new_n943), .ZN(new_n947));
  AND3_X1   g0747(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n946), .B1(new_n945), .B2(new_n947), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n680), .B(KEYINPUT41), .Z(new_n951));
  XNOR2_X1  g0751(.A(new_n671), .B(new_n676), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(new_n667), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n717), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT88), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n672), .B(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n677), .A2(new_n674), .A3(new_n932), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT45), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n957), .A2(new_n958), .ZN(new_n960));
  OR2_X1    g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n677), .A2(new_n674), .ZN(new_n962));
  AND3_X1   g0762(.A1(new_n962), .A2(KEYINPUT44), .A3(new_n933), .ZN(new_n963));
  AOI21_X1  g0763(.A(KEYINPUT44), .B1(new_n962), .B2(new_n933), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n956), .A2(new_n961), .A3(new_n965), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n960), .A2(new_n959), .B1(new_n963), .B2(new_n964), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n673), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n954), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT102), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n951), .B1(new_n970), .B2(new_n717), .ZN(new_n971));
  OAI211_X1 g0771(.A(KEYINPUT103), .B(new_n950), .C1(new_n971), .C2(new_n723), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT103), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n969), .A2(KEYINPUT102), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT102), .ZN(new_n975));
  AOI211_X1 g0775(.A(new_n975), .B(new_n954), .C1(new_n966), .C2(new_n968), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n717), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n951), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n723), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n950), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n973), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n972), .A2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n734), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n731), .B1(new_n212), .B2(new_n325), .C1(new_n983), .C2(new_n238), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n724), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT104), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n742), .A2(new_n225), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT46), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n988), .B1(G107), .B2(new_n752), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n375), .B1(new_n767), .B2(new_n415), .ZN(new_n990));
  INV_X1    g0790(.A(G317), .ZN(new_n991));
  INV_X1    g0791(.A(G283), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n762), .A2(new_n991), .B1(new_n747), .B2(new_n992), .ZN(new_n993));
  AOI211_X1 g0793(.A(new_n990), .B(new_n993), .C1(G294), .C2(new_n808), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n755), .A2(new_n743), .B1(new_n765), .B2(new_n748), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT105), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n989), .A2(new_n994), .A3(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n808), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n998), .A2(new_n771), .B1(new_n223), .B2(new_n747), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(KEYINPUT106), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n768), .A2(G77), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n1001), .B(new_n263), .C1(new_n811), .C2(new_n762), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(G68), .B2(new_n752), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n818), .A2(G58), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n766), .A2(G143), .B1(G150), .B2(new_n754), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n1000), .A2(new_n1003), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n999), .A2(KEYINPUT106), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n997), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT47), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n730), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n986), .B1(new_n1010), .B2(new_n1012), .C1(new_n940), .C2(new_n728), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1013), .B(KEYINPUT107), .Z(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n982), .A2(new_n1015), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n1016), .A2(KEYINPUT108), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(KEYINPUT108), .ZN(new_n1018));
  AND2_X1   g0818(.A1(new_n1017), .A2(new_n1018), .ZN(G387));
  OAI22_X1  g0819(.A1(new_n751), .A2(new_n992), .B1(new_n742), .B2(new_n799), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n754), .A2(G317), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1021), .B1(new_n747), .B2(new_n743), .C1(new_n756), .C2(new_n765), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(G311), .B2(new_n808), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1020), .B1(new_n1023), .B2(KEYINPUT48), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n1024), .B(KEYINPUT110), .Z(new_n1025));
  OR2_X1    g0825(.A1(new_n1023), .A2(KEYINPUT48), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT111), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1025), .A2(KEYINPUT111), .A3(new_n1026), .ZN(new_n1030));
  AND3_X1   g0830(.A1(new_n1029), .A2(KEYINPUT49), .A3(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(KEYINPUT49), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n463), .B1(new_n763), .B2(G326), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n225), .B2(new_n767), .ZN(new_n1034));
  OR3_X1    g0834(.A1(new_n1031), .A2(new_n1032), .A3(new_n1034), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n765), .A2(new_n771), .B1(new_n759), .B2(new_n293), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n375), .B(new_n1036), .C1(G97), .C2(new_n768), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n747), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(G150), .A2(new_n763), .B1(new_n1038), .B2(G68), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n818), .A2(G77), .B1(G50), .B2(new_n754), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n751), .A2(new_n325), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n1037), .A2(new_n1039), .A3(new_n1040), .A4(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n739), .B1(new_n1035), .B2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n671), .A2(new_n728), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n734), .B1(new_n235), .B2(new_n456), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n736), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1045), .B1(new_n682), .B2(new_n1046), .ZN(new_n1047));
  OR3_X1    g0847(.A1(new_n293), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1048));
  OAI21_X1  g0848(.A(KEYINPUT50), .B1(new_n293), .B2(G50), .ZN(new_n1049));
  AOI21_X1  g0849(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n1048), .A2(new_n682), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n1047), .A2(new_n1051), .B1(new_n219), .B2(new_n679), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n724), .B1(new_n1052), .B2(new_n732), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT109), .Z(new_n1054));
  NOR3_X1   g0854(.A1(new_n1043), .A2(new_n1044), .A3(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(new_n723), .B2(new_n953), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n953), .A2(new_n717), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n954), .A2(new_n680), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1056), .B1(new_n1057), .B2(new_n1058), .ZN(G393));
  INV_X1    g0859(.A(new_n954), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n966), .A2(new_n968), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n680), .B1(new_n1060), .B2(new_n1061), .C1(new_n974), .C2(new_n976), .ZN(new_n1062));
  AND2_X1   g0862(.A1(new_n734), .A2(new_n246), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n731), .B1(new_n212), .B2(new_n415), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n742), .A2(new_n290), .B1(new_n762), .B2(new_n814), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n375), .B(new_n1065), .C1(G87), .C2(new_n768), .ZN(new_n1066));
  XOR2_X1   g0866(.A(new_n1066), .B(KEYINPUT112), .Z(new_n1067));
  OAI22_X1  g0867(.A1(new_n755), .A2(new_n771), .B1(new_n765), .B2(new_n295), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT51), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n751), .A2(new_n266), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n293), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1070), .B1(new_n1071), .B2(new_n1038), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1069), .B(new_n1072), .C1(new_n223), .C2(new_n998), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n766), .A2(G317), .B1(G311), .B2(new_n754), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT52), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n767), .A2(new_n219), .B1(new_n747), .B2(new_n799), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n742), .A2(new_n992), .B1(new_n762), .B2(new_n756), .ZN(new_n1078));
  NOR4_X1   g0878(.A1(new_n1076), .A2(new_n263), .A3(new_n1077), .A4(new_n1078), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n808), .A2(G303), .B1(G116), .B2(new_n752), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT113), .Z(new_n1081));
  AOI22_X1  g0881(.A1(new_n1067), .A2(new_n1074), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n724), .B1(new_n1063), .B2(new_n1064), .C1(new_n1082), .C2(new_n739), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(new_n933), .B2(new_n729), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(new_n1061), .B2(new_n723), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1062), .A2(new_n1085), .ZN(G390));
  INV_X1    g0886(.A(KEYINPUT114), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n705), .A2(new_n793), .A3(new_n901), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n894), .B1(new_n712), .B2(new_n825), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n704), .A2(G330), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n902), .B1(new_n1090), .B2(new_n794), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1088), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1092));
  AND2_X1   g0892(.A1(new_n1088), .A2(new_n1091), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1087), .B(new_n1092), .C1(new_n1093), .C2(new_n896), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n454), .A2(new_n705), .ZN(new_n1095));
  AND3_X1   g0895(.A1(new_n908), .A2(new_n637), .A3(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1093), .A2(KEYINPUT114), .A3(new_n1089), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1094), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n844), .B1(new_n896), .B2(new_n902), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n887), .A2(new_n892), .A3(new_n1099), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n844), .B(new_n889), .C1(new_n1089), .C2(new_n902), .ZN(new_n1101));
  AND3_X1   g0901(.A1(new_n1100), .A2(new_n1088), .A3(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1088), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1098), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1088), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1100), .A2(new_n1088), .A3(new_n1101), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1098), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1107), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1104), .A2(new_n1110), .A3(new_n680), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(KEYINPUT54), .B(G143), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n752), .A2(G159), .B1(new_n1038), .B2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n998), .B2(new_n811), .ZN(new_n1115));
  XOR2_X1   g0915(.A(new_n1115), .B(KEYINPUT115), .Z(new_n1116));
  NOR2_X1   g0916(.A1(new_n742), .A2(new_n295), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT53), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n263), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(G50), .A2(new_n768), .B1(new_n763), .B2(G125), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n766), .A2(G128), .B1(G132), .B2(new_n754), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  AOI211_X1 g0922(.A(new_n1119), .B(new_n1122), .C1(new_n1118), .C2(new_n1117), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n808), .A2(G107), .B1(G97), .B2(new_n1038), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT116), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n765), .A2(new_n992), .B1(new_n767), .B2(new_n290), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n755), .A2(new_n225), .B1(new_n762), .B2(new_n799), .ZN(new_n1128));
  NOR4_X1   g0928(.A1(new_n1126), .A2(new_n1070), .A3(new_n1127), .A4(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n263), .B1(G87), .B2(new_n818), .ZN(new_n1130));
  OR2_X1    g0930(.A1(new_n1130), .A2(KEYINPUT117), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(KEYINPUT117), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n1131), .A2(new_n1132), .B1(new_n1125), .B2(new_n1124), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n1116), .A2(new_n1123), .B1(new_n1129), .B2(new_n1133), .ZN(new_n1134));
  OAI221_X1 g0934(.A(new_n724), .B1(new_n1071), .B2(new_n797), .C1(new_n1134), .C2(new_n739), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n892), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n891), .B1(new_n890), .B2(new_n871), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1135), .B1(new_n1138), .B2(new_n727), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1139), .B1(new_n1140), .B2(new_n723), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1111), .A2(new_n1141), .ZN(G378));
  NAND3_X1  g0942(.A1(new_n914), .A2(G330), .A3(new_n916), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n300), .A2(new_n660), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n349), .A2(new_n302), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1147), .B1(new_n349), .B2(new_n302), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1145), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1150), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1152), .A2(new_n1148), .A3(new_n1144), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1143), .A2(new_n1155), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1154), .A2(new_n914), .A3(G330), .A4(new_n916), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(KEYINPUT122), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n843), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n906), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1159), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT122), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1164), .B1(new_n893), .B2(new_n906), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1162), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(new_n723), .ZN(new_n1167));
  AOI211_X1 g0967(.A(G41), .B(new_n463), .C1(new_n818), .C2(G77), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n325), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(G58), .A2(new_n768), .B1(new_n1038), .B2(new_n1169), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1168), .B(new_n1170), .C1(new_n290), .C2(new_n751), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n755), .A2(new_n219), .B1(new_n762), .B2(new_n992), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n765), .A2(new_n225), .B1(new_n759), .B2(new_n415), .ZN(new_n1173));
  NOR3_X1   g0973(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  OR2_X1    g0974(.A1(new_n1174), .A2(KEYINPUT58), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(KEYINPUT58), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(G33), .A2(G41), .ZN(new_n1177));
  XOR2_X1   g0977(.A(new_n1177), .B(KEYINPUT118), .Z(new_n1178));
  OAI211_X1 g0978(.A(new_n1178), .B(new_n223), .C1(G41), .C2(new_n463), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1175), .A2(new_n1176), .A3(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(G132), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n1181), .A2(new_n759), .B1(new_n742), .B2(new_n1112), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n766), .A2(G125), .B1(G128), .B2(new_n754), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1183), .B1(new_n811), .B2(new_n747), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n1182), .B(new_n1184), .C1(G150), .C2(new_n752), .ZN(new_n1185));
  XOR2_X1   g0985(.A(new_n1185), .B(KEYINPUT59), .Z(new_n1186));
  OR2_X1    g0986(.A1(new_n1186), .A2(KEYINPUT119), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(G159), .A2(new_n768), .B1(new_n763), .B2(G124), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1178), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1190), .B(KEYINPUT120), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(new_n1186), .B2(KEYINPUT119), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1180), .B1(new_n1187), .B2(new_n1192), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1193), .A2(new_n739), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1194), .B(KEYINPUT121), .ZN(new_n1195));
  AOI211_X1 g0995(.A(new_n782), .B(new_n1195), .C1(new_n223), .C2(new_n796), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1155), .A2(new_n727), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1167), .A2(KEYINPUT123), .A3(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT123), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n722), .B1(new_n1162), .B2(new_n1165), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1198), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1200), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1199), .A2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT57), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1160), .A2(new_n1161), .A3(new_n1157), .A4(new_n1156), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1158), .B1(new_n893), .B2(new_n906), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1205), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  NOR3_X1   g1008(.A1(new_n1102), .A2(new_n1103), .A3(new_n1098), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1096), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1208), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(new_n680), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1110), .A2(new_n1096), .ZN(new_n1213));
  AOI21_X1  g1013(.A(KEYINPUT57), .B1(new_n1213), .B2(new_n1166), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1204), .B1(new_n1212), .B2(new_n1214), .ZN(G375));
  AOI21_X1  g1015(.A(new_n1096), .B1(new_n1094), .B2(new_n1097), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1217), .A2(new_n978), .A3(new_n1098), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1092), .A2(new_n1087), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n896), .B1(new_n1088), .B2(new_n1091), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1097), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n902), .A2(new_n727), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n724), .B1(new_n797), .B2(G68), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(G128), .A2(new_n763), .B1(new_n1038), .B2(G150), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n1225), .B1(new_n811), .B2(new_n755), .C1(new_n998), .C2(new_n1112), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(G132), .A2(new_n766), .B1(new_n818), .B2(G159), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n375), .B1(new_n768), .B2(G58), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n1227), .B(new_n1228), .C1(new_n223), .C2(new_n751), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n766), .A2(G294), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1041), .A2(new_n330), .A3(new_n1230), .A4(new_n1001), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n1038), .A2(G107), .B1(G283), .B2(new_n754), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(G97), .A2(new_n818), .B1(new_n763), .B2(G303), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1232), .B(new_n1233), .C1(new_n998), .C2(new_n225), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n1226), .A2(new_n1229), .B1(new_n1231), .B2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1224), .B1(new_n1235), .B2(new_n730), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n1222), .A2(new_n723), .B1(new_n1223), .B2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1218), .A2(new_n1237), .ZN(G381));
  NOR4_X1   g1038(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1239));
  INV_X1    g1039(.A(G378), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1239), .A2(new_n1240), .A3(new_n1237), .A4(new_n1218), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1242));
  XOR2_X1   g1042(.A(G375), .B(KEYINPUT124), .Z(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(G407));
  AND2_X1   g1044(.A1(new_n661), .A2(G213), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1243), .A2(new_n1240), .A3(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(G407), .A2(G213), .A3(new_n1246), .ZN(G409));
  OAI211_X1 g1047(.A(new_n1204), .B(G378), .C1(new_n1212), .C2(new_n1214), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1213), .A2(new_n978), .A3(new_n1166), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1202), .B1(new_n1250), .B2(new_n723), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1249), .A2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(new_n1240), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1245), .B1(new_n1248), .B2(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1216), .B1(KEYINPUT60), .B2(new_n1098), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1221), .A2(new_n1210), .A3(KEYINPUT60), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(new_n680), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1237), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(G384), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  OAI211_X1 g1060(.A(G384), .B(new_n1237), .C1(new_n1255), .C2(new_n1257), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1260), .A2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1254), .A2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT63), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1267), .A2(KEYINPUT125), .A3(new_n1261), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1245), .A2(G2897), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1268), .A2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT125), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1272), .B1(new_n1260), .B2(new_n1262), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1271), .A2(new_n1273), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1272), .B(new_n1270), .C1(new_n1260), .C2(new_n1262), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  OR2_X1    g1076(.A1(new_n1254), .A2(new_n1276), .ZN(new_n1277));
  XNOR2_X1  g1077(.A(G393), .B(new_n785), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n1062), .B(new_n1085), .C1(new_n1278), .C2(KEYINPUT108), .ZN(new_n1279));
  INV_X1    g1079(.A(G390), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1279), .B1(new_n1280), .B2(new_n1278), .ZN(new_n1281));
  AND3_X1   g1081(.A1(new_n982), .A2(new_n1281), .A3(new_n1015), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1281), .B1(new_n982), .B2(new_n1015), .ZN(new_n1283));
  NOR3_X1   g1083(.A1(new_n1282), .A2(new_n1283), .A3(KEYINPUT61), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1254), .A2(KEYINPUT63), .A3(new_n1263), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1266), .A2(new_n1277), .A3(new_n1284), .A4(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT62), .ZN(new_n1287));
  AND3_X1   g1087(.A1(new_n1254), .A2(new_n1287), .A3(new_n1263), .ZN(new_n1288));
  XOR2_X1   g1088(.A(KEYINPUT126), .B(KEYINPUT61), .Z(new_n1289));
  OAI21_X1  g1089(.A(new_n1289), .B1(new_n1254), .B2(new_n1276), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1287), .B1(new_n1254), .B2(new_n1263), .ZN(new_n1291));
  NOR3_X1   g1091(.A1(new_n1288), .A2(new_n1290), .A3(new_n1291), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1286), .B1(new_n1292), .B2(new_n1293), .ZN(G405));
  INV_X1    g1094(.A(KEYINPUT127), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1263), .A2(new_n1295), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1296), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1281), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1016), .A2(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n982), .A2(new_n1281), .A3(new_n1015), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1296), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1299), .A2(new_n1300), .A3(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1297), .A2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1263), .A2(new_n1295), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1248), .A2(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1305), .B1(new_n1240), .B2(G375), .ZN(new_n1306));
  XNOR2_X1  g1106(.A(new_n1303), .B(new_n1306), .ZN(G402));
endmodule


