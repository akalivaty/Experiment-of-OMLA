//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 1 0 1 0 1 1 1 1 1 1 1 1 0 1 1 0 1 1 0 0 0 0 0 1 1 1 0 1 0 1 1 1 0 0 0 1 0 1 1 1 1 1 1 1 0 0 1 0 0 1 0 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:51 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n882, new_n883, new_n884,
    new_n885, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964;
  INV_X1    g000(.A(G953), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G227), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(G140), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT77), .B(G110), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT12), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT11), .ZN(new_n194));
  INV_X1    g008(.A(G134), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n194), .B1(new_n195), .B2(G137), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(G137), .ZN(new_n197));
  INV_X1    g011(.A(G137), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n198), .A2(KEYINPUT11), .A3(G134), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n196), .A2(new_n197), .A3(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G131), .ZN(new_n201));
  INV_X1    g015(.A(G131), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n196), .A2(new_n199), .A3(new_n202), .A4(new_n197), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  XNOR2_X1  g019(.A(G143), .B(G146), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT1), .ZN(new_n207));
  AND3_X1   g021(.A1(new_n206), .A2(new_n207), .A3(G128), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G143), .ZN(new_n210));
  INV_X1    g024(.A(G143), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G146), .ZN(new_n212));
  AOI21_X1  g026(.A(G128), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  NOR3_X1   g027(.A1(new_n207), .A2(new_n209), .A3(G143), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT67), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n209), .A2(G143), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(KEYINPUT1), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT67), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n217), .B(new_n218), .C1(new_n206), .C2(G128), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n208), .B1(new_n215), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT78), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n222), .A2(G107), .ZN(new_n223));
  INV_X1    g037(.A(G107), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n224), .A2(KEYINPUT78), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n221), .B(G104), .C1(new_n223), .C2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G101), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n224), .A2(G104), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n224), .A2(G104), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n228), .B1(KEYINPUT3), .B2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n226), .A2(new_n227), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n224), .A2(KEYINPUT78), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n222), .A2(G107), .ZN(new_n233));
  INV_X1    g047(.A(G104), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(new_n229), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G101), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n231), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n220), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n206), .A2(new_n207), .A3(G128), .ZN(new_n240));
  INV_X1    g054(.A(G128), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n211), .A2(G146), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n241), .B1(new_n242), .B2(new_n216), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n240), .A2(new_n243), .A3(new_n217), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n244), .A2(new_n231), .A3(new_n237), .ZN(new_n245));
  AOI211_X1 g059(.A(new_n193), .B(new_n205), .C1(new_n239), .C2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT82), .ZN(new_n247));
  AND3_X1   g061(.A1(new_n239), .A2(KEYINPUT81), .A3(new_n245), .ZN(new_n248));
  AOI21_X1  g062(.A(KEYINPUT81), .B1(new_n239), .B2(new_n245), .ZN(new_n249));
  NOR3_X1   g063(.A1(new_n248), .A2(new_n249), .A3(new_n205), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n247), .B1(new_n250), .B2(KEYINPUT12), .ZN(new_n251));
  INV_X1    g065(.A(new_n249), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n239), .A2(KEYINPUT81), .A3(new_n245), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n252), .A2(new_n204), .A3(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n254), .A2(KEYINPUT82), .A3(new_n193), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n246), .B1(new_n251), .B2(new_n255), .ZN(new_n256));
  XNOR2_X1  g070(.A(KEYINPUT78), .B(G107), .ZN(new_n257));
  NOR3_X1   g071(.A1(new_n257), .A2(KEYINPUT3), .A3(new_n234), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n229), .A2(KEYINPUT3), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n259), .B1(G104), .B2(new_n224), .ZN(new_n260));
  OAI21_X1  g074(.A(G101), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n261), .A2(KEYINPUT4), .A3(new_n231), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT0), .B(G128), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT64), .ZN(new_n264));
  OR3_X1    g078(.A1(new_n206), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n206), .A2(KEYINPUT0), .A3(G128), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n264), .B1(new_n206), .B2(new_n263), .ZN(new_n267));
  AND3_X1   g081(.A1(new_n265), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT4), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n269), .B(G101), .C1(new_n258), .C2(new_n260), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n262), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n218), .B1(new_n243), .B2(new_n217), .ZN(new_n272));
  NOR3_X1   g086(.A1(new_n213), .A2(KEYINPUT67), .A3(new_n214), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n240), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n231), .A2(new_n237), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n274), .A2(new_n275), .A3(KEYINPUT10), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT80), .ZN(new_n277));
  XOR2_X1   g091(.A(KEYINPUT79), .B(KEYINPUT10), .Z(new_n278));
  AND3_X1   g092(.A1(new_n245), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n277), .B1(new_n245), .B2(new_n278), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n271), .B(new_n276), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n281), .A2(new_n204), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n192), .B1(new_n256), .B2(new_n282), .ZN(new_n283));
  OR2_X1    g097(.A1(new_n281), .A2(new_n204), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n191), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(KEYINPUT83), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n281), .A2(new_n204), .ZN(new_n287));
  OR3_X1    g101(.A1(new_n282), .A2(KEYINPUT83), .A3(new_n192), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n283), .A2(new_n289), .A3(G469), .ZN(new_n290));
  INV_X1    g104(.A(G469), .ZN(new_n291));
  XNOR2_X1  g105(.A(KEYINPUT72), .B(G902), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n251), .A2(new_n255), .ZN(new_n294));
  INV_X1    g108(.A(new_n246), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n285), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n191), .B1(new_n284), .B2(new_n287), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n291), .B(new_n293), .C1(new_n296), .C2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(G469), .A2(G902), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n290), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G221), .ZN(new_n301));
  XOR2_X1   g115(.A(KEYINPUT9), .B(G234), .Z(new_n302));
  INV_X1    g116(.A(G902), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  AND2_X1   g119(.A1(new_n300), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(G214), .B1(G237), .B2(G902), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n265), .A2(new_n266), .A3(new_n267), .ZN(new_n309));
  XNOR2_X1  g123(.A(KEYINPUT74), .B(G125), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n311), .B1(new_n274), .B2(new_n310), .ZN(new_n312));
  INV_X1    g126(.A(G224), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n313), .A2(G953), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n312), .B(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT6), .ZN(new_n316));
  NOR2_X1   g130(.A1(KEYINPUT2), .A2(G113), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n317), .B(KEYINPUT69), .ZN(new_n318));
  NAND2_X1  g132(.A1(KEYINPUT2), .A2(G113), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n319), .B(KEYINPUT70), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g135(.A(G116), .B(G119), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n318), .A2(new_n322), .A3(new_n320), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n262), .A2(new_n270), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT85), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n322), .A2(KEYINPUT5), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT5), .ZN(new_n330));
  INV_X1    g144(.A(G119), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n330), .A2(new_n331), .A3(G116), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT84), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n330), .A2(new_n331), .A3(KEYINPUT84), .A4(G116), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n329), .A2(G113), .A3(new_n334), .A4(new_n335), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n275), .A2(new_n328), .A3(new_n325), .A4(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n325), .ZN(new_n338));
  OAI21_X1  g152(.A(KEYINPUT85), .B1(new_n338), .B2(new_n238), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n327), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  XNOR2_X1  g154(.A(G110), .B(G122), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n341), .B(KEYINPUT86), .ZN(new_n342));
  XOR2_X1   g156(.A(new_n342), .B(KEYINPUT87), .Z(new_n343));
  NAND2_X1  g157(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n327), .A2(new_n337), .A3(new_n342), .A4(new_n339), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n316), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(KEYINPUT6), .B1(new_n340), .B2(new_n343), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n315), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n338), .B(new_n238), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n342), .B(KEYINPUT8), .ZN(new_n350));
  AOI22_X1  g164(.A1(new_n349), .A2(new_n350), .B1(new_n312), .B2(new_n314), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT7), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT88), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n352), .B1(new_n314), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n354), .B1(new_n353), .B2(new_n314), .ZN(new_n355));
  OR2_X1    g169(.A1(new_n312), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n312), .A2(new_n352), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n351), .A2(new_n356), .A3(new_n357), .A4(new_n345), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n348), .A2(new_n303), .A3(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(G210), .B1(G237), .B2(G902), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n348), .A2(new_n303), .A3(new_n360), .A4(new_n358), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n308), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(KEYINPUT96), .B(G952), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n365), .A2(G953), .ZN(new_n366));
  NAND2_X1  g180(.A1(G234), .A2(G237), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n292), .A2(G953), .A3(new_n367), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  XOR2_X1   g185(.A(KEYINPUT21), .B(G898), .Z(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n369), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n364), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(G116), .ZN(new_n378));
  OAI21_X1  g192(.A(KEYINPUT94), .B1(new_n378), .B2(G122), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT94), .ZN(new_n380));
  INV_X1    g194(.A(G122), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n381), .A3(G116), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n378), .A2(G122), .ZN(new_n384));
  AND2_X1   g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n257), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  XNOR2_X1  g201(.A(G128), .B(G143), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n388), .B(new_n195), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT95), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n384), .A2(KEYINPUT14), .ZN(new_n391));
  AND3_X1   g205(.A1(new_n383), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n390), .B1(new_n383), .B2(new_n391), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n384), .A2(KEYINPUT14), .ZN(new_n394));
  NOR3_X1   g208(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n387), .B(new_n389), .C1(new_n395), .C2(new_n224), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n388), .A2(KEYINPUT13), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n211), .A2(G128), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n397), .B(G134), .C1(KEYINPUT13), .C2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n388), .A2(new_n195), .ZN(new_n400));
  INV_X1    g214(.A(new_n387), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n385), .A2(new_n386), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n399), .B(new_n400), .C1(new_n401), .C2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n396), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n302), .A2(G217), .A3(new_n187), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n405), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n396), .A2(new_n403), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n292), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(G478), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n410), .A2(KEYINPUT15), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n409), .B(new_n411), .ZN(new_n412));
  NOR2_X1   g226(.A1(G125), .A2(G140), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n413), .B1(new_n310), .B2(G140), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(G146), .ZN(new_n415));
  XOR2_X1   g229(.A(G125), .B(G140), .Z(new_n416));
  OR2_X1    g230(.A1(new_n416), .A2(G146), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g232(.A1(G237), .A2(G953), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n419), .A2(G143), .A3(G214), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(G143), .B1(new_n419), .B2(G214), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT89), .ZN(new_n424));
  AOI22_X1  g238(.A1(new_n423), .A2(new_n424), .B1(KEYINPUT18), .B2(G131), .ZN(new_n425));
  NAND2_X1  g239(.A1(KEYINPUT18), .A2(G131), .ZN(new_n426));
  NOR4_X1   g240(.A1(new_n421), .A2(new_n422), .A3(KEYINPUT89), .A4(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n418), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n310), .A2(G140), .ZN(new_n429));
  INV_X1    g243(.A(new_n413), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n429), .A2(KEYINPUT19), .A3(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT90), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n432), .B1(new_n416), .B2(KEYINPUT19), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n414), .A2(new_n432), .A3(KEYINPUT19), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n434), .A2(new_n209), .A3(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(G131), .B1(new_n421), .B2(new_n422), .ZN(new_n437));
  INV_X1    g251(.A(new_n422), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(new_n202), .A3(new_n420), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT16), .ZN(new_n441));
  INV_X1    g255(.A(G140), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n310), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  OAI211_X1 g257(.A(G146), .B(new_n443), .C1(new_n414), .C2(new_n441), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n440), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n428), .B1(new_n436), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(KEYINPUT91), .ZN(new_n447));
  XNOR2_X1  g261(.A(G113), .B(G122), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n448), .B(new_n234), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT91), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n428), .B(new_n451), .C1(new_n436), .C2(new_n445), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n447), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n443), .B1(new_n414), .B2(new_n441), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n209), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n444), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT92), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT17), .ZN(new_n459));
  OR2_X1    g273(.A1(new_n437), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n455), .A2(KEYINPUT92), .A3(new_n444), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n437), .A2(new_n439), .A3(new_n459), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n458), .A2(new_n460), .A3(new_n461), .A4(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n463), .A2(new_n449), .A3(new_n428), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n453), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(G475), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n465), .A2(new_n466), .A3(new_n303), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT20), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n464), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n449), .B1(new_n463), .B2(new_n428), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n303), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(G475), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n465), .A2(KEYINPUT20), .A3(new_n466), .A4(new_n303), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n469), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT93), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n469), .A2(new_n473), .A3(KEYINPUT93), .A4(new_n474), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AND3_X1   g293(.A1(new_n377), .A2(new_n412), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n241), .A2(G119), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT23), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n331), .A2(G128), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n241), .A2(KEYINPUT23), .A3(G119), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(G110), .ZN(new_n487));
  XNOR2_X1  g301(.A(KEYINPUT24), .B(G110), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n488), .B(KEYINPUT73), .ZN(new_n489));
  AND2_X1   g303(.A1(new_n484), .A2(new_n481), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n456), .A2(new_n487), .A3(new_n491), .ZN(new_n492));
  OAI22_X1  g306(.A1(new_n489), .A2(new_n490), .B1(G110), .B2(new_n486), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n493), .A2(new_n444), .A3(new_n417), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT75), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n492), .A2(KEYINPUT75), .A3(new_n494), .ZN(new_n498));
  XNOR2_X1  g312(.A(KEYINPUT22), .B(G137), .ZN(new_n499));
  AND3_X1   g313(.A1(new_n187), .A2(G221), .A3(G234), .ZN(new_n500));
  XOR2_X1   g314(.A(new_n499), .B(new_n500), .Z(new_n501));
  NAND3_X1  g315(.A1(new_n497), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n501), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n492), .A2(KEYINPUT75), .A3(new_n494), .A4(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n293), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(KEYINPUT25), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT25), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n505), .A2(new_n508), .A3(new_n293), .ZN(new_n509));
  AND2_X1   g323(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(G217), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n511), .B1(new_n293), .B2(G234), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n512), .A2(G902), .ZN(new_n513));
  AOI22_X1  g327(.A1(new_n510), .A2(new_n512), .B1(new_n513), .B2(new_n505), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n309), .A2(new_n205), .ZN(new_n516));
  OAI21_X1  g330(.A(KEYINPUT65), .B1(new_n195), .B2(G137), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT65), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n518), .A2(new_n198), .A3(G134), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n517), .A2(new_n519), .A3(new_n197), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n520), .A2(KEYINPUT66), .A3(G131), .ZN(new_n521));
  AOI22_X1  g335(.A1(KEYINPUT66), .A2(new_n203), .B1(new_n520), .B2(G131), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n274), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT68), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n215), .A2(new_n219), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n522), .B1(new_n527), .B2(new_n240), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n528), .A2(KEYINPUT68), .A3(new_n521), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n516), .B1(new_n526), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n326), .ZN(new_n531));
  OAI21_X1  g345(.A(KEYINPUT71), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n268), .A2(new_n204), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n524), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n534), .A2(new_n326), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(KEYINPUT68), .B1(new_n528), .B2(new_n521), .ZN(new_n537));
  INV_X1    g351(.A(new_n521), .ZN(new_n538));
  NOR4_X1   g352(.A1(new_n220), .A2(new_n522), .A3(new_n538), .A4(new_n525), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n533), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT71), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n540), .A2(new_n541), .A3(new_n326), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n532), .A2(new_n536), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(KEYINPUT28), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n535), .A2(KEYINPUT28), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n419), .A2(G210), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n548), .B(new_n227), .ZN(new_n549));
  XNOR2_X1  g363(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n550));
  XOR2_X1   g364(.A(new_n549), .B(new_n550), .Z(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n516), .B1(new_n521), .B2(new_n528), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(KEYINPUT30), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n326), .B(new_n554), .C1(new_n530), .C2(KEYINPUT30), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n555), .A2(new_n536), .A3(new_n551), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT31), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n555), .A2(KEYINPUT31), .A3(new_n536), .A4(new_n551), .ZN(new_n559));
  AOI22_X1  g373(.A1(new_n547), .A2(new_n552), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NOR2_X1   g374(.A1(G472), .A2(G902), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  OAI21_X1  g376(.A(KEYINPUT32), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT28), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n540), .A2(new_n326), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n535), .B1(new_n565), .B2(KEYINPUT71), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n564), .B1(new_n566), .B2(new_n542), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n552), .B1(new_n567), .B2(new_n545), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n558), .A2(new_n559), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT32), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n570), .A2(new_n571), .A3(new_n561), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n563), .A2(new_n572), .ZN(new_n573));
  AOI211_X1 g387(.A(new_n545), .B(new_n552), .C1(new_n543), .C2(KEYINPUT28), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT29), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT30), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n534), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n577), .B1(new_n576), .B2(new_n540), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n535), .B1(new_n578), .B2(new_n326), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n575), .B1(new_n579), .B2(new_n551), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n293), .B1(new_n574), .B2(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n534), .B(new_n326), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(KEYINPUT28), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(new_n546), .ZN(new_n584));
  NOR3_X1   g398(.A1(new_n584), .A2(new_n575), .A3(new_n552), .ZN(new_n585));
  OAI21_X1  g399(.A(G472), .B1(new_n581), .B2(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n515), .B1(new_n573), .B2(new_n586), .ZN(new_n587));
  AND2_X1   g401(.A1(new_n587), .A2(KEYINPUT76), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n587), .A2(KEYINPUT76), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n306), .B(new_n480), .C1(new_n588), .C2(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(G101), .ZN(G3));
  NAND2_X1  g405(.A1(new_n570), .A2(new_n293), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT97), .ZN(new_n593));
  OAI21_X1  g407(.A(G472), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(KEYINPUT97), .B1(new_n570), .B2(new_n293), .ZN(new_n595));
  OAI22_X1  g409(.A1(new_n594), .A2(new_n595), .B1(new_n560), .B2(new_n562), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n597), .A2(new_n306), .A3(new_n514), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(KEYINPUT98), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n406), .A2(new_n408), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(KEYINPUT33), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT33), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n406), .A2(new_n602), .A3(new_n408), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n604), .A2(G478), .A3(new_n293), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT100), .ZN(new_n606));
  XNOR2_X1  g420(.A(KEYINPUT99), .B(G478), .ZN(new_n607));
  OAI211_X1 g421(.A(new_n605), .B(new_n606), .C1(new_n409), .C2(new_n607), .ZN(new_n608));
  AOI211_X1 g422(.A(new_n410), .B(new_n292), .C1(new_n601), .C2(new_n603), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n409), .A2(new_n607), .ZN(new_n610));
  OAI21_X1  g424(.A(KEYINPUT100), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n612), .A2(new_n477), .A3(new_n478), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n613), .A2(new_n376), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n599), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(new_n234), .ZN(new_n616));
  XNOR2_X1  g430(.A(KEYINPUT101), .B(KEYINPUT34), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G6));
  NOR3_X1   g432(.A1(new_n376), .A2(new_n412), .A3(new_n475), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n599), .A2(new_n619), .ZN(new_n620));
  XOR2_X1   g434(.A(KEYINPUT35), .B(G107), .Z(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G9));
  NAND3_X1  g436(.A1(new_n507), .A2(new_n512), .A3(new_n509), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n503), .A2(KEYINPUT36), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n495), .B(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(new_n513), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  AND4_X1   g441(.A1(new_n412), .A2(new_n479), .A3(new_n375), .A4(new_n627), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n597), .A2(new_n306), .A3(new_n364), .A4(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT37), .B(G110), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G12));
  AOI21_X1  g445(.A(new_n571), .B1(new_n570), .B2(new_n561), .ZN(new_n632));
  AOI211_X1 g446(.A(KEYINPUT32), .B(new_n562), .C1(new_n568), .C2(new_n569), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n586), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  AND3_X1   g448(.A1(new_n300), .A2(new_n305), .A3(new_n627), .ZN(new_n635));
  INV_X1    g449(.A(G900), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n371), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n368), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n475), .A2(new_n412), .A3(new_n639), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n634), .A2(new_n635), .A3(new_n364), .A4(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT102), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n364), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n644), .B1(new_n573), .B2(new_n586), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n645), .A2(KEYINPUT102), .A3(new_n640), .A4(new_n635), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G128), .ZN(G30));
  NAND2_X1  g462(.A1(new_n582), .A2(new_n552), .ZN(new_n649));
  OR2_X1    g463(.A1(new_n649), .A2(KEYINPUT103), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(KEYINPUT103), .ZN(new_n651));
  AND3_X1   g465(.A1(new_n650), .A2(new_n556), .A3(new_n651), .ZN(new_n652));
  OAI21_X1  g466(.A(G472), .B1(new_n652), .B2(G902), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n573), .A2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n655), .A2(new_n627), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n362), .A2(new_n363), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(KEYINPUT38), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NOR4_X1   g473(.A1(new_n659), .A2(new_n412), .A3(new_n479), .A4(new_n308), .ZN(new_n660));
  XOR2_X1   g474(.A(new_n638), .B(KEYINPUT39), .Z(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n306), .A2(new_n662), .ZN(new_n663));
  OR2_X1    g477(.A1(new_n663), .A2(KEYINPUT40), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(KEYINPUT40), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n656), .A2(new_n660), .A3(new_n664), .A4(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G143), .ZN(G45));
  NAND4_X1  g481(.A1(new_n612), .A2(new_n477), .A3(new_n478), .A4(new_n638), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n634), .A2(new_n635), .A3(new_n669), .A4(new_n364), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G146), .ZN(G48));
  NOR2_X1   g485(.A1(new_n296), .A2(new_n297), .ZN(new_n672));
  OAI21_X1  g486(.A(G469), .B1(new_n672), .B2(new_n292), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n673), .A2(new_n305), .A3(new_n298), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n587), .A2(new_n614), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(KEYINPUT41), .B(G113), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G15));
  NAND3_X1  g492(.A1(new_n587), .A2(new_n619), .A3(new_n675), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G116), .ZN(G18));
  NAND4_X1  g494(.A1(new_n628), .A2(new_n634), .A3(new_n364), .A4(new_n675), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT104), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n645), .A2(KEYINPUT104), .A3(new_n628), .A4(new_n675), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G119), .ZN(G21));
  NOR3_X1   g500(.A1(new_n674), .A2(new_n479), .A3(new_n412), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n584), .A2(new_n552), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n562), .B1(new_n569), .B2(new_n688), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n689), .B1(new_n592), .B2(G472), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n687), .A2(new_n514), .A3(new_n377), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G122), .ZN(G24));
  NOR2_X1   g506(.A1(new_n668), .A2(new_n674), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n693), .A2(new_n364), .A3(new_n627), .A4(new_n690), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G125), .ZN(G27));
  NAND3_X1  g509(.A1(new_n362), .A2(new_n307), .A3(new_n363), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT106), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n362), .A2(KEYINPUT106), .A3(new_n307), .A4(new_n363), .ZN(new_n699));
  AND2_X1   g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n299), .B(KEYINPUT105), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n290), .A2(new_n298), .A3(new_n701), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n702), .A2(new_n305), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n700), .A2(new_n703), .A3(KEYINPUT107), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n698), .A2(new_n702), .A3(new_n305), .A4(new_n699), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT107), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n668), .B1(new_n704), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n587), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT42), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n708), .A2(KEYINPUT42), .A3(new_n587), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G131), .ZN(G33));
  XNOR2_X1  g528(.A(new_n705), .B(KEYINPUT107), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n587), .A2(new_n640), .ZN(new_n716));
  OAI21_X1  g530(.A(KEYINPUT108), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n704), .A2(new_n707), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT108), .ZN(new_n719));
  AND3_X1   g533(.A1(new_n634), .A2(new_n514), .A3(new_n640), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n718), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n717), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G134), .ZN(G36));
  NAND2_X1  g537(.A1(new_n479), .A2(new_n612), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT43), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n479), .A2(KEYINPUT43), .A3(new_n612), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n728), .A2(new_n596), .A3(new_n627), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT44), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(KEYINPUT110), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT110), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n729), .A2(new_n733), .A3(new_n730), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(new_n298), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT109), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n283), .A2(new_n289), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n737), .B(G469), .C1(new_n738), .C2(KEYINPUT45), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(KEYINPUT45), .ZN(new_n740));
  AOI21_X1  g554(.A(KEYINPUT45), .B1(new_n283), .B2(new_n289), .ZN(new_n741));
  OAI21_X1  g555(.A(KEYINPUT109), .B1(new_n741), .B2(new_n291), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n739), .A2(new_n740), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n701), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT46), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n736), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n743), .A2(KEYINPUT46), .A3(new_n701), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n304), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n729), .A2(new_n730), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n698), .A2(new_n699), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n735), .A2(new_n662), .A3(new_n748), .A4(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G137), .ZN(G39));
  NOR4_X1   g567(.A1(new_n634), .A2(new_n750), .A3(new_n514), .A4(new_n668), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n748), .A2(KEYINPUT47), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT47), .ZN(new_n756));
  AOI211_X1 g570(.A(new_n756), .B(new_n304), .C1(new_n746), .C2(new_n747), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n754), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G140), .ZN(G42));
  AND2_X1   g573(.A1(new_n726), .A2(new_n727), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n690), .A2(new_n514), .A3(new_n369), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n748), .B(KEYINPUT47), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n673), .A2(new_n298), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n764), .A2(new_n305), .ZN(new_n765));
  OAI211_X1 g579(.A(new_n700), .B(new_n762), .C1(new_n763), .C2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT51), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n760), .A2(new_n674), .A3(new_n761), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n768), .A2(new_n308), .A3(new_n659), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT50), .ZN(new_n770));
  OR2_X1    g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n769), .A2(new_n770), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n767), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n750), .A2(new_n674), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n774), .A2(KEYINPUT114), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(KEYINPUT114), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n775), .A2(new_n369), .A3(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(new_n612), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n479), .ZN(new_n779));
  NOR4_X1   g593(.A1(new_n777), .A2(new_n515), .A3(new_n654), .A4(new_n779), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n775), .A2(new_n369), .A3(new_n728), .A4(new_n776), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n690), .A2(new_n627), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n782), .A2(KEYINPUT115), .A3(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT115), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n786), .B1(new_n781), .B2(new_n783), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n780), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n788), .A2(KEYINPUT116), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT116), .ZN(new_n790));
  AOI211_X1 g604(.A(new_n790), .B(new_n780), .C1(new_n787), .C2(new_n785), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n766), .B(new_n773), .C1(new_n789), .C2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n771), .A2(new_n772), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n766), .A2(new_n793), .A3(new_n788), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n767), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n782), .A2(new_n587), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n796), .A2(KEYINPUT48), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(KEYINPUT48), .ZN(new_n798));
  OR4_X1    g612(.A1(new_n515), .A2(new_n777), .A3(new_n613), .A4(new_n654), .ZN(new_n799));
  AND4_X1   g613(.A1(new_n366), .A2(new_n797), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n792), .A2(new_n795), .A3(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT53), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n694), .A2(new_n670), .ZN(new_n803));
  INV_X1    g617(.A(new_n627), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n804), .A2(new_n702), .A3(new_n305), .A4(new_n638), .ZN(new_n805));
  OR2_X1    g619(.A1(new_n805), .A2(KEYINPUT112), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(KEYINPUT112), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n644), .A2(new_n479), .A3(new_n412), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n806), .A2(new_n654), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n647), .A2(new_n803), .A3(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT52), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n647), .A2(new_n803), .A3(KEYINPUT52), .A4(new_n809), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  MUX2_X1   g628(.A(new_n778), .B(new_n412), .S(new_n479), .Z(new_n815));
  NOR2_X1   g629(.A1(new_n815), .A2(new_n376), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n816), .A2(new_n306), .A3(new_n514), .A4(new_n597), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n590), .A2(new_n817), .A3(new_n629), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n475), .A2(new_n639), .ZN(new_n820));
  AND4_X1   g634(.A1(new_n634), .A2(new_n700), .A3(new_n412), .A4(new_n820), .ZN(new_n821));
  AOI22_X1  g635(.A1(new_n708), .A2(new_n784), .B1(new_n821), .B2(new_n635), .ZN(new_n822));
  INV_X1    g636(.A(new_n721), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n719), .B1(new_n718), .B2(new_n720), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n822), .B(KEYINPUT111), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(KEYINPUT111), .B1(new_n722), .B2(new_n822), .ZN(new_n827));
  OAI211_X1 g641(.A(new_n814), .B(new_n819), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(new_n713), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n676), .A2(new_n691), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n685), .A2(new_n830), .A3(new_n679), .ZN(new_n831));
  OR2_X1    g645(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n802), .B1(new_n828), .B2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT54), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n831), .A2(KEYINPUT113), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT113), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n685), .A2(new_n830), .A3(new_n836), .A4(new_n679), .ZN(new_n837));
  AND4_X1   g651(.A1(KEYINPUT53), .A2(new_n835), .A3(new_n713), .A4(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n722), .A2(new_n822), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT111), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n818), .B1(new_n841), .B2(new_n825), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n838), .A2(new_n842), .A3(new_n814), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n833), .A2(new_n834), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n768), .A2(new_n364), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n829), .A2(new_n831), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n842), .A2(KEYINPUT53), .A3(new_n846), .A4(new_n814), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n833), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT54), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n801), .A2(new_n844), .A3(new_n845), .A4(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n850), .B1(G952), .B2(G953), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n764), .B(KEYINPUT49), .ZN(new_n852));
  NOR4_X1   g666(.A1(new_n852), .A2(new_n515), .A3(new_n308), .A4(new_n658), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n853), .A2(new_n305), .A3(new_n655), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n851), .B1(new_n724), .B2(new_n854), .ZN(G75));
  NAND2_X1  g669(.A1(new_n833), .A2(new_n843), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n856), .A2(new_n292), .A3(new_n361), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT56), .ZN(new_n858));
  AOI21_X1  g672(.A(KEYINPUT118), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n857), .A2(KEYINPUT118), .A3(new_n858), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n346), .A2(new_n347), .ZN(new_n861));
  XOR2_X1   g675(.A(new_n861), .B(KEYINPUT117), .Z(new_n862));
  XOR2_X1   g676(.A(new_n315), .B(KEYINPUT55), .Z(new_n863));
  XNOR2_X1  g677(.A(new_n862), .B(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n859), .B1(new_n860), .B2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT118), .ZN(new_n866));
  AOI211_X1 g680(.A(new_n293), .B(new_n360), .C1(new_n833), .C2(new_n843), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n866), .B(new_n864), .C1(new_n867), .C2(KEYINPUT56), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n187), .A2(G952), .ZN(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n865), .A2(new_n871), .ZN(G51));
  INV_X1    g686(.A(new_n844), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n834), .B1(new_n833), .B2(new_n843), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n701), .B(KEYINPUT57), .ZN(new_n876));
  OAI22_X1  g690(.A1(new_n875), .A2(new_n876), .B1(new_n297), .B2(new_n296), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n293), .B1(new_n833), .B2(new_n843), .ZN(new_n878));
  INV_X1    g692(.A(new_n743), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n869), .B1(new_n877), .B2(new_n880), .ZN(G54));
  NAND3_X1  g695(.A1(new_n878), .A2(KEYINPUT58), .A3(G475), .ZN(new_n882));
  INV_X1    g696(.A(new_n465), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n882), .A2(new_n883), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n884), .A2(new_n885), .A3(new_n869), .ZN(G60));
  XNOR2_X1  g700(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n410), .A2(new_n303), .ZN(new_n888));
  XOR2_X1   g702(.A(new_n887), .B(new_n888), .Z(new_n889));
  OAI211_X1 g703(.A(new_n604), .B(new_n889), .C1(new_n873), .C2(new_n874), .ZN(new_n890));
  INV_X1    g704(.A(new_n889), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n891), .B1(new_n849), .B2(new_n844), .ZN(new_n892));
  OAI211_X1 g706(.A(new_n890), .B(new_n870), .C1(new_n892), .C2(new_n604), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(G63));
  NAND2_X1  g708(.A1(G217), .A2(G902), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT120), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT60), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n856), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n505), .B(KEYINPUT121), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n856), .A2(new_n625), .A3(new_n897), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n900), .A2(new_n870), .A3(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT61), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n900), .A2(KEYINPUT61), .A3(new_n870), .A4(new_n901), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(G66));
  OAI21_X1  g720(.A(G953), .B1(new_n373), .B2(new_n313), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n818), .A2(new_n831), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n907), .B1(new_n908), .B2(G953), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n909), .B(KEYINPUT122), .Z(new_n910));
  OAI21_X1  g724(.A(new_n862), .B1(G898), .B2(new_n187), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n910), .B(new_n911), .ZN(G69));
  AOI21_X1  g726(.A(new_n187), .B1(G227), .B2(G900), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n752), .A2(new_n758), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n748), .A2(new_n587), .A3(new_n662), .A4(new_n808), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n647), .A2(new_n803), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n713), .A2(new_n916), .A3(new_n722), .A4(new_n917), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n187), .B1(new_n915), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n636), .A2(G953), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n919), .A2(KEYINPUT124), .A3(new_n920), .ZN(new_n921));
  OR2_X1    g735(.A1(new_n920), .A2(KEYINPUT124), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n921), .A2(KEYINPUT125), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(KEYINPUT125), .B1(new_n921), .B2(new_n922), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n434), .A2(new_n435), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n578), .B(new_n925), .Z(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n923), .A2(new_n924), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n917), .A2(new_n666), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT123), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n930), .A2(KEYINPUT62), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n929), .B(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(new_n915), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n588), .A2(new_n589), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n934), .A2(new_n663), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n815), .A2(new_n750), .ZN(new_n936));
  AOI22_X1  g750(.A1(new_n935), .A2(new_n936), .B1(new_n930), .B2(KEYINPUT62), .ZN(new_n937));
  AND3_X1   g751(.A1(new_n932), .A2(new_n933), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n927), .A2(new_n187), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n914), .B1(new_n928), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n921), .A2(new_n922), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT125), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n921), .A2(KEYINPUT125), .A3(new_n922), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n944), .A2(new_n926), .A3(new_n945), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n946), .B(new_n913), .C1(new_n938), .C2(new_n939), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n941), .A2(new_n947), .ZN(G72));
  NAND2_X1  g762(.A1(new_n938), .A2(new_n908), .ZN(new_n949));
  NAND2_X1  g763(.A1(G472), .A2(G902), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(KEYINPUT63), .Z(new_n951));
  AOI21_X1  g765(.A(new_n552), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n579), .B(KEYINPUT126), .Z(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n869), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n951), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n915), .A2(new_n918), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n956), .B1(new_n957), .B2(new_n908), .ZN(new_n958));
  OR2_X1    g772(.A1(new_n958), .A2(KEYINPUT127), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(KEYINPUT127), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n959), .A2(new_n552), .A3(new_n953), .A4(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n556), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n579), .A2(new_n551), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n848), .B(new_n951), .C1(new_n962), .C2(new_n963), .ZN(new_n964));
  AND3_X1   g778(.A1(new_n955), .A2(new_n961), .A3(new_n964), .ZN(G57));
endmodule


