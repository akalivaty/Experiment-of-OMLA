//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 1 1 0 0 1 1 1 0 1 0 1 1 0 0 1 0 0 0 0 0 0 0 0 0 0 1 1 0 1 0 0 0 1 0 1 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n843, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1011, new_n1012, new_n1013, new_n1015, new_n1016,
    new_n1017, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1064, new_n1065;
  INV_X1    g000(.A(KEYINPUT5), .ZN(new_n202));
  NOR2_X1   g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT72), .ZN(new_n204));
  INV_X1    g003(.A(G141gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G148gat), .ZN(new_n206));
  INV_X1    g005(.A(G148gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G141gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT2), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n204), .A2(new_n212), .A3(new_n210), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT73), .ZN(new_n214));
  XNOR2_X1  g013(.A(G155gat), .B(G162gat), .ZN(new_n215));
  AND4_X1   g014(.A1(new_n214), .A2(new_n209), .A3(new_n215), .A4(new_n211), .ZN(new_n216));
  AOI22_X1  g015(.A1(new_n206), .A2(new_n208), .B1(KEYINPUT2), .B2(new_n210), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n214), .B1(new_n217), .B2(new_n215), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n213), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G134gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G127gat), .ZN(new_n221));
  INV_X1    g020(.A(G127gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G134gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT1), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n221), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G120gat), .ZN(new_n226));
  NOR3_X1   g025(.A1(new_n226), .A2(KEYINPUT67), .A3(G113gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(G113gat), .B(G120gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(KEYINPUT67), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(G113gat), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n232), .A2(G120gat), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n226), .A2(G113gat), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n224), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n221), .A2(new_n223), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n231), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n219), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n209), .A2(new_n215), .A3(new_n211), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(KEYINPUT73), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n217), .A2(new_n214), .A3(new_n215), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  AOI22_X1  g042(.A1(new_n228), .A2(new_n230), .B1(new_n235), .B2(new_n236), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n243), .A2(new_n244), .A3(new_n213), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n239), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(G225gat), .A2(G233gat), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n202), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n219), .A2(KEYINPUT75), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT75), .ZN(new_n251));
  OAI211_X1 g050(.A(new_n251), .B(new_n213), .C1(new_n216), .C2(new_n218), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n250), .A2(new_n244), .A3(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT76), .ZN(new_n254));
  AND3_X1   g053(.A1(new_n253), .A2(new_n254), .A3(KEYINPUT4), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n254), .B1(new_n253), .B2(KEYINPUT4), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n245), .A2(KEYINPUT4), .ZN(new_n257));
  NOR3_X1   g056(.A1(new_n255), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n219), .A2(KEYINPUT3), .ZN(new_n259));
  XOR2_X1   g058(.A(KEYINPUT74), .B(KEYINPUT3), .Z(new_n260));
  OAI211_X1 g059(.A(new_n213), .B(new_n260), .C1(new_n216), .C2(new_n218), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n259), .A2(new_n238), .A3(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n263), .A2(new_n248), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n249), .B1(new_n258), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT6), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT77), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n269));
  AOI22_X1  g068(.A1(new_n209), .A2(new_n211), .B1(G155gat), .B2(G162gat), .ZN(new_n270));
  AOI22_X1  g069(.A1(new_n241), .A2(new_n242), .B1(new_n204), .B2(new_n270), .ZN(new_n271));
  AOI211_X1 g070(.A(new_n268), .B(new_n269), .C1(new_n271), .C2(new_n244), .ZN(new_n272));
  AOI21_X1  g071(.A(KEYINPUT77), .B1(new_n245), .B2(KEYINPUT4), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n250), .A2(new_n269), .A3(new_n244), .A4(new_n252), .ZN(new_n275));
  AOI21_X1  g074(.A(KEYINPUT78), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g075(.A(KEYINPUT4), .B1(new_n219), .B2(new_n238), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(new_n268), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n245), .A2(KEYINPUT77), .A3(KEYINPUT4), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n278), .A2(new_n275), .A3(KEYINPUT78), .A4(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  OAI211_X1 g080(.A(new_n202), .B(new_n264), .C1(new_n276), .C2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G1gat), .B(G29gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n283), .B(KEYINPUT0), .ZN(new_n284));
  XNOR2_X1  g083(.A(G57gat), .B(G85gat), .ZN(new_n285));
  XOR2_X1   g084(.A(new_n284), .B(new_n285), .Z(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n266), .A2(new_n267), .A3(new_n282), .A4(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n286), .A2(KEYINPUT6), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n287), .A2(new_n267), .ZN(new_n290));
  INV_X1    g089(.A(new_n249), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n253), .A2(KEYINPUT4), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT76), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n253), .A2(new_n254), .A3(KEYINPUT4), .ZN(new_n294));
  INV_X1    g093(.A(new_n257), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n293), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n291), .B1(new_n296), .B2(new_n264), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n262), .A2(new_n202), .A3(new_n247), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n278), .A2(new_n275), .A3(new_n279), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT78), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n298), .B1(new_n301), .B2(new_n280), .ZN(new_n302));
  OAI211_X1 g101(.A(new_n289), .B(new_n290), .C1(new_n297), .C2(new_n302), .ZN(new_n303));
  AND2_X1   g102(.A1(new_n288), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT37), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT22), .ZN(new_n306));
  INV_X1    g105(.A(G211gat), .ZN(new_n307));
  INV_X1    g106(.A(G218gat), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n306), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NOR2_X1   g108(.A1(G197gat), .A2(G204gat), .ZN(new_n310));
  AND2_X1   g109(.A1(G197gat), .A2(G204gat), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(G211gat), .B(G218gat), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  OR2_X1    g114(.A1(new_n311), .A2(new_n310), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n316), .A2(new_n313), .A3(new_n309), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT69), .ZN(new_n320));
  INV_X1    g119(.A(G226gat), .ZN(new_n321));
  INV_X1    g120(.A(G233gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  AND2_X1   g123(.A1(G183gat), .A2(G190gat), .ZN(new_n325));
  INV_X1    g124(.A(G183gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(KEYINPUT27), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT27), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(G183gat), .ZN(new_n329));
  INV_X1    g128(.A(G190gat), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n327), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT28), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(KEYINPUT65), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n325), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(KEYINPUT27), .B(G183gat), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n335), .A2(KEYINPUT65), .A3(new_n332), .A4(new_n330), .ZN(new_n336));
  AND2_X1   g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(G169gat), .ZN(new_n338));
  INV_X1    g137(.A(G176gat), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n338), .A2(new_n339), .A3(KEYINPUT66), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(KEYINPUT26), .ZN(new_n341));
  NAND2_X1  g140(.A1(G169gat), .A2(G176gat), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT64), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(KEYINPUT64), .A2(G169gat), .A3(G176gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT26), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n347), .A2(new_n338), .A3(new_n339), .A4(KEYINPUT66), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n341), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT25), .ZN(new_n350));
  XNOR2_X1  g149(.A(G183gat), .B(G190gat), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT24), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n346), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT23), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n354), .A2(new_n338), .A3(new_n339), .ZN(new_n355));
  OAI21_X1  g154(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n325), .A2(new_n352), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n350), .B1(new_n353), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n326), .A2(G190gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n330), .A2(G183gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI22_X1  g162(.A1(new_n363), .A2(KEYINPUT24), .B1(new_n344), .B2(new_n345), .ZN(new_n364));
  AOI22_X1  g163(.A1(new_n355), .A2(new_n356), .B1(new_n352), .B2(new_n325), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n364), .A2(KEYINPUT25), .A3(new_n365), .ZN(new_n366));
  AOI22_X1  g165(.A1(new_n337), .A2(new_n349), .B1(new_n360), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n324), .B1(new_n367), .B2(KEYINPUT29), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n360), .A2(new_n366), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n334), .A2(new_n349), .A3(new_n336), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n324), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n320), .B1(new_n368), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n363), .A2(KEYINPUT24), .ZN(new_n374));
  AND4_X1   g173(.A1(KEYINPUT25), .A2(new_n374), .A3(new_n365), .A4(new_n346), .ZN(new_n375));
  AOI21_X1  g174(.A(KEYINPUT25), .B1(new_n364), .B2(new_n365), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n370), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT29), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n323), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n379), .A2(KEYINPUT69), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n319), .B1(new_n373), .B2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT70), .ZN(new_n382));
  NOR3_X1   g181(.A1(new_n379), .A2(new_n319), .A3(new_n371), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n381), .A2(new_n382), .A3(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(KEYINPUT69), .B1(new_n379), .B2(new_n371), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n368), .A2(new_n320), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n318), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(KEYINPUT70), .B1(new_n388), .B2(new_n383), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n305), .B1(new_n385), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n386), .A2(new_n387), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n383), .B1(new_n391), .B2(new_n319), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(new_n305), .ZN(new_n393));
  XNOR2_X1  g192(.A(G8gat), .B(G36gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n394), .B(KEYINPUT71), .ZN(new_n395));
  XNOR2_X1  g194(.A(G64gat), .B(G92gat), .ZN(new_n396));
  XOR2_X1   g195(.A(new_n395), .B(new_n396), .Z(new_n397));
  NAND2_X1  g196(.A1(new_n393), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(KEYINPUT38), .B1(new_n390), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n397), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n381), .A2(new_n400), .A3(new_n384), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n391), .A2(new_n318), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n379), .A2(new_n371), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n305), .B1(new_n403), .B2(new_n319), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT38), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n393), .A2(new_n405), .A3(new_n397), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n304), .A2(new_n399), .A3(new_n401), .A4(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(G78gat), .B(G106gat), .ZN(new_n408));
  INV_X1    g207(.A(G50gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n408), .B(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT29), .B1(new_n315), .B2(new_n317), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n219), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(G228gat), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n413), .A2(new_n322), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n259), .A2(new_n412), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n318), .B1(new_n261), .B2(new_n378), .ZN(new_n416));
  OAI21_X1  g215(.A(KEYINPUT80), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n261), .A2(new_n378), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(new_n319), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT80), .ZN(new_n420));
  INV_X1    g219(.A(new_n414), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n421), .B1(new_n219), .B2(KEYINPUT3), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n419), .A2(new_n420), .A3(new_n412), .A4(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n417), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(G22gat), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n312), .A2(new_n314), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n313), .B1(new_n316), .B2(new_n309), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n378), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  AOI22_X1  g227(.A1(new_n250), .A2(new_n252), .B1(new_n260), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n421), .B1(new_n429), .B2(new_n416), .ZN(new_n430));
  AND3_X1   g229(.A1(new_n424), .A2(new_n425), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n425), .B1(new_n424), .B2(new_n430), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n410), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT3), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n414), .B1(new_n271), .B2(new_n434), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n271), .A2(new_n428), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n420), .B1(new_n437), .B2(new_n419), .ZN(new_n438));
  NOR3_X1   g237(.A1(new_n415), .A2(KEYINPUT80), .A3(new_n416), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n430), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(G22gat), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n424), .A2(new_n425), .A3(new_n430), .ZN(new_n442));
  INV_X1    g241(.A(new_n410), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  XNOR2_X1  g243(.A(KEYINPUT79), .B(KEYINPUT31), .ZN(new_n445));
  AND3_X1   g244(.A1(new_n433), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n445), .B1(new_n433), .B2(new_n444), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n287), .B1(new_n297), .B2(new_n302), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT40), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n301), .A2(new_n280), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n247), .B1(new_n451), .B2(new_n262), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT39), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n287), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n246), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n453), .B1(new_n455), .B2(new_n247), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n263), .B1(new_n301), .B2(new_n280), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n456), .B1(new_n457), .B2(new_n247), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n450), .B1(new_n454), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n262), .B1(new_n276), .B2(new_n281), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n460), .A2(new_n453), .A3(new_n248), .ZN(new_n461));
  AND4_X1   g260(.A1(new_n450), .A2(new_n461), .A3(new_n458), .A4(new_n286), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n449), .B1(new_n459), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT30), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n464), .B1(new_n392), .B2(new_n400), .ZN(new_n465));
  NOR4_X1   g264(.A1(new_n388), .A2(KEYINPUT30), .A3(new_n397), .A4(new_n383), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n400), .B1(new_n385), .B2(new_n389), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT81), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n401), .A2(KEYINPUT30), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n392), .A2(new_n464), .A3(new_n400), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n382), .B1(new_n381), .B2(new_n384), .ZN(new_n473));
  NOR3_X1   g272(.A1(new_n388), .A2(KEYINPUT70), .A3(new_n383), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n397), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT81), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n472), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n469), .A2(new_n477), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n407), .B(new_n448), .C1(new_n463), .C2(new_n478), .ZN(new_n479));
  XNOR2_X1  g278(.A(new_n377), .B(new_n244), .ZN(new_n480));
  AND2_X1   g279(.A1(G227gat), .A2(G233gat), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT32), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT33), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n484), .B1(new_n480), .B2(new_n482), .ZN(new_n485));
  XOR2_X1   g284(.A(G15gat), .B(G43gat), .Z(new_n486));
  XNOR2_X1  g285(.A(G71gat), .B(G99gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n486), .B(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n483), .A2(new_n485), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n367), .A2(new_n244), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n377), .A2(new_n238), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n490), .A2(new_n482), .A3(new_n491), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n492), .B(KEYINPUT34), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n482), .B1(new_n490), .B2(new_n491), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n488), .B1(new_n494), .B2(KEYINPUT33), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT32), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  AND3_X1   g297(.A1(new_n489), .A2(new_n493), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n493), .B1(new_n489), .B2(new_n498), .ZN(new_n500));
  NOR3_X1   g299(.A1(new_n499), .A2(new_n500), .A3(KEYINPUT36), .ZN(new_n501));
  INV_X1    g300(.A(new_n498), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n495), .A2(new_n497), .ZN(new_n503));
  INV_X1    g302(.A(new_n493), .ZN(new_n504));
  OAI22_X1  g303(.A1(new_n502), .A2(new_n503), .B1(new_n504), .B2(KEYINPUT68), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n489), .A2(new_n493), .A3(new_n498), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n505), .B1(KEYINPUT68), .B2(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n501), .B1(new_n507), .B2(KEYINPUT36), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n433), .A2(new_n444), .ZN(new_n509));
  INV_X1    g308(.A(new_n445), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n433), .A2(new_n444), .A3(new_n445), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n288), .A2(new_n303), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n514), .A2(new_n475), .A3(new_n472), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n508), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n511), .A2(new_n507), .A3(new_n512), .ZN(new_n517));
  OAI21_X1  g316(.A(KEYINPUT35), .B1(new_n517), .B2(new_n515), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n504), .B1(new_n502), .B2(new_n503), .ZN(new_n519));
  AOI21_X1  g318(.A(KEYINPUT35), .B1(new_n519), .B2(new_n506), .ZN(new_n520));
  AND2_X1   g319(.A1(new_n520), .A2(new_n514), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n478), .A2(new_n521), .A3(new_n448), .ZN(new_n522));
  AOI22_X1  g321(.A1(new_n479), .A2(new_n516), .B1(new_n518), .B2(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(G15gat), .B(G22gat), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT16), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n524), .B1(new_n525), .B2(G1gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT86), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT86), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n524), .B(new_n528), .C1(new_n525), .C2(G1gat), .ZN(new_n529));
  XOR2_X1   g328(.A(G15gat), .B(G22gat), .Z(new_n530));
  INV_X1    g329(.A(G1gat), .ZN(new_n531));
  AOI21_X1  g330(.A(G8gat), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n527), .A2(new_n529), .A3(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT87), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n527), .A2(KEYINPUT87), .A3(new_n532), .A4(new_n529), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n526), .B1(G1gat), .B2(new_n524), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(G8gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT88), .ZN(new_n541));
  NOR2_X1   g340(.A1(G29gat), .A2(G36gat), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT14), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n542), .B1(KEYINPUT82), .B2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(KEYINPUT82), .B(KEYINPUT14), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n544), .B1(new_n545), .B2(new_n542), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT15), .ZN(new_n547));
  OR2_X1    g346(.A1(G43gat), .A2(G50gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(G43gat), .A2(G50gat), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(G29gat), .A2(G36gat), .ZN(new_n552));
  AND3_X1   g351(.A1(new_n546), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(KEYINPUT84), .B(G43gat), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n554), .A2(G50gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(KEYINPUT85), .B(G50gat), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n556), .A2(G43gat), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n547), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  AND2_X1   g357(.A1(new_n553), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT83), .ZN(new_n560));
  AOI22_X1  g359(.A1(new_n546), .A2(new_n560), .B1(G29gat), .B2(G36gat), .ZN(new_n561));
  OAI211_X1 g360(.A(KEYINPUT83), .B(new_n544), .C1(new_n545), .C2(new_n542), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n551), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  OAI211_X1 g362(.A(new_n541), .B(KEYINPUT17), .C1(new_n559), .C2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n546), .A2(new_n560), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n565), .A2(new_n562), .A3(new_n552), .ZN(new_n566));
  AOI22_X1  g365(.A1(new_n566), .A2(new_n550), .B1(new_n553), .B2(new_n558), .ZN(new_n567));
  OR2_X1    g366(.A1(new_n541), .A2(KEYINPUT17), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n541), .A2(KEYINPUT17), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n540), .B1(new_n564), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(G229gat), .A2(G233gat), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  AOI22_X1  g372(.A1(new_n535), .A2(new_n536), .B1(G8gat), .B2(new_n538), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n574), .A2(new_n567), .ZN(new_n575));
  NOR3_X1   g374(.A1(new_n571), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  OAI21_X1  g375(.A(KEYINPUT89), .B1(new_n576), .B2(KEYINPUT18), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n570), .A2(new_n564), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(new_n574), .ZN(new_n579));
  INV_X1    g378(.A(new_n575), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n579), .A2(new_n572), .A3(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT89), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT18), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  AND2_X1   g383(.A1(new_n577), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n579), .A2(KEYINPUT18), .A3(new_n572), .A4(new_n580), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n574), .B(new_n567), .ZN(new_n587));
  XOR2_X1   g386(.A(new_n572), .B(KEYINPUT13), .Z(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(G113gat), .B(G141gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(G197gat), .ZN(new_n591));
  XOR2_X1   g390(.A(KEYINPUT11), .B(G169gat), .Z(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT12), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n586), .A2(new_n589), .A3(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  AOI22_X1  g395(.A1(new_n576), .A2(KEYINPUT18), .B1(new_n587), .B2(new_n588), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n575), .B1(new_n578), .B2(new_n574), .ZN(new_n598));
  AOI21_X1  g397(.A(KEYINPUT18), .B1(new_n598), .B2(new_n572), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n594), .ZN(new_n602));
  AOI22_X1  g401(.A1(new_n585), .A2(new_n596), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n523), .A2(new_n603), .ZN(new_n604));
  AND2_X1   g403(.A1(G232gat), .A2(G233gat), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n605), .A2(KEYINPUT41), .ZN(new_n606));
  XNOR2_X1  g405(.A(G134gat), .B(G162gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  XOR2_X1   g408(.A(G190gat), .B(G218gat), .Z(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  OR2_X1    g410(.A1(G99gat), .A2(G106gat), .ZN(new_n612));
  NAND2_X1  g411(.A1(G99gat), .A2(G106gat), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(G85gat), .A2(G92gat), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT7), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n613), .A2(KEYINPUT8), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n618), .B1(G85gat), .B2(G92gat), .ZN(new_n619));
  OAI211_X1 g418(.A(KEYINPUT94), .B(new_n614), .C1(new_n617), .C2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n614), .A2(KEYINPUT94), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n615), .B(KEYINPUT7), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT94), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n612), .A2(new_n623), .A3(new_n613), .ZN(new_n624));
  INV_X1    g423(.A(G85gat), .ZN(new_n625));
  INV_X1    g424(.A(G92gat), .ZN(new_n626));
  AOI22_X1  g425(.A1(KEYINPUT8), .A2(new_n613), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n621), .A2(new_n622), .A3(new_n624), .A4(new_n627), .ZN(new_n628));
  AND3_X1   g427(.A1(new_n620), .A2(new_n628), .A3(KEYINPUT95), .ZN(new_n629));
  AOI21_X1  g428(.A(KEYINPUT95), .B1(new_n620), .B2(new_n628), .ZN(new_n630));
  OR2_X1    g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n578), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n605), .A2(KEYINPUT41), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n633), .B1(new_n631), .B2(new_n567), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n611), .B1(new_n632), .B2(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n629), .A2(new_n630), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n637), .B1(new_n570), .B2(new_n564), .ZN(new_n638));
  NOR3_X1   g437(.A1(new_n638), .A2(new_n610), .A3(new_n634), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n609), .B1(new_n636), .B2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n632), .A2(new_n635), .A3(new_n611), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n610), .B1(new_n638), .B2(new_n634), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n641), .A2(new_n608), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(G57gat), .ZN(new_n645));
  OAI21_X1  g444(.A(G64gat), .B1(new_n645), .B2(KEYINPUT91), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT91), .ZN(new_n647));
  INV_X1    g446(.A(G64gat), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n647), .A2(new_n648), .A3(G57gat), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(G71gat), .ZN(new_n651));
  INV_X1    g450(.A(G78gat), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n651), .A2(new_n652), .A3(KEYINPUT9), .ZN(new_n653));
  NAND2_X1  g452(.A1(G71gat), .A2(G78gat), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n650), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT90), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n658), .A2(new_n651), .A3(new_n652), .ZN(new_n659));
  OAI21_X1  g458(.A(KEYINPUT90), .B1(G71gat), .B2(G78gat), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n659), .A2(new_n654), .A3(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT9), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n648), .A2(G57gat), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n645), .A2(G64gat), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n662), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n657), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n667), .A2(KEYINPUT21), .ZN(new_n668));
  XNOR2_X1  g467(.A(G127gat), .B(G155gat), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n668), .B(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n656), .B1(new_n665), .B2(new_n661), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT93), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  OAI211_X1 g473(.A(new_n656), .B(KEYINPUT93), .C1(new_n665), .C2(new_n661), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n674), .A2(KEYINPUT21), .A3(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n671), .A2(new_n676), .A3(new_n574), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n668), .B(new_n669), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n574), .A2(new_n676), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(G231gat), .A2(G233gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT92), .ZN(new_n683));
  XOR2_X1   g482(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(G183gat), .B(G211gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n681), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n677), .A2(new_n680), .A3(new_n687), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n667), .A2(new_n620), .A3(new_n628), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n620), .A2(new_n628), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(new_n672), .ZN(new_n695));
  INV_X1    g494(.A(G230gat), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n696), .A2(new_n322), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n693), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT97), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g499(.A1(new_n693), .A2(new_n695), .A3(KEYINPUT97), .A4(new_n697), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g501(.A(G120gat), .B(G148gat), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT98), .ZN(new_n704));
  XNOR2_X1  g503(.A(G176gat), .B(G204gat), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n704), .B(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n702), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT10), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n695), .ZN(new_n710));
  AND3_X1   g509(.A1(new_n674), .A2(KEYINPUT10), .A3(new_n675), .ZN(new_n711));
  AOI22_X1  g510(.A1(new_n709), .A2(new_n710), .B1(new_n637), .B2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(KEYINPUT96), .B1(new_n712), .B2(new_n697), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT96), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n674), .A2(KEYINPUT10), .A3(new_n675), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n715), .A2(new_n629), .A3(new_n630), .ZN(new_n716));
  AOI21_X1  g515(.A(KEYINPUT10), .B1(new_n693), .B2(new_n695), .ZN(new_n717));
  OAI221_X1 g516(.A(new_n714), .B1(new_n696), .B2(new_n322), .C1(new_n716), .C2(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n708), .A2(new_n713), .A3(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n712), .A2(new_n697), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n707), .B1(new_n720), .B2(new_n702), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  AND3_X1   g522(.A1(new_n644), .A2(new_n692), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n604), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n725), .A2(new_n514), .ZN(new_n726));
  XNOR2_X1  g525(.A(KEYINPUT99), .B(G1gat), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(G1324gat));
  INV_X1    g527(.A(G8gat), .ZN(new_n729));
  INV_X1    g528(.A(new_n725), .ZN(new_n730));
  INV_X1    g529(.A(new_n478), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  XNOR2_X1  g531(.A(KEYINPUT16), .B(G8gat), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n725), .A2(new_n478), .A3(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(KEYINPUT42), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n735), .B1(KEYINPUT42), .B2(new_n734), .ZN(G1325gat));
  NOR2_X1   g535(.A1(new_n499), .A2(new_n500), .ZN(new_n737));
  OR3_X1    g536(.A1(new_n725), .A2(G15gat), .A3(new_n737), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n506), .A2(KEYINPUT68), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT68), .ZN(new_n740));
  AOI22_X1  g539(.A1(new_n489), .A2(new_n498), .B1(new_n493), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(KEYINPUT36), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n737), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n742), .B1(new_n743), .B2(KEYINPUT36), .ZN(new_n744));
  OAI21_X1  g543(.A(G15gat), .B1(new_n725), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n738), .A2(new_n745), .ZN(G1326gat));
  INV_X1    g545(.A(KEYINPUT100), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n730), .A2(new_n747), .A3(new_n513), .ZN(new_n748));
  OAI21_X1  g547(.A(KEYINPUT100), .B1(new_n725), .B2(new_n448), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g549(.A(KEYINPUT43), .B(G22gat), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n748), .A2(new_n749), .A3(new_n751), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(G1327gat));
  INV_X1    g554(.A(KEYINPUT44), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n756), .B1(new_n523), .B2(new_n644), .ZN(new_n757));
  INV_X1    g556(.A(new_n644), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n472), .A2(new_n475), .ZN(new_n759));
  OAI22_X1  g558(.A1(new_n304), .A2(new_n759), .B1(new_n446), .B2(new_n447), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(new_n744), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n461), .A2(new_n458), .A3(new_n286), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(KEYINPUT40), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n454), .A2(new_n450), .A3(new_n458), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n765), .A2(new_n469), .A3(new_n477), .A4(new_n449), .ZN(new_n766));
  AND4_X1   g565(.A1(new_n288), .A2(new_n406), .A3(new_n303), .A4(new_n401), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n513), .B1(new_n767), .B2(new_n399), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n761), .B1(new_n766), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n304), .A2(new_n759), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n770), .A2(new_n448), .A3(new_n507), .ZN(new_n771));
  AND4_X1   g570(.A1(new_n514), .A2(new_n511), .A3(new_n520), .A4(new_n512), .ZN(new_n772));
  AOI22_X1  g571(.A1(new_n771), .A2(KEYINPUT35), .B1(new_n772), .B2(new_n478), .ZN(new_n773));
  OAI211_X1 g572(.A(KEYINPUT44), .B(new_n758), .C1(new_n769), .C2(new_n773), .ZN(new_n774));
  XOR2_X1   g573(.A(new_n722), .B(KEYINPUT101), .Z(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n776), .A2(new_n603), .A3(new_n692), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n757), .A2(new_n774), .A3(new_n777), .ZN(new_n778));
  OAI21_X1  g577(.A(G29gat), .B1(new_n778), .B2(new_n514), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT45), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n644), .A2(new_n692), .A3(new_n722), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n604), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n514), .A2(G29gat), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n780), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n604), .A2(KEYINPUT45), .A3(new_n781), .A4(new_n783), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n779), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT102), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n779), .A2(new_n785), .A3(KEYINPUT102), .A4(new_n786), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(G1328gat));
  NOR3_X1   g590(.A1(new_n782), .A2(G36gat), .A3(new_n478), .ZN(new_n792));
  NAND2_X1  g591(.A1(KEYINPUT103), .A2(KEYINPUT46), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(G36gat), .B1(new_n778), .B2(new_n478), .ZN(new_n795));
  XOR2_X1   g594(.A(KEYINPUT103), .B(KEYINPUT46), .Z(new_n796));
  OAI211_X1 g595(.A(new_n794), .B(new_n795), .C1(new_n792), .C2(new_n796), .ZN(G1329gat));
  OAI21_X1  g596(.A(new_n554), .B1(new_n782), .B2(new_n737), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n744), .A2(new_n554), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n757), .A2(new_n774), .A3(new_n777), .A4(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT104), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(KEYINPUT47), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n798), .A2(new_n800), .A3(new_n802), .ZN(new_n803));
  OR2_X1    g602(.A1(new_n801), .A2(KEYINPUT47), .ZN(new_n804));
  XNOR2_X1  g603(.A(new_n803), .B(new_n804), .ZN(G1330gat));
  NAND4_X1  g604(.A1(new_n757), .A2(new_n513), .A3(new_n774), .A4(new_n777), .ZN(new_n806));
  INV_X1    g605(.A(new_n556), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n448), .A2(new_n807), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(KEYINPUT106), .ZN(new_n810));
  INV_X1    g609(.A(new_n781), .ZN(new_n811));
  NOR4_X1   g610(.A1(new_n523), .A2(new_n810), .A3(new_n603), .A4(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n808), .A2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT105), .ZN(new_n815));
  AOI21_X1  g614(.A(KEYINPUT48), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n812), .B1(new_n806), .B2(new_n807), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT48), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n817), .A2(KEYINPUT105), .A3(new_n818), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n816), .A2(new_n819), .ZN(G1331gat));
  AOI21_X1  g619(.A(new_n691), .B1(new_n640), .B2(new_n643), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n776), .A2(new_n603), .A3(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n523), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(new_n304), .ZN(new_n824));
  XNOR2_X1  g623(.A(new_n824), .B(G57gat), .ZN(G1332gat));
  NOR3_X1   g624(.A1(new_n523), .A2(new_n478), .A3(new_n822), .ZN(new_n826));
  NOR2_X1   g625(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n827));
  AND2_X1   g626(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n826), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n829), .B1(new_n826), .B2(new_n827), .ZN(G1333gat));
  NAND2_X1  g629(.A1(new_n823), .A2(new_n743), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(KEYINPUT107), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT107), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n823), .A2(new_n833), .A3(new_n743), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n832), .A2(new_n651), .A3(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n823), .A2(G71gat), .A3(new_n508), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g636(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n835), .A2(new_n836), .A3(new_n838), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(G1334gat));
  NAND2_X1  g641(.A1(new_n823), .A2(new_n513), .ZN(new_n843));
  XNOR2_X1  g642(.A(new_n843), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g643(.A1(new_n586), .A2(new_n589), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n602), .B1(new_n845), .B2(new_n599), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n577), .A2(new_n584), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n846), .B1(new_n847), .B2(new_n595), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n848), .A2(new_n692), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n850), .A2(new_n723), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n757), .A2(new_n774), .A3(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(G85gat), .B1(new_n852), .B2(new_n514), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n523), .A2(new_n644), .A3(new_n850), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n854), .A2(KEYINPUT51), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n758), .B(new_n849), .C1(new_n769), .C2(new_n773), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT51), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n304), .A2(new_n625), .A3(new_n722), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n853), .B1(new_n859), .B2(new_n860), .ZN(G1336gat));
  NOR3_X1   g660(.A1(new_n854), .A2(KEYINPUT110), .A3(new_n857), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT110), .ZN(new_n863));
  AOI21_X1  g662(.A(KEYINPUT51), .B1(new_n856), .B2(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n731), .A2(new_n626), .A3(new_n776), .ZN(new_n865));
  XNOR2_X1  g664(.A(new_n865), .B(KEYINPUT109), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n862), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n757), .A2(new_n731), .A3(new_n774), .A4(new_n851), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(G92gat), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(KEYINPUT52), .B1(new_n867), .B2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT52), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n872), .B(new_n869), .C1(new_n859), .C2(new_n865), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n871), .A2(new_n873), .ZN(G1337gat));
  NOR2_X1   g673(.A1(new_n723), .A2(G99gat), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n743), .B(new_n875), .C1(new_n855), .C2(new_n858), .ZN(new_n876));
  OAI21_X1  g675(.A(G99gat), .B1(new_n852), .B2(new_n744), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(KEYINPUT111), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT111), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n876), .A2(new_n880), .A3(new_n877), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n879), .A2(new_n881), .ZN(G1338gat));
  NOR3_X1   g681(.A1(new_n448), .A2(new_n775), .A3(G106gat), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n862), .A2(new_n864), .A3(new_n884), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n757), .A2(new_n513), .A3(new_n774), .A4(new_n851), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(G106gat), .ZN(new_n887));
  INV_X1    g686(.A(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(KEYINPUT53), .B1(new_n885), .B2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT53), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n890), .B(new_n887), .C1(new_n859), .C2(new_n884), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n889), .A2(new_n891), .ZN(G1339gat));
  INV_X1    g691(.A(KEYINPUT54), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n893), .B1(new_n712), .B2(new_n697), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n713), .A2(new_n894), .A3(new_n718), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n706), .B1(new_n720), .B2(new_n893), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(KEYINPUT55), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT55), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n895), .A2(new_n896), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n848), .A2(new_n644), .A3(new_n901), .A4(new_n719), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n644), .B1(new_n901), .B2(new_n719), .ZN(new_n903));
  AND3_X1   g702(.A1(new_n641), .A2(new_n608), .A3(new_n642), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n608), .B1(new_n641), .B2(new_n642), .ZN(new_n905));
  OAI211_X1 g704(.A(new_n721), .B(new_n719), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(KEYINPUT112), .B1(new_n598), .B2(new_n572), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT112), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n908), .B(new_n573), .C1(new_n571), .C2(new_n575), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n907), .B(new_n909), .C1(new_n587), .C2(new_n588), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(new_n593), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n597), .A2(new_n577), .A3(new_n594), .A4(new_n584), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n906), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n902), .B1(new_n903), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(new_n691), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n821), .A2(new_n912), .A3(new_n846), .A4(new_n723), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(new_n448), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n478), .A2(new_n304), .A3(new_n743), .ZN(new_n919));
  OR2_X1    g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n920), .A2(new_n232), .A3(new_n603), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n917), .A2(new_n304), .A3(new_n478), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n922), .A2(new_n517), .ZN(new_n923));
  AOI21_X1  g722(.A(G113gat), .B1(new_n923), .B2(new_n848), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n921), .A2(new_n924), .ZN(G1340gat));
  NOR3_X1   g724(.A1(new_n920), .A2(new_n226), .A3(new_n775), .ZN(new_n926));
  AOI21_X1  g725(.A(G120gat), .B1(new_n923), .B2(new_n722), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n926), .A2(new_n927), .ZN(G1341gat));
  OAI21_X1  g727(.A(G127gat), .B1(new_n920), .B2(new_n691), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n923), .A2(new_n222), .A3(new_n692), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(G1342gat));
  OAI21_X1  g730(.A(G134gat), .B1(new_n920), .B2(new_n644), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT56), .ZN(new_n933));
  NOR4_X1   g732(.A1(new_n922), .A2(G134gat), .A3(new_n517), .A4(new_n644), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n934), .A2(KEYINPUT113), .A3(new_n933), .ZN(new_n935));
  AOI21_X1  g734(.A(KEYINPUT113), .B1(new_n934), .B2(new_n933), .ZN(new_n936));
  OAI221_X1 g735(.A(new_n932), .B1(new_n933), .B2(new_n934), .C1(new_n935), .C2(new_n936), .ZN(G1343gat));
  XOR2_X1   g736(.A(KEYINPUT115), .B(KEYINPUT57), .Z(new_n938));
  AND3_X1   g737(.A1(new_n906), .A2(new_n911), .A3(new_n912), .ZN(new_n939));
  INV_X1    g738(.A(new_n900), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n899), .B1(new_n895), .B2(new_n896), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n719), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(new_n758), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n939), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n692), .B1(new_n944), .B2(new_n902), .ZN(new_n945));
  INV_X1    g744(.A(new_n916), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n938), .B1(new_n947), .B2(new_n448), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT57), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n917), .A2(new_n949), .A3(new_n513), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n744), .A2(new_n478), .A3(new_n304), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT114), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n951), .A2(new_n952), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n948), .A2(new_n950), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g755(.A(G141gat), .B1(new_n956), .B2(new_n603), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT58), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n508), .A2(new_n448), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n917), .A2(new_n304), .A3(new_n959), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT117), .ZN(new_n961));
  OR2_X1    g760(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n960), .A2(new_n961), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n962), .A2(new_n478), .A3(new_n963), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n603), .A2(G141gat), .ZN(new_n965));
  INV_X1    g764(.A(new_n965), .ZN(new_n966));
  OAI211_X1 g765(.A(new_n957), .B(new_n958), .C1(new_n964), .C2(new_n966), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT116), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n959), .A2(new_n965), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n968), .B1(new_n922), .B2(new_n969), .ZN(new_n970));
  OR3_X1    g769(.A1(new_n922), .A2(new_n968), .A3(new_n969), .ZN(new_n971));
  AND3_X1   g770(.A1(new_n957), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n967), .B1(new_n972), .B2(new_n958), .ZN(G1344gat));
  INV_X1    g772(.A(KEYINPUT59), .ZN(new_n974));
  OAI211_X1 g773(.A(new_n974), .B(G148gat), .C1(new_n956), .C2(new_n723), .ZN(new_n975));
  OAI211_X1 g774(.A(new_n513), .B(new_n938), .C1(new_n945), .C2(new_n946), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT118), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n603), .A2(new_n724), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n916), .A2(KEYINPUT118), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g779(.A(new_n980), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n448), .B1(new_n915), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n976), .B1(new_n982), .B2(KEYINPUT57), .ZN(new_n983));
  NOR3_X1   g782(.A1(new_n953), .A2(new_n954), .A3(new_n723), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n985), .A2(G148gat), .ZN(new_n986));
  AOI21_X1  g785(.A(KEYINPUT119), .B1(new_n986), .B2(KEYINPUT59), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n207), .B1(new_n983), .B2(new_n984), .ZN(new_n988));
  INV_X1    g787(.A(KEYINPUT119), .ZN(new_n989));
  NOR3_X1   g788(.A1(new_n988), .A2(new_n989), .A3(new_n974), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n975), .B1(new_n987), .B2(new_n990), .ZN(new_n991));
  INV_X1    g790(.A(new_n964), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n992), .A2(new_n207), .A3(new_n722), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n991), .A2(new_n993), .ZN(G1345gat));
  OAI21_X1  g793(.A(G155gat), .B1(new_n956), .B2(new_n691), .ZN(new_n995));
  OR2_X1    g794(.A1(new_n691), .A2(G155gat), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n995), .B1(new_n964), .B2(new_n996), .ZN(G1346gat));
  INV_X1    g796(.A(G162gat), .ZN(new_n998));
  NOR3_X1   g797(.A1(new_n956), .A2(new_n998), .A3(new_n644), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n992), .A2(new_n758), .ZN(new_n1000));
  AOI21_X1  g799(.A(new_n999), .B1(new_n1000), .B2(new_n998), .ZN(G1347gat));
  NOR2_X1   g800(.A1(new_n478), .A2(new_n517), .ZN(new_n1002));
  XNOR2_X1  g801(.A(new_n1002), .B(KEYINPUT120), .ZN(new_n1003));
  NOR3_X1   g802(.A1(new_n1003), .A2(new_n947), .A3(new_n304), .ZN(new_n1004));
  AOI21_X1  g803(.A(G169gat), .B1(new_n1004), .B2(new_n848), .ZN(new_n1005));
  NOR3_X1   g804(.A1(new_n478), .A2(new_n304), .A3(new_n737), .ZN(new_n1006));
  XNOR2_X1  g805(.A(new_n1006), .B(KEYINPUT121), .ZN(new_n1007));
  NOR2_X1   g806(.A1(new_n918), .A2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g807(.A1(new_n603), .A2(new_n338), .ZN(new_n1009));
  AOI21_X1  g808(.A(new_n1005), .B1(new_n1008), .B2(new_n1009), .ZN(G1348gat));
  NAND3_X1  g809(.A1(new_n1004), .A2(new_n339), .A3(new_n722), .ZN(new_n1011));
  NOR3_X1   g810(.A1(new_n918), .A2(new_n1007), .A3(new_n775), .ZN(new_n1012));
  OAI21_X1  g811(.A(new_n1011), .B1(new_n339), .B2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g812(.A(new_n1013), .B(KEYINPUT122), .ZN(G1349gat));
  NAND3_X1  g813(.A1(new_n1004), .A2(new_n335), .A3(new_n692), .ZN(new_n1015));
  NOR3_X1   g814(.A1(new_n918), .A2(new_n1007), .A3(new_n691), .ZN(new_n1016));
  OAI21_X1  g815(.A(new_n1015), .B1(new_n326), .B2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g816(.A(new_n1017), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g817(.A1(new_n1004), .A2(new_n330), .A3(new_n758), .ZN(new_n1019));
  INV_X1    g818(.A(KEYINPUT61), .ZN(new_n1020));
  NAND2_X1  g819(.A1(new_n1008), .A2(new_n758), .ZN(new_n1021));
  AOI21_X1  g820(.A(new_n1020), .B1(new_n1021), .B2(G190gat), .ZN(new_n1022));
  AOI211_X1 g821(.A(KEYINPUT61), .B(new_n330), .C1(new_n1008), .C2(new_n758), .ZN(new_n1023));
  OAI21_X1  g822(.A(new_n1019), .B1(new_n1022), .B2(new_n1023), .ZN(G1351gat));
  NOR3_X1   g823(.A1(new_n508), .A2(new_n478), .A3(new_n448), .ZN(new_n1025));
  AND3_X1   g824(.A1(new_n917), .A2(new_n514), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g825(.A(G197gat), .ZN(new_n1027));
  NAND3_X1  g826(.A1(new_n1026), .A2(new_n1027), .A3(new_n848), .ZN(new_n1028));
  XNOR2_X1  g827(.A(new_n1028), .B(KEYINPUT123), .ZN(new_n1029));
  NAND3_X1  g828(.A1(new_n731), .A2(new_n514), .A3(new_n744), .ZN(new_n1030));
  INV_X1    g829(.A(new_n1030), .ZN(new_n1031));
  NAND2_X1  g830(.A1(new_n983), .A2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g831(.A(G197gat), .B1(new_n1032), .B2(new_n603), .ZN(new_n1033));
  NAND2_X1  g832(.A1(new_n1029), .A2(new_n1033), .ZN(G1352gat));
  OAI21_X1  g833(.A(G204gat), .B1(new_n1032), .B2(new_n775), .ZN(new_n1035));
  INV_X1    g834(.A(KEYINPUT62), .ZN(new_n1036));
  NOR2_X1   g835(.A1(new_n723), .A2(G204gat), .ZN(new_n1037));
  NAND4_X1  g836(.A1(new_n1026), .A2(KEYINPUT124), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  INV_X1    g837(.A(KEYINPUT124), .ZN(new_n1039));
  NAND4_X1  g838(.A1(new_n917), .A2(new_n514), .A3(new_n1025), .A4(new_n1037), .ZN(new_n1040));
  OAI21_X1  g839(.A(new_n1039), .B1(new_n1040), .B2(KEYINPUT62), .ZN(new_n1041));
  NAND2_X1  g840(.A1(new_n1038), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g841(.A1(new_n1040), .A2(KEYINPUT62), .ZN(new_n1043));
  NAND3_X1  g842(.A1(new_n1035), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g843(.A(KEYINPUT125), .ZN(new_n1045));
  NAND2_X1  g844(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND4_X1  g845(.A1(new_n1035), .A2(new_n1042), .A3(KEYINPUT125), .A4(new_n1043), .ZN(new_n1047));
  NAND2_X1  g846(.A1(new_n1046), .A2(new_n1047), .ZN(G1353gat));
  INV_X1    g847(.A(KEYINPUT63), .ZN(new_n1049));
  NAND4_X1  g848(.A1(new_n983), .A2(KEYINPUT126), .A3(new_n692), .A4(new_n1031), .ZN(new_n1050));
  NAND2_X1  g849(.A1(new_n1050), .A2(G211gat), .ZN(new_n1051));
  AOI21_X1  g850(.A(new_n980), .B1(new_n691), .B2(new_n914), .ZN(new_n1052));
  OAI21_X1  g851(.A(new_n949), .B1(new_n1052), .B2(new_n448), .ZN(new_n1053));
  AOI21_X1  g852(.A(new_n1030), .B1(new_n1053), .B2(new_n976), .ZN(new_n1054));
  AOI21_X1  g853(.A(KEYINPUT126), .B1(new_n1054), .B2(new_n692), .ZN(new_n1055));
  OAI21_X1  g854(.A(new_n1049), .B1(new_n1051), .B2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g855(.A1(new_n983), .A2(new_n692), .A3(new_n1031), .ZN(new_n1057));
  INV_X1    g856(.A(KEYINPUT126), .ZN(new_n1058));
  NAND2_X1  g857(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND4_X1  g858(.A1(new_n1059), .A2(KEYINPUT63), .A3(G211gat), .A4(new_n1050), .ZN(new_n1060));
  NAND2_X1  g859(.A1(new_n1056), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g860(.A1(new_n1026), .A2(new_n307), .A3(new_n692), .ZN(new_n1062));
  NAND2_X1  g861(.A1(new_n1061), .A2(new_n1062), .ZN(G1354gat));
  OAI21_X1  g862(.A(G218gat), .B1(new_n1032), .B2(new_n644), .ZN(new_n1064));
  NAND3_X1  g863(.A1(new_n1026), .A2(new_n308), .A3(new_n758), .ZN(new_n1065));
  NAND2_X1  g864(.A1(new_n1064), .A2(new_n1065), .ZN(G1355gat));
endmodule


