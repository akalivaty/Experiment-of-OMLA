

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786;

  INV_X2 U377 ( .A(G953), .ZN(n773) );
  XNOR2_X1 U378 ( .A(n489), .B(n488), .ZN(n566) );
  AND2_X2 U379 ( .A1(n716), .A2(n405), .ZN(n401) );
  XNOR2_X1 U380 ( .A(n673), .B(KEYINPUT66), .ZN(n678) );
  XNOR2_X2 U381 ( .A(G119), .B(KEYINPUT71), .ZN(n469) );
  XNOR2_X2 U382 ( .A(n438), .B(G146), .ZN(n412) );
  XNOR2_X2 U383 ( .A(G116), .B(G113), .ZN(n470) );
  XNOR2_X2 U384 ( .A(n480), .B(n358), .ZN(n438) );
  XNOR2_X2 U385 ( .A(n585), .B(n584), .ZN(n621) );
  NOR2_X2 U386 ( .A1(n621), .A2(n781), .ZN(n623) );
  INV_X2 U387 ( .A(G125), .ZN(n403) );
  AND2_X1 U388 ( .A1(n375), .A2(n380), .ZN(n379) );
  NAND2_X1 U389 ( .A1(n712), .A2(n698), .ZN(n659) );
  NOR2_X1 U390 ( .A1(n727), .A2(n637), .ZN(n653) );
  NOR2_X1 U391 ( .A1(n722), .A2(n592), .ZN(n593) );
  XNOR2_X1 U392 ( .A(n432), .B(n431), .ZN(n640) );
  NAND2_X1 U393 ( .A1(n379), .A2(n376), .ZN(n662) );
  XNOR2_X1 U394 ( .A(n668), .B(KEYINPUT84), .ZN(n772) );
  AND2_X1 U395 ( .A1(n646), .A2(n649), .ZN(n644) );
  AND2_X1 U396 ( .A1(n391), .A2(n361), .ZN(n388) );
  OR2_X1 U397 ( .A1(n439), .A2(KEYINPUT35), .ZN(n361) );
  NOR2_X1 U398 ( .A1(n568), .A2(n564), .ZN(n587) );
  NAND2_X1 U399 ( .A1(n464), .A2(n461), .ZN(n596) );
  AND2_X1 U400 ( .A1(n467), .A2(n465), .ZN(n464) );
  BUF_X1 U401 ( .A(n572), .Z(n719) );
  XNOR2_X1 U402 ( .A(n434), .B(n433), .ZN(n602) );
  XNOR2_X1 U403 ( .A(n545), .B(n544), .ZN(n572) );
  XNOR2_X1 U404 ( .A(n396), .B(n395), .ZN(n546) );
  XNOR2_X1 U405 ( .A(n470), .B(n468), .ZN(n396) );
  XNOR2_X1 U406 ( .A(n469), .B(n482), .ZN(n395) );
  INV_X1 U407 ( .A(n453), .ZN(n355) );
  XNOR2_X1 U408 ( .A(n573), .B(n529), .ZN(n716) );
  NAND2_X1 U409 ( .A1(n678), .A2(n750), .ZN(n409) );
  INV_X1 U410 ( .A(n566), .ZN(n586) );
  XNOR2_X1 U411 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U412 ( .A(n650), .B(n558), .ZN(n635) );
  NAND2_X1 U413 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U414 ( .A1(n457), .A2(n362), .ZN(n592) );
  INV_X1 U415 ( .A(n572), .ZN(n457) );
  INV_X1 U416 ( .A(n574), .ZN(n456) );
  XNOR2_X1 U417 ( .A(n502), .B(n532), .ZN(n508) );
  XNOR2_X1 U418 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U419 ( .A(n374), .B(KEYINPUT0), .ZN(n636) );
  NAND2_X1 U420 ( .A1(n596), .A2(n497), .ZN(n374) );
  XNOR2_X1 U421 ( .A(n496), .B(KEYINPUT94), .ZN(n497) );
  AND2_X1 U422 ( .A1(n572), .A2(n720), .ZN(n717) );
  AND2_X1 U423 ( .A1(n586), .A2(n367), .ZN(n451) );
  NOR2_X1 U424 ( .A1(G953), .A2(G237), .ZN(n547) );
  NAND2_X1 U425 ( .A1(n381), .A2(KEYINPUT44), .ZN(n380) );
  XNOR2_X1 U426 ( .A(n377), .B(KEYINPUT107), .ZN(n376) );
  NAND2_X1 U427 ( .A1(n660), .A2(n378), .ZN(n377) );
  NAND2_X1 U428 ( .A1(n659), .A2(n658), .ZN(n378) );
  NOR2_X1 U429 ( .A1(n615), .A2(n614), .ZN(n625) );
  INV_X1 U430 ( .A(G237), .ZN(n484) );
  NOR2_X1 U431 ( .A1(n734), .A2(n563), .ZN(n521) );
  INV_X1 U432 ( .A(KEYINPUT4), .ZN(n404) );
  NAND2_X1 U433 ( .A1(n602), .A2(n430), .ZN(n734) );
  INV_X1 U434 ( .A(n640), .ZN(n430) );
  NAND2_X1 U435 ( .A1(n714), .A2(KEYINPUT34), .ZN(n439) );
  INV_X1 U436 ( .A(KEYINPUT19), .ZN(n463) );
  NAND2_X1 U437 ( .A1(n466), .A2(KEYINPUT19), .ZN(n465) );
  NOR2_X1 U438 ( .A1(n768), .A2(G902), .ZN(n545) );
  INV_X1 U439 ( .A(KEYINPUT70), .ZN(n482) );
  XNOR2_X1 U440 ( .A(n429), .B(n428), .ZN(n539) );
  INV_X1 U441 ( .A(KEYINPUT8), .ZN(n428) );
  NAND2_X1 U442 ( .A1(n773), .A2(G234), .ZN(n429) );
  XNOR2_X1 U443 ( .A(n532), .B(n460), .ZN(n771) );
  INV_X1 U444 ( .A(n531), .ZN(n460) );
  XNOR2_X1 U445 ( .A(n579), .B(KEYINPUT39), .ZN(n581) );
  NAND2_X1 U446 ( .A1(n578), .A2(n732), .ZN(n579) );
  NOR2_X1 U447 ( .A1(n453), .A2(n450), .ZN(n449) );
  NOR2_X1 U448 ( .A1(n586), .A2(n367), .ZN(n450) );
  NOR2_X1 U449 ( .A1(n708), .A2(n466), .ZN(n454) );
  INV_X1 U450 ( .A(n592), .ZN(n455) );
  NAND2_X1 U451 ( .A1(n439), .A2(KEYINPUT35), .ZN(n390) );
  INV_X1 U452 ( .A(n637), .ZN(n445) );
  AND2_X1 U453 ( .A1(n417), .A2(n416), .ZN(n415) );
  NAND2_X1 U454 ( .A1(n676), .A2(n674), .ZN(n416) );
  NAND2_X1 U455 ( .A1(n409), .A2(n676), .ZN(n417) );
  NAND2_X1 U456 ( .A1(n766), .A2(n357), .ZN(n414) );
  INV_X2 U457 ( .A(n409), .ZN(n766) );
  XNOR2_X1 U458 ( .A(KEYINPUT68), .B(G131), .ZN(n526) );
  AND2_X1 U459 ( .A1(n719), .A2(n720), .ZN(n405) );
  XNOR2_X1 U460 ( .A(G140), .B(KEYINPUT11), .ZN(n498) );
  XNOR2_X1 U461 ( .A(G113), .B(n427), .ZN(n503) );
  XNOR2_X1 U462 ( .A(n504), .B(n526), .ZN(n505) );
  XOR2_X1 U463 ( .A(G104), .B(G122), .Z(n504) );
  XNOR2_X1 U464 ( .A(KEYINPUT5), .B(G137), .ZN(n548) );
  XOR2_X1 U465 ( .A(KEYINPUT90), .B(KEYINPUT77), .Z(n475) );
  XNOR2_X1 U466 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n474) );
  AND2_X1 U467 ( .A1(n631), .A2(n630), .ZN(n668) );
  NAND2_X1 U468 ( .A1(G234), .A2(G237), .ZN(n491) );
  XNOR2_X1 U469 ( .A(n521), .B(n520), .ZN(n522) );
  XOR2_X1 U470 ( .A(G107), .B(G122), .Z(n511) );
  INV_X1 U471 ( .A(G128), .ZN(n478) );
  NOR2_X1 U472 ( .A1(n734), .A2(n736), .ZN(n617) );
  INV_X1 U473 ( .A(KEYINPUT30), .ZN(n436) );
  NAND2_X1 U474 ( .A1(n586), .A2(n462), .ZN(n461) );
  AND2_X1 U475 ( .A1(n473), .A2(n463), .ZN(n462) );
  OR2_X1 U476 ( .A1(n679), .A2(G902), .ZN(n556) );
  INV_X1 U477 ( .A(G478), .ZN(n433) );
  NAND2_X1 U478 ( .A1(n435), .A2(n485), .ZN(n434) );
  XNOR2_X1 U479 ( .A(n509), .B(G475), .ZN(n431) );
  OR2_X1 U480 ( .A1(n675), .A2(G902), .ZN(n432) );
  XNOR2_X1 U481 ( .A(n546), .B(n393), .ZN(n691) );
  XNOR2_X1 U482 ( .A(n527), .B(n359), .ZN(n393) );
  XNOR2_X1 U483 ( .A(n459), .B(n458), .ZN(n768) );
  XNOR2_X1 U484 ( .A(n540), .B(n360), .ZN(n458) );
  XNOR2_X1 U485 ( .A(n771), .B(n538), .ZN(n459) );
  XNOR2_X1 U486 ( .A(n412), .B(n406), .ZN(n761) );
  XNOR2_X1 U487 ( .A(n408), .B(n407), .ZN(n406) );
  XNOR2_X1 U488 ( .A(n364), .B(n528), .ZN(n407) );
  XNOR2_X1 U489 ( .A(n452), .B(KEYINPUT112), .ZN(n782) );
  NAND2_X1 U490 ( .A1(n447), .A2(n446), .ZN(n452) );
  AND2_X1 U491 ( .A1(n448), .A2(n449), .ZN(n447) );
  NOR2_X1 U492 ( .A1(n441), .A2(n390), .ZN(n389) );
  NAND2_X1 U493 ( .A1(n582), .A2(n570), .ZN(n571) );
  NOR2_X1 U494 ( .A1(n453), .A2(n719), .ZN(n570) );
  INV_X1 U495 ( .A(KEYINPUT60), .ZN(n418) );
  INV_X1 U496 ( .A(KEYINPUT56), .ZN(n424) );
  XOR2_X1 U497 ( .A(n530), .B(KEYINPUT108), .Z(n356) );
  AND2_X1 U498 ( .A1(n419), .A2(G475), .ZN(n357) );
  XOR2_X1 U499 ( .A(n526), .B(G134), .Z(n358) );
  NAND2_X1 U500 ( .A1(n442), .A2(n641), .ZN(n441) );
  XOR2_X1 U501 ( .A(KEYINPUT16), .B(G122), .Z(n359) );
  XOR2_X1 U502 ( .A(n537), .B(n536), .Z(n360) );
  AND2_X1 U503 ( .A1(n720), .A2(n456), .ZN(n362) );
  AND2_X1 U504 ( .A1(n453), .A2(n719), .ZN(n363) );
  AND2_X1 U505 ( .A1(G227), .A2(n773), .ZN(n364) );
  NOR2_X1 U506 ( .A1(n719), .A2(n650), .ZN(n365) );
  INV_X1 U507 ( .A(n473), .ZN(n466) );
  XNOR2_X1 U508 ( .A(KEYINPUT109), .B(KEYINPUT33), .ZN(n366) );
  XNOR2_X1 U509 ( .A(KEYINPUT111), .B(KEYINPUT36), .ZN(n367) );
  XOR2_X1 U510 ( .A(n682), .B(n681), .Z(n368) );
  INV_X1 U511 ( .A(n676), .ZN(n419) );
  XNOR2_X1 U512 ( .A(n675), .B(KEYINPUT59), .ZN(n676) );
  XOR2_X1 U513 ( .A(n679), .B(KEYINPUT62), .Z(n369) );
  XOR2_X1 U514 ( .A(KEYINPUT113), .B(KEYINPUT63), .Z(n370) );
  AND2_X1 U515 ( .A1(n677), .A2(G953), .ZN(n770) );
  INV_X1 U516 ( .A(n770), .ZN(n421) );
  INV_X1 U517 ( .A(G475), .ZN(n674) );
  XNOR2_X1 U518 ( .A(n371), .B(n372), .ZN(n762) );
  NAND2_X1 U519 ( .A1(n766), .A2(G469), .ZN(n371) );
  XOR2_X1 U520 ( .A(n761), .B(n760), .Z(n372) );
  XNOR2_X1 U521 ( .A(n662), .B(n661), .ZN(n666) );
  BUF_X1 U522 ( .A(G143), .Z(n427) );
  NAND2_X1 U523 ( .A1(n422), .A2(n421), .ZN(n420) );
  XNOR2_X1 U524 ( .A(n423), .B(n369), .ZN(n422) );
  NAND2_X1 U525 ( .A1(n426), .A2(n421), .ZN(n425) );
  XNOR2_X1 U526 ( .A(n683), .B(n368), .ZN(n426) );
  XNOR2_X1 U527 ( .A(n525), .B(n524), .ZN(n373) );
  XNOR2_X1 U528 ( .A(n525), .B(n524), .ZN(n569) );
  NAND2_X1 U529 ( .A1(n633), .A2(n634), .ZN(n646) );
  NAND2_X1 U530 ( .A1(n382), .A2(n383), .ZN(n375) );
  XNOR2_X1 U531 ( .A(n384), .B(n476), .ZN(n402) );
  NAND2_X2 U532 ( .A1(n388), .A2(n387), .ZN(n785) );
  XNOR2_X2 U533 ( .A(n410), .B(KEYINPUT106), .ZN(n660) );
  INV_X1 U534 ( .A(n785), .ZN(n381) );
  NAND2_X1 U535 ( .A1(n643), .A2(n644), .ZN(n382) );
  NAND2_X1 U536 ( .A1(n648), .A2(n647), .ZN(n383) );
  XNOR2_X1 U537 ( .A(n384), .B(n501), .ZN(n532) );
  XNOR2_X2 U538 ( .A(n403), .B(G146), .ZN(n384) );
  NAND2_X1 U539 ( .A1(n385), .A2(n642), .ZN(n391) );
  NAND2_X1 U540 ( .A1(n443), .A2(n440), .ZN(n385) );
  XNOR2_X1 U541 ( .A(n402), .B(n477), .ZN(n481) );
  NAND2_X1 U542 ( .A1(n386), .A2(n421), .ZN(n413) );
  NAND2_X1 U543 ( .A1(n415), .A2(n414), .ZN(n386) );
  XNOR2_X2 U544 ( .A(n512), .B(n404), .ZN(n480) );
  NAND2_X1 U545 ( .A1(n389), .A2(n443), .ZN(n387) );
  XNOR2_X2 U546 ( .A(n392), .B(n758), .ZN(n573) );
  OR2_X2 U547 ( .A1(n761), .A2(G902), .ZN(n392) );
  XNOR2_X2 U548 ( .A(n394), .B(G110), .ZN(n527) );
  XNOR2_X2 U549 ( .A(G107), .B(G104), .ZN(n394) );
  NAND2_X1 U550 ( .A1(n597), .A2(n397), .ZN(n601) );
  INV_X1 U551 ( .A(n706), .ZN(n397) );
  XNOR2_X2 U552 ( .A(n398), .B(KEYINPUT78), .ZN(n706) );
  NAND2_X1 U553 ( .A1(n399), .A2(n596), .ZN(n398) );
  INV_X1 U554 ( .A(n618), .ZN(n399) );
  XNOR2_X2 U555 ( .A(n400), .B(n366), .ZN(n714) );
  NAND2_X1 U556 ( .A1(n401), .A2(n635), .ZN(n400) );
  XNOR2_X2 U557 ( .A(n556), .B(n555), .ZN(n650) );
  XNOR2_X1 U558 ( .A(n527), .B(n531), .ZN(n408) );
  NAND2_X1 U559 ( .A1(n411), .A2(n363), .ZN(n410) );
  XNOR2_X1 U560 ( .A(n582), .B(KEYINPUT88), .ZN(n411) );
  AND2_X2 U561 ( .A1(n569), .A2(n568), .ZN(n582) );
  XNOR2_X1 U562 ( .A(n412), .B(n553), .ZN(n679) );
  XNOR2_X1 U563 ( .A(n413), .B(n418), .ZN(G60) );
  XNOR2_X1 U564 ( .A(n420), .B(n370), .ZN(G57) );
  NAND2_X1 U565 ( .A1(n680), .A2(G472), .ZN(n423) );
  AND2_X2 U566 ( .A1(n678), .A2(n750), .ZN(n680) );
  XNOR2_X1 U567 ( .A(n425), .B(n424), .ZN(G51) );
  INV_X1 U568 ( .A(n441), .ZN(n440) );
  INV_X1 U569 ( .A(n650), .ZN(n722) );
  NAND2_X2 U570 ( .A1(n523), .A2(n522), .ZN(n525) );
  NAND2_X1 U571 ( .A1(n566), .A2(KEYINPUT19), .ZN(n467) );
  NAND2_X1 U572 ( .A1(n356), .A2(n365), .ZN(n633) );
  INV_X1 U573 ( .A(n602), .ZN(n639) );
  INV_X1 U574 ( .A(n763), .ZN(n435) );
  XNOR2_X1 U575 ( .A(n437), .B(n436), .ZN(n575) );
  NAND2_X1 U576 ( .A1(n650), .A2(n473), .ZN(n437) );
  XNOR2_X1 U577 ( .A(n438), .B(n771), .ZN(n775) );
  NAND2_X1 U578 ( .A1(n637), .A2(KEYINPUT34), .ZN(n442) );
  OR2_X2 U579 ( .A1(n714), .A2(n444), .ZN(n443) );
  NAND2_X1 U580 ( .A1(n445), .A2(n638), .ZN(n444) );
  OR2_X1 U581 ( .A1(n587), .A2(n367), .ZN(n446) );
  NAND2_X1 U582 ( .A1(n587), .A2(n451), .ZN(n448) );
  INV_X1 U583 ( .A(n716), .ZN(n453) );
  NAND2_X1 U584 ( .A1(n455), .A2(n454), .ZN(n564) );
  NAND2_X1 U585 ( .A1(n640), .A2(n602), .ZN(n708) );
  XNOR2_X2 U586 ( .A(G101), .B(KEYINPUT3), .ZN(n468) );
  XNOR2_X2 U587 ( .A(n571), .B(KEYINPUT32), .ZN(n634) );
  XOR2_X1 U588 ( .A(n622), .B(KEYINPUT46), .Z(n471) );
  AND2_X1 U589 ( .A1(G214), .A2(n547), .ZN(n472) );
  NAND2_X1 U590 ( .A1(n490), .A2(G214), .ZN(n473) );
  XNOR2_X1 U591 ( .A(n623), .B(n471), .ZN(n624) );
  INV_X1 U592 ( .A(KEYINPUT10), .ZN(n501) );
  XNOR2_X1 U593 ( .A(n500), .B(n472), .ZN(n502) );
  XNOR2_X1 U594 ( .A(n475), .B(n474), .ZN(n477) );
  NAND2_X1 U595 ( .A1(n773), .A2(G224), .ZN(n476) );
  XNOR2_X2 U596 ( .A(KEYINPUT65), .B(G143), .ZN(n479) );
  XNOR2_X2 U597 ( .A(n479), .B(n478), .ZN(n512) );
  XNOR2_X1 U598 ( .A(n481), .B(n480), .ZN(n483) );
  XNOR2_X1 U599 ( .A(n483), .B(n691), .ZN(n682) );
  XNOR2_X1 U600 ( .A(G902), .B(KEYINPUT15), .ZN(n665) );
  NAND2_X1 U601 ( .A1(n682), .A2(n665), .ZN(n489) );
  INV_X1 U602 ( .A(G902), .ZN(n485) );
  NAND2_X1 U603 ( .A1(n485), .A2(n484), .ZN(n490) );
  NAND2_X1 U604 ( .A1(n490), .A2(G210), .ZN(n487) );
  INV_X1 U605 ( .A(KEYINPUT91), .ZN(n486) );
  XNOR2_X1 U606 ( .A(n491), .B(KEYINPUT14), .ZN(n493) );
  NAND2_X1 U607 ( .A1(n493), .A2(G952), .ZN(n492) );
  XOR2_X1 U608 ( .A(KEYINPUT92), .B(n492), .Z(n744) );
  NAND2_X1 U609 ( .A1(n744), .A2(n773), .ZN(n562) );
  NAND2_X1 U610 ( .A1(n493), .A2(G902), .ZN(n494) );
  XNOR2_X1 U611 ( .A(n494), .B(KEYINPUT93), .ZN(n559) );
  NOR2_X1 U612 ( .A1(G898), .A2(n773), .ZN(n692) );
  NAND2_X1 U613 ( .A1(n559), .A2(n692), .ZN(n495) );
  NAND2_X1 U614 ( .A1(n562), .A2(n495), .ZN(n496) );
  INV_X1 U615 ( .A(n636), .ZN(n523) );
  XOR2_X1 U616 ( .A(KEYINPUT101), .B(KEYINPUT12), .Z(n499) );
  XNOR2_X1 U617 ( .A(n499), .B(n498), .ZN(n500) );
  XOR2_X1 U618 ( .A(n503), .B(KEYINPUT102), .Z(n506) );
  XNOR2_X1 U619 ( .A(n508), .B(n507), .ZN(n675) );
  XNOR2_X1 U620 ( .A(KEYINPUT103), .B(KEYINPUT13), .ZN(n509) );
  XNOR2_X1 U621 ( .A(G116), .B(G134), .ZN(n510) );
  XNOR2_X1 U622 ( .A(n511), .B(n510), .ZN(n513) );
  XNOR2_X1 U623 ( .A(n512), .B(n513), .ZN(n517) );
  NAND2_X1 U624 ( .A1(G217), .A2(n539), .ZN(n515) );
  XOR2_X1 U625 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n514) );
  XNOR2_X1 U626 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U627 ( .A(n517), .B(n516), .ZN(n763) );
  NAND2_X1 U628 ( .A1(n665), .A2(G234), .ZN(n518) );
  XNOR2_X1 U629 ( .A(n518), .B(KEYINPUT20), .ZN(n541) );
  NAND2_X1 U630 ( .A1(n541), .A2(G221), .ZN(n519) );
  XNOR2_X1 U631 ( .A(KEYINPUT21), .B(n519), .ZN(n563) );
  INV_X1 U632 ( .A(KEYINPUT105), .ZN(n520) );
  INV_X1 U633 ( .A(KEYINPUT22), .ZN(n524) );
  XNOR2_X1 U634 ( .A(G101), .B(KEYINPUT95), .ZN(n528) );
  XOR2_X1 U635 ( .A(G137), .B(G140), .Z(n531) );
  INV_X1 U636 ( .A(G469), .ZN(n758) );
  XNOR2_X1 U637 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n529) );
  NAND2_X1 U638 ( .A1(n373), .A2(n453), .ZN(n530) );
  XOR2_X1 U639 ( .A(KEYINPUT76), .B(KEYINPUT82), .Z(n534) );
  XNOR2_X1 U640 ( .A(G119), .B(G110), .ZN(n533) );
  XNOR2_X1 U641 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U642 ( .A(n535), .B(KEYINPUT96), .Z(n538) );
  XOR2_X1 U643 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n537) );
  XNOR2_X1 U644 ( .A(G128), .B(KEYINPUT72), .ZN(n536) );
  NAND2_X1 U645 ( .A1(n539), .A2(G221), .ZN(n540) );
  NAND2_X1 U646 ( .A1(n541), .A2(G217), .ZN(n543) );
  XOR2_X1 U647 ( .A(KEYINPUT97), .B(KEYINPUT25), .Z(n542) );
  XNOR2_X1 U648 ( .A(n543), .B(n542), .ZN(n544) );
  NAND2_X1 U649 ( .A1(n547), .A2(G210), .ZN(n549) );
  XNOR2_X1 U650 ( .A(n549), .B(n548), .ZN(n551) );
  XNOR2_X1 U651 ( .A(KEYINPUT75), .B(KEYINPUT99), .ZN(n550) );
  XNOR2_X1 U652 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U653 ( .A(n546), .B(n552), .ZN(n553) );
  INV_X1 U654 ( .A(KEYINPUT73), .ZN(n554) );
  XNOR2_X1 U655 ( .A(n554), .B(G472), .ZN(n555) );
  XNOR2_X1 U656 ( .A(G110), .B(KEYINPUT116), .ZN(n557) );
  XNOR2_X1 U657 ( .A(n633), .B(n557), .ZN(G12) );
  INV_X1 U658 ( .A(KEYINPUT6), .ZN(n558) );
  INV_X1 U659 ( .A(n635), .ZN(n568) );
  NAND2_X1 U660 ( .A1(G953), .A2(n559), .ZN(n560) );
  OR2_X1 U661 ( .A1(n560), .A2(G900), .ZN(n561) );
  AND2_X1 U662 ( .A1(n562), .A2(n561), .ZN(n574) );
  INV_X1 U663 ( .A(n563), .ZN(n720) );
  NAND2_X1 U664 ( .A1(n453), .A2(n587), .ZN(n565) );
  XNOR2_X1 U665 ( .A(n565), .B(KEYINPUT43), .ZN(n567) );
  INV_X1 U666 ( .A(n586), .ZN(n603) );
  AND2_X1 U667 ( .A1(n567), .A2(n603), .ZN(n629) );
  XOR2_X1 U668 ( .A(n629), .B(G140), .Z(G42) );
  XNOR2_X1 U669 ( .A(n634), .B(G119), .ZN(G21) );
  INV_X1 U670 ( .A(n573), .ZN(n594) );
  NAND2_X1 U671 ( .A1(n717), .A2(n594), .ZN(n654) );
  NOR2_X1 U672 ( .A1(n654), .A2(n574), .ZN(n576) );
  NAND2_X1 U673 ( .A1(n576), .A2(n575), .ZN(n606) );
  INV_X1 U674 ( .A(n606), .ZN(n578) );
  INV_X1 U675 ( .A(KEYINPUT38), .ZN(n577) );
  XNOR2_X1 U676 ( .A(n603), .B(n577), .ZN(n616) );
  OR2_X1 U677 ( .A1(n640), .A2(n602), .ZN(n711) );
  INV_X1 U678 ( .A(n711), .ZN(n580) );
  AND2_X1 U679 ( .A1(n581), .A2(n580), .ZN(n628) );
  XOR2_X1 U680 ( .A(G134), .B(n628), .Z(G36) );
  XNOR2_X1 U681 ( .A(n660), .B(G101), .ZN(G3) );
  INV_X1 U682 ( .A(n708), .ZN(n583) );
  NAND2_X1 U683 ( .A1(n581), .A2(n583), .ZN(n585) );
  INV_X1 U684 ( .A(KEYINPUT40), .ZN(n584) );
  XOR2_X1 U685 ( .A(G131), .B(n621), .Z(G33) );
  XNOR2_X1 U686 ( .A(n782), .B(KEYINPUT87), .ZN(n615) );
  NAND2_X1 U687 ( .A1(n711), .A2(n708), .ZN(n589) );
  INV_X1 U688 ( .A(KEYINPUT104), .ZN(n588) );
  XNOR2_X1 U689 ( .A(n589), .B(n588), .ZN(n737) );
  NOR2_X1 U690 ( .A1(KEYINPUT47), .A2(n737), .ZN(n590) );
  XNOR2_X1 U691 ( .A(n590), .B(KEYINPUT74), .ZN(n591) );
  NOR2_X1 U692 ( .A1(KEYINPUT81), .A2(n591), .ZN(n597) );
  XNOR2_X1 U693 ( .A(n593), .B(KEYINPUT28), .ZN(n595) );
  NAND2_X1 U694 ( .A1(n595), .A2(n594), .ZN(n618) );
  INV_X1 U695 ( .A(KEYINPUT81), .ZN(n598) );
  NAND2_X1 U696 ( .A1(n598), .A2(KEYINPUT47), .ZN(n599) );
  NAND2_X1 U697 ( .A1(n706), .A2(n599), .ZN(n600) );
  NAND2_X1 U698 ( .A1(n601), .A2(n600), .ZN(n613) );
  NOR2_X1 U699 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U700 ( .A1(n640), .A2(n604), .ZN(n605) );
  OR2_X1 U701 ( .A1(n606), .A2(n605), .ZN(n705) );
  NAND2_X1 U702 ( .A1(n737), .A2(KEYINPUT47), .ZN(n607) );
  NAND2_X1 U703 ( .A1(n705), .A2(n607), .ZN(n608) );
  XNOR2_X1 U704 ( .A(n608), .B(KEYINPUT79), .ZN(n611) );
  INV_X1 U705 ( .A(KEYINPUT47), .ZN(n609) );
  NAND2_X1 U706 ( .A1(n609), .A2(KEYINPUT81), .ZN(n610) );
  AND2_X1 U707 ( .A1(n611), .A2(n610), .ZN(n612) );
  NAND2_X1 U708 ( .A1(n613), .A2(n612), .ZN(n614) );
  INV_X1 U709 ( .A(n616), .ZN(n732) );
  NAND2_X1 U710 ( .A1(n732), .A2(n473), .ZN(n736) );
  XNOR2_X1 U711 ( .A(KEYINPUT41), .B(n617), .ZN(n731) );
  NOR2_X1 U712 ( .A1(n731), .A2(n618), .ZN(n620) );
  XNOR2_X1 U713 ( .A(KEYINPUT110), .B(KEYINPUT42), .ZN(n619) );
  XNOR2_X1 U714 ( .A(n620), .B(n619), .ZN(n781) );
  INV_X1 U715 ( .A(KEYINPUT86), .ZN(n622) );
  NAND2_X1 U716 ( .A1(n625), .A2(n624), .ZN(n627) );
  XNOR2_X1 U717 ( .A(KEYINPUT69), .B(KEYINPUT48), .ZN(n626) );
  XNOR2_X1 U718 ( .A(n627), .B(n626), .ZN(n631) );
  NOR2_X1 U719 ( .A1(n629), .A2(n628), .ZN(n630) );
  NAND2_X1 U720 ( .A1(n668), .A2(KEYINPUT2), .ZN(n632) );
  XNOR2_X1 U721 ( .A(n632), .B(KEYINPUT85), .ZN(n664) );
  INV_X1 U722 ( .A(KEYINPUT44), .ZN(n649) );
  BUF_X1 U723 ( .A(n636), .Z(n637) );
  INV_X1 U724 ( .A(KEYINPUT34), .ZN(n638) );
  AND2_X1 U725 ( .A1(n640), .A2(n639), .ZN(n641) );
  INV_X1 U726 ( .A(KEYINPUT35), .ZN(n642) );
  NAND2_X1 U727 ( .A1(n785), .A2(KEYINPUT89), .ZN(n643) );
  NOR2_X1 U728 ( .A1(KEYINPUT89), .A2(KEYINPUT44), .ZN(n645) );
  NAND2_X1 U729 ( .A1(n785), .A2(n645), .ZN(n648) );
  INV_X1 U730 ( .A(n646), .ZN(n647) );
  NAND2_X1 U731 ( .A1(n717), .A2(n650), .ZN(n651) );
  OR2_X1 U732 ( .A1(n651), .A2(n453), .ZN(n727) );
  XNOR2_X1 U733 ( .A(KEYINPUT31), .B(KEYINPUT100), .ZN(n652) );
  XNOR2_X1 U734 ( .A(n653), .B(n652), .ZN(n712) );
  OR2_X1 U735 ( .A1(n637), .A2(n654), .ZN(n656) );
  INV_X1 U736 ( .A(KEYINPUT98), .ZN(n655) );
  XNOR2_X1 U737 ( .A(n656), .B(n655), .ZN(n657) );
  NAND2_X1 U738 ( .A1(n657), .A2(n722), .ZN(n698) );
  INV_X1 U739 ( .A(n737), .ZN(n658) );
  XNOR2_X1 U740 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n661) );
  BUF_X1 U741 ( .A(n666), .Z(n663) );
  NAND2_X1 U742 ( .A1(n664), .A2(n663), .ZN(n750) );
  INV_X1 U743 ( .A(n665), .ZN(n670) );
  NAND2_X1 U744 ( .A1(n666), .A2(n670), .ZN(n667) );
  XNOR2_X1 U745 ( .A(n667), .B(KEYINPUT83), .ZN(n669) );
  NAND2_X1 U746 ( .A1(n669), .A2(n772), .ZN(n672) );
  NAND2_X1 U747 ( .A1(n670), .A2(KEYINPUT2), .ZN(n671) );
  INV_X1 U748 ( .A(G952), .ZN(n677) );
  NAND2_X1 U749 ( .A1(n680), .A2(G210), .ZN(n683) );
  XNOR2_X1 U750 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n681) );
  NAND2_X1 U751 ( .A1(n663), .A2(n773), .ZN(n684) );
  XOR2_X1 U752 ( .A(KEYINPUT125), .B(n684), .Z(n690) );
  XOR2_X1 U753 ( .A(KEYINPUT61), .B(KEYINPUT124), .Z(n686) );
  NAND2_X1 U754 ( .A1(G224), .A2(G953), .ZN(n685) );
  XNOR2_X1 U755 ( .A(n686), .B(n685), .ZN(n687) );
  XNOR2_X1 U756 ( .A(KEYINPUT123), .B(n687), .ZN(n688) );
  NAND2_X1 U757 ( .A1(n688), .A2(G898), .ZN(n689) );
  NAND2_X1 U758 ( .A1(n690), .A2(n689), .ZN(n695) );
  INV_X1 U759 ( .A(n691), .ZN(n693) );
  NOR2_X1 U760 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U761 ( .A(n695), .B(n694), .ZN(G69) );
  NOR2_X1 U762 ( .A1(n698), .A2(n708), .ZN(n696) );
  XOR2_X1 U763 ( .A(KEYINPUT114), .B(n696), .Z(n697) );
  XNOR2_X1 U764 ( .A(G104), .B(n697), .ZN(G6) );
  NOR2_X1 U765 ( .A1(n698), .A2(n711), .ZN(n702) );
  XOR2_X1 U766 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n700) );
  XNOR2_X1 U767 ( .A(G107), .B(KEYINPUT115), .ZN(n699) );
  XNOR2_X1 U768 ( .A(n700), .B(n699), .ZN(n701) );
  XNOR2_X1 U769 ( .A(n702), .B(n701), .ZN(G9) );
  NOR2_X1 U770 ( .A1(n706), .A2(n711), .ZN(n704) );
  XNOR2_X1 U771 ( .A(G128), .B(KEYINPUT29), .ZN(n703) );
  XNOR2_X1 U772 ( .A(n704), .B(n703), .ZN(G30) );
  XNOR2_X1 U773 ( .A(n427), .B(n705), .ZN(G45) );
  NOR2_X1 U774 ( .A1(n706), .A2(n708), .ZN(n707) );
  XOR2_X1 U775 ( .A(G146), .B(n707), .Z(G48) );
  NOR2_X1 U776 ( .A1(n712), .A2(n708), .ZN(n710) );
  XNOR2_X1 U777 ( .A(G113), .B(KEYINPUT117), .ZN(n709) );
  XNOR2_X1 U778 ( .A(n710), .B(n709), .ZN(G15) );
  NOR2_X1 U779 ( .A1(n712), .A2(n711), .ZN(n713) );
  XOR2_X1 U780 ( .A(G116), .B(n713), .Z(G18) );
  BUF_X1 U781 ( .A(n714), .Z(n715) );
  OR2_X1 U782 ( .A1(n731), .A2(n715), .ZN(n747) );
  NOR2_X1 U783 ( .A1(n717), .A2(n355), .ZN(n718) );
  XNOR2_X1 U784 ( .A(n718), .B(KEYINPUT50), .ZN(n725) );
  NOR2_X1 U785 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U786 ( .A(n721), .B(KEYINPUT49), .ZN(n723) );
  NAND2_X1 U787 ( .A1(n723), .A2(n722), .ZN(n724) );
  NOR2_X1 U788 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U789 ( .A(n726), .B(KEYINPUT119), .ZN(n728) );
  NAND2_X1 U790 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U791 ( .A(KEYINPUT51), .B(n729), .ZN(n730) );
  NOR2_X1 U792 ( .A1(n731), .A2(n730), .ZN(n742) );
  NOR2_X1 U793 ( .A1(n732), .A2(n473), .ZN(n733) );
  NOR2_X1 U794 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U795 ( .A(n735), .B(KEYINPUT120), .ZN(n739) );
  NOR2_X1 U796 ( .A1(n737), .A2(n736), .ZN(n738) );
  NOR2_X1 U797 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X1 U798 ( .A1(n740), .A2(n715), .ZN(n741) );
  NOR2_X1 U799 ( .A1(n742), .A2(n741), .ZN(n743) );
  XOR2_X1 U800 ( .A(KEYINPUT52), .B(n743), .Z(n745) );
  NAND2_X1 U801 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U802 ( .A1(n747), .A2(n746), .ZN(n754) );
  AND2_X1 U803 ( .A1(n772), .A2(n663), .ZN(n749) );
  XNOR2_X1 U804 ( .A(KEYINPUT80), .B(KEYINPUT2), .ZN(n748) );
  NOR2_X1 U805 ( .A1(n749), .A2(n748), .ZN(n752) );
  INV_X1 U806 ( .A(n750), .ZN(n751) );
  NOR2_X1 U807 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U808 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U809 ( .A(n755), .B(KEYINPUT121), .ZN(n756) );
  NOR2_X1 U810 ( .A1(G953), .A2(n756), .ZN(n757) );
  XNOR2_X1 U811 ( .A(KEYINPUT53), .B(n757), .ZN(G75) );
  XNOR2_X1 U812 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n759) );
  XNOR2_X1 U813 ( .A(n759), .B(KEYINPUT57), .ZN(n760) );
  NOR2_X1 U814 ( .A1(n770), .A2(n762), .ZN(G54) );
  NAND2_X1 U815 ( .A1(n766), .A2(G478), .ZN(n764) );
  XNOR2_X1 U816 ( .A(n764), .B(n763), .ZN(n765) );
  NOR2_X1 U817 ( .A1(n770), .A2(n765), .ZN(G63) );
  NAND2_X1 U818 ( .A1(n766), .A2(G217), .ZN(n767) );
  XNOR2_X1 U819 ( .A(n768), .B(n767), .ZN(n769) );
  NOR2_X1 U820 ( .A1(n770), .A2(n769), .ZN(G66) );
  XNOR2_X1 U821 ( .A(n772), .B(n775), .ZN(n774) );
  NAND2_X1 U822 ( .A1(n774), .A2(n773), .ZN(n780) );
  XOR2_X1 U823 ( .A(n775), .B(G227), .Z(n776) );
  NAND2_X1 U824 ( .A1(n776), .A2(G900), .ZN(n777) );
  XNOR2_X1 U825 ( .A(KEYINPUT126), .B(n777), .ZN(n778) );
  NAND2_X1 U826 ( .A1(n778), .A2(G953), .ZN(n779) );
  NAND2_X1 U827 ( .A1(n780), .A2(n779), .ZN(G72) );
  XOR2_X1 U828 ( .A(G137), .B(n781), .Z(G39) );
  XOR2_X1 U829 ( .A(KEYINPUT37), .B(KEYINPUT118), .Z(n784) );
  XNOR2_X1 U830 ( .A(G125), .B(n782), .ZN(n783) );
  XNOR2_X1 U831 ( .A(n784), .B(n783), .ZN(G27) );
  BUF_X1 U832 ( .A(n785), .Z(n786) );
  XNOR2_X1 U833 ( .A(G122), .B(n786), .ZN(G24) );
endmodule

