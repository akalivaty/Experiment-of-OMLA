//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 1 1 0 1 0 0 1 0 1 1 1 0 1 0 1 1 0 1 0 1 0 1 0 1 0 1 0 1 1 1 0 1 0 0 1 1 1 0 1 0 1 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:00 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1286, new_n1287, new_n1288, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  OAI21_X1  g0012(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NOR3_X1   g0014(.A1(KEYINPUT64), .A2(G58), .A3(G68), .ZN(new_n215));
  OAI21_X1  g0015(.A(G50), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT65), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(new_n207), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT67), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT66), .Z(new_n227));
  OAI21_X1  g0027(.A(new_n209), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n212), .B(new_n220), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(KEYINPUT68), .Z(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G226), .ZN(new_n234));
  INV_X1    g0034(.A(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G250), .B(G257), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT69), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n236), .B(new_n240), .Z(G358));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(KEYINPUT77), .ZN(new_n249));
  OR2_X1    g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G1698), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n252), .A2(G226), .A3(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n252), .A2(G232), .A3(G1698), .ZN(new_n255));
  AND3_X1   g0055(.A1(KEYINPUT75), .A2(G33), .A3(G97), .ZN(new_n256));
  AOI21_X1  g0056(.A(KEYINPUT75), .B1(G33), .B2(G97), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n254), .A2(new_n255), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G33), .A2(G41), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n260), .A2(G1), .A3(G13), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n264));
  INV_X1    g0064(.A(G274), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n261), .A2(new_n264), .ZN(new_n268));
  INV_X1    g0068(.A(G238), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n263), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n272), .A2(KEYINPUT76), .A3(KEYINPUT13), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT76), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n270), .B1(new_n259), .B2(new_n262), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT13), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n275), .A2(new_n276), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n273), .A2(new_n277), .A3(G190), .A4(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  AOI211_X1 g0080(.A(KEYINPUT13), .B(new_n270), .C1(new_n262), .C2(new_n259), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n276), .B1(new_n263), .B2(new_n271), .ZN(new_n282));
  OAI21_X1  g0082(.A(G200), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(new_n218), .ZN(new_n287));
  OAI21_X1  g0087(.A(KEYINPUT72), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT72), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n284), .A2(new_n289), .A3(new_n218), .A4(new_n286), .ZN(new_n290));
  AND2_X1   g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n206), .A2(G20), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n291), .A2(G68), .A3(new_n292), .ZN(new_n293));
  NOR2_X1   g0093(.A1(G20), .A2(G33), .ZN(new_n294));
  INV_X1    g0094(.A(G68), .ZN(new_n295));
  AOI22_X1  g0095(.A1(new_n294), .A2(G50), .B1(G20), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G77), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n207), .A2(G33), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n296), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n299), .A2(KEYINPUT11), .A3(new_n287), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n287), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT11), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G13), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n304), .A2(G1), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n305), .A2(G20), .A3(new_n295), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n306), .B(KEYINPUT12), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n293), .A2(new_n300), .A3(new_n303), .A4(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n283), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n249), .B1(new_n280), .B2(new_n310), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n279), .A2(KEYINPUT77), .A3(new_n283), .A4(new_n309), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g0113(.A(G169), .B1(new_n281), .B2(new_n282), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n314), .A2(KEYINPUT78), .A3(KEYINPUT14), .ZN(new_n315));
  NAND2_X1  g0115(.A1(KEYINPUT78), .A2(KEYINPUT14), .ZN(new_n316));
  OAI211_X1 g0116(.A(G169), .B(new_n316), .C1(new_n281), .C2(new_n282), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n273), .A2(new_n277), .A3(G179), .A4(new_n278), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n315), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(new_n308), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n313), .A2(new_n320), .ZN(new_n321));
  MUX2_X1   g0121(.A(G222), .B(G223), .S(G1698), .Z(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n252), .ZN(new_n323));
  AND2_X1   g0123(.A1(KEYINPUT3), .A2(G33), .ZN(new_n324));
  NOR2_X1   g0124(.A1(KEYINPUT3), .A2(G33), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(G77), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n261), .B1(new_n323), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G226), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n267), .B1(new_n268), .B2(new_n329), .ZN(new_n330));
  OR2_X1    g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g0131(.A(KEYINPUT73), .B(G200), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G190), .ZN(new_n335));
  OR3_X1    g0135(.A1(new_n328), .A2(new_n330), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n285), .A2(new_n287), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n339), .A2(G50), .A3(new_n292), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n340), .B1(G50), .B2(new_n284), .ZN(new_n341));
  INV_X1    g0141(.A(new_n287), .ZN(new_n342));
  XNOR2_X1  g0142(.A(KEYINPUT8), .B(G58), .ZN(new_n343));
  OR2_X1    g0143(.A1(new_n343), .A2(new_n298), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n294), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n342), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n341), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(KEYINPUT9), .ZN(new_n348));
  OR2_X1    g0148(.A1(new_n347), .A2(KEYINPUT9), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n338), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT10), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT74), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n350), .B(new_n351), .C1(new_n352), .C2(new_n337), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n351), .B1(new_n337), .B2(new_n352), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n354), .A2(new_n338), .A3(new_n348), .A4(new_n349), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n331), .A2(G169), .ZN(new_n356));
  INV_X1    g0156(.A(G179), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n356), .B1(new_n357), .B2(new_n331), .ZN(new_n358));
  INV_X1    g0158(.A(new_n347), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n353), .A2(new_n355), .A3(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n291), .A2(G77), .A3(new_n292), .ZN(new_n362));
  INV_X1    g0162(.A(new_n294), .ZN(new_n363));
  OR2_X1    g0163(.A1(new_n363), .A2(KEYINPUT70), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(KEYINPUT70), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n343), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  XNOR2_X1  g0166(.A(KEYINPUT15), .B(G87), .ZN(new_n367));
  OAI22_X1  g0167(.A1(new_n367), .A2(new_n298), .B1(new_n207), .B2(new_n297), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n287), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n284), .A2(G77), .ZN(new_n370));
  XNOR2_X1  g0170(.A(new_n370), .B(KEYINPUT71), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n362), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n252), .A2(G238), .A3(G1698), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n252), .A2(G232), .A3(new_n253), .ZN(new_n375));
  INV_X1    g0175(.A(G107), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n374), .B(new_n375), .C1(new_n376), .C2(new_n252), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n262), .ZN(new_n378));
  INV_X1    g0178(.A(new_n268), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n266), .B1(new_n379), .B2(G244), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n381), .A2(G190), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n333), .B1(new_n378), .B2(new_n380), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n373), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n381), .A2(new_n357), .ZN(new_n385));
  INV_X1    g0185(.A(G169), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n386), .B1(new_n378), .B2(new_n380), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n372), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n384), .A2(new_n388), .ZN(new_n389));
  NOR3_X1   g0189(.A1(new_n321), .A2(new_n361), .A3(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT80), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n250), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n251), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT79), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NOR3_X1   g0194(.A1(new_n324), .A2(new_n325), .A3(G20), .ZN(new_n395));
  OAI21_X1  g0195(.A(KEYINPUT79), .B1(new_n395), .B2(KEYINPUT7), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n394), .B1(new_n396), .B2(new_n392), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n391), .B1(new_n397), .B2(new_n295), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n250), .A2(new_n207), .A3(new_n251), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT7), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n393), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n392), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  OAI211_X1 g0203(.A(KEYINPUT80), .B(G68), .C1(new_n403), .C2(new_n394), .ZN(new_n404));
  XNOR2_X1  g0204(.A(G58), .B(G68), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n405), .A2(G20), .B1(G159), .B2(new_n294), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n398), .A2(KEYINPUT16), .A3(new_n404), .A4(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(KEYINPUT7), .B1(new_n326), .B2(new_n207), .ZN(new_n408));
  OAI21_X1  g0208(.A(G68), .B1(new_n408), .B2(new_n402), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(new_n406), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT16), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n342), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n407), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n339), .ZN(new_n414));
  INV_X1    g0214(.A(new_n343), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n292), .ZN(new_n416));
  OAI22_X1  g0216(.A1(new_n414), .A2(new_n416), .B1(new_n284), .B2(new_n415), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n266), .B1(new_n379), .B2(G232), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n252), .A2(G226), .A3(G1698), .ZN(new_n419));
  INV_X1    g0219(.A(G33), .ZN(new_n420));
  INV_X1    g0220(.A(G87), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n419), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT81), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n253), .A2(G223), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n425), .B1(new_n326), .B2(new_n426), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n252), .A2(KEYINPUT81), .A3(G223), .A4(new_n253), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n424), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n335), .B(new_n418), .C1(new_n429), .C2(new_n261), .ZN(new_n430));
  INV_X1    g0230(.A(G200), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n326), .A2(new_n329), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n422), .B1(new_n432), .B2(G1698), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n428), .A2(new_n427), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n261), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n418), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n431), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n417), .B1(new_n430), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n413), .A2(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n439), .A2(KEYINPUT17), .ZN(new_n440));
  AND3_X1   g0240(.A1(new_n413), .A2(new_n438), .A3(KEYINPUT82), .ZN(new_n441));
  AOI21_X1  g0241(.A(KEYINPUT82), .B1(new_n413), .B2(new_n438), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n440), .B1(new_n443), .B2(KEYINPUT17), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n357), .B(new_n418), .C1(new_n429), .C2(new_n261), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n386), .B1(new_n435), .B2(new_n436), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n417), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n447), .B1(new_n413), .B2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT18), .ZN(new_n450));
  XNOR2_X1  g0250(.A(new_n449), .B(new_n450), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n444), .A2(new_n451), .ZN(new_n452));
  AND2_X1   g0252(.A1(new_n390), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n206), .A2(G33), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n288), .A2(new_n290), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(G116), .ZN(new_n456));
  INV_X1    g0256(.A(G116), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n284), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n286), .A2(new_n218), .B1(G20), .B2(new_n457), .ZN(new_n460));
  AOI21_X1  g0260(.A(G20), .B1(G33), .B2(G283), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n420), .A2(G97), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT88), .ZN(new_n463));
  AND3_X1   g0263(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n463), .B1(new_n461), .B2(new_n462), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n460), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT20), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI211_X1 g0268(.A(KEYINPUT20), .B(new_n460), .C1(new_n464), .C2(new_n465), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n459), .A2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT5), .ZN(new_n472));
  OAI21_X1  g0272(.A(G274), .B1(new_n472), .B2(G41), .ZN(new_n473));
  INV_X1    g0273(.A(new_n218), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n473), .B1(new_n474), .B2(new_n260), .ZN(new_n475));
  INV_X1    g0275(.A(G41), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n206), .B(G45), .C1(new_n476), .C2(KEYINPUT5), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n477), .A2(KEYINPUT84), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT84), .ZN(new_n479));
  INV_X1    g0279(.A(G45), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n480), .A2(G1), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n472), .A2(G41), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n479), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n475), .B1(new_n478), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n472), .A2(G41), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n261), .B(G270), .C1(new_n477), .C2(new_n485), .ZN(new_n486));
  AND2_X1   g0286(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  OAI211_X1 g0287(.A(G264), .B(G1698), .C1(new_n324), .C2(new_n325), .ZN(new_n488));
  OAI211_X1 g0288(.A(G257), .B(new_n253), .C1(new_n324), .C2(new_n325), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n250), .A2(G303), .A3(new_n251), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n262), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n386), .B1(new_n487), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n471), .A2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT21), .ZN(new_n495));
  OAI21_X1  g0295(.A(KEYINPUT89), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n456), .A2(new_n458), .B1(new_n468), .B2(new_n469), .ZN(new_n497));
  AND2_X1   g0297(.A1(new_n491), .A2(new_n262), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n484), .A2(new_n486), .ZN(new_n499));
  OAI21_X1  g0299(.A(G169), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT89), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n501), .A2(new_n502), .A3(KEYINPUT21), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n496), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n498), .A2(new_n499), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n335), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n506), .B1(G200), .B2(new_n505), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n497), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n492), .A2(G179), .A3(new_n484), .A4(new_n486), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n509), .B1(new_n459), .B2(new_n470), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n510), .B1(new_n494), .B2(new_n495), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n504), .A2(new_n508), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n305), .A2(G20), .A3(new_n376), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(KEYINPUT25), .ZN(new_n514));
  OR2_X1    g0314(.A1(new_n513), .A2(KEYINPUT25), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n339), .A2(new_n454), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n514), .B(new_n515), .C1(new_n516), .C2(new_n376), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT23), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n519), .B1(new_n207), .B2(G107), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n376), .A2(KEYINPUT23), .A3(G20), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n420), .A2(new_n457), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n207), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT22), .ZN(new_n527));
  AOI21_X1  g0327(.A(G20), .B1(new_n250), .B2(new_n251), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n527), .B1(new_n528), .B2(G87), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n207), .B(G87), .C1(new_n324), .C2(new_n325), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n530), .A2(KEYINPUT22), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n526), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT24), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n287), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n528), .A2(new_n527), .A3(G87), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n530), .A2(KEYINPUT22), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n525), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n537), .A2(KEYINPUT24), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n518), .B1(new_n534), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(KEYINPUT90), .ZN(new_n540));
  OAI211_X1 g0340(.A(G250), .B(new_n253), .C1(new_n324), .C2(new_n325), .ZN(new_n541));
  OAI211_X1 g0341(.A(G257), .B(G1698), .C1(new_n324), .C2(new_n325), .ZN(new_n542));
  NAND2_X1  g0342(.A1(G33), .A2(G294), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n261), .B1(new_n477), .B2(new_n485), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n262), .A2(new_n544), .B1(new_n546), .B2(G264), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n547), .A2(KEYINPUT91), .A3(G179), .A4(new_n484), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT91), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n544), .A2(new_n262), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n261), .B(G264), .C1(new_n477), .C2(new_n485), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n550), .A2(new_n484), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n549), .B1(new_n552), .B2(G169), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n552), .A2(new_n357), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n548), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n342), .B1(new_n537), .B2(KEYINPUT24), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n532), .A2(new_n533), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n517), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT90), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n540), .A2(new_n555), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n552), .A2(new_n431), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n562), .B1(G190), .B2(new_n552), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n558), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n516), .ZN(new_n566));
  INV_X1    g0366(.A(G97), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n285), .A2(G97), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(G107), .B1(new_n408), .B2(new_n402), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT6), .ZN(new_n572));
  AND2_X1   g0372(.A1(G97), .A2(G107), .ZN(new_n573));
  NOR2_X1   g0373(.A1(G97), .A2(G107), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n376), .A2(KEYINPUT6), .A3(G97), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n577), .A2(G20), .B1(G77), .B2(new_n294), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n571), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n287), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT83), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n342), .B1(new_n571), .B2(new_n578), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(KEYINPUT83), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n570), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n252), .A2(G244), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT4), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(G33), .A2(G283), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n252), .A2(KEYINPUT4), .A3(G244), .A4(new_n253), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n252), .A2(G250), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n253), .B1(new_n592), .B2(KEYINPUT4), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n262), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n546), .A2(G257), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n484), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n594), .A2(new_n597), .A3(new_n335), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n586), .A2(new_n587), .B1(G33), .B2(G283), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n587), .B1(new_n252), .B2(G250), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n599), .B(new_n590), .C1(new_n253), .C2(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n596), .B1(new_n601), .B2(new_n262), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n598), .B1(new_n602), .B2(G200), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n585), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n583), .A2(KEYINPUT83), .ZN(new_n605));
  AOI211_X1 g0405(.A(new_n581), .B(new_n342), .C1(new_n571), .C2(new_n578), .ZN(new_n606));
  OAI22_X1  g0406(.A1(new_n605), .A2(new_n606), .B1(new_n569), .B2(new_n568), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n594), .A2(new_n597), .A3(G179), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n608), .B1(new_n602), .B2(new_n386), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n604), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n252), .A2(new_n207), .ZN(new_n612));
  NAND2_X1  g0412(.A1(G33), .A2(G97), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n613), .A2(G20), .ZN(new_n614));
  OAI22_X1  g0414(.A1(new_n612), .A2(new_n295), .B1(KEYINPUT19), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(KEYINPUT19), .B1(new_n256), .B2(new_n257), .ZN(new_n616));
  NOR2_X1   g0416(.A1(G87), .A2(G97), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n616), .A2(new_n207), .B1(new_n376), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n287), .B1(new_n615), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n367), .A2(new_n285), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n619), .B(new_n620), .C1(new_n421), .C2(new_n516), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n481), .A2(G274), .ZN(new_n622));
  OAI21_X1  g0422(.A(G250), .B1(new_n480), .B2(G1), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n262), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  OAI211_X1 g0424(.A(G244), .B(G1698), .C1(new_n324), .C2(new_n325), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT85), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n252), .A2(KEYINPUT85), .A3(G244), .A4(G1698), .ZN(new_n628));
  INV_X1    g0428(.A(new_n523), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n252), .A2(G238), .A3(new_n253), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n627), .A2(new_n628), .A3(new_n629), .A4(new_n630), .ZN(new_n631));
  AOI211_X1 g0431(.A(new_n335), .B(new_n624), .C1(new_n631), .C2(new_n262), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n621), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n624), .B1(new_n631), .B2(new_n262), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n333), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n634), .A2(new_n357), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(KEYINPUT86), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n635), .A2(new_n386), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n367), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n566), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n619), .A2(new_n620), .A3(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT87), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT86), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n634), .A2(new_n647), .A3(new_n357), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n619), .A2(new_n643), .A3(KEYINPUT87), .A4(new_n620), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n646), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n637), .B1(new_n641), .B2(new_n650), .ZN(new_n651));
  NOR4_X1   g0451(.A1(new_n512), .A2(new_n565), .A3(new_n611), .A4(new_n651), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n453), .A2(new_n652), .ZN(G372));
  XNOR2_X1  g0453(.A(new_n449), .B(KEYINPUT18), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n388), .B1(new_n311), .B2(new_n312), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n655), .B1(new_n308), .B2(new_n319), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n654), .B1(new_n656), .B2(new_n444), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n355), .A2(new_n353), .ZN(new_n658));
  AOI22_X1  g0458(.A1(new_n657), .A2(new_n658), .B1(new_n359), .B2(new_n358), .ZN(new_n659));
  INV_X1    g0459(.A(new_n453), .ZN(new_n660));
  INV_X1    g0460(.A(new_n651), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT26), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n610), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g0464(.A(new_n624), .B(KEYINPUT92), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n631), .A2(new_n262), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n333), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n633), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n604), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n555), .A2(new_n539), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n502), .B1(new_n501), .B2(KEYINPUT21), .ZN(new_n672));
  NOR4_X1   g0472(.A1(new_n497), .A2(new_n500), .A3(KEYINPUT89), .A4(new_n495), .ZN(new_n673));
  OAI211_X1 g0473(.A(new_n671), .B(new_n511), .C1(new_n672), .C2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(new_n564), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n670), .B1(new_n675), .B2(new_n610), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n664), .B1(new_n676), .B2(KEYINPUT26), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n667), .A2(new_n386), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n678), .A2(new_n638), .A3(new_n644), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n659), .B1(new_n660), .B2(new_n680), .ZN(G369));
  INV_X1    g0481(.A(new_n305), .ZN(new_n682));
  OR3_X1    g0482(.A1(new_n682), .A2(KEYINPUT27), .A3(G20), .ZN(new_n683));
  OAI21_X1  g0483(.A(KEYINPUT27), .B1(new_n682), .B2(G20), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(G213), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(G343), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n497), .A2(new_n688), .ZN(new_n689));
  OAI22_X1  g0489(.A1(new_n501), .A2(KEYINPUT21), .B1(new_n497), .B2(new_n509), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n690), .B1(new_n503), .B2(new_n496), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n689), .B1(new_n691), .B2(new_n508), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n692), .B1(new_n691), .B2(new_n689), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(G330), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n561), .A2(new_n688), .ZN(new_n695));
  INV_X1    g0495(.A(new_n565), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n540), .A2(new_n560), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n697), .A2(KEYINPUT93), .A3(new_n687), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n697), .A2(new_n687), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT93), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n695), .B1(new_n699), .B2(new_n702), .ZN(new_n703));
  OR3_X1    g0503(.A1(new_n694), .A2(KEYINPUT94), .A3(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(KEYINPUT94), .B1(new_n694), .B2(new_n703), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n691), .A2(new_n687), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n707), .A2(new_n702), .A3(new_n696), .A4(new_n698), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n555), .A2(new_n539), .A3(new_n688), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n706), .A2(new_n711), .ZN(G399));
  INV_X1    g0512(.A(KEYINPUT95), .ZN(new_n713));
  INV_X1    g0513(.A(new_n210), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n713), .B1(new_n714), .B2(G41), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n210), .A2(KEYINPUT95), .A3(new_n476), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n617), .A2(new_n376), .A3(new_n457), .ZN(new_n719));
  NOR3_X1   g0519(.A1(new_n718), .A2(new_n206), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n720), .B1(new_n217), .B2(new_n718), .ZN(new_n721));
  XOR2_X1   g0521(.A(new_n721), .B(KEYINPUT28), .Z(new_n722));
  NOR3_X1   g0522(.A1(new_n565), .A2(new_n611), .A3(new_n651), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n723), .A2(new_n691), .A3(new_n508), .A4(new_n688), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT30), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n602), .A2(new_n547), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n505), .A2(G179), .A3(new_n634), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n635), .A2(new_n509), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n729), .A2(KEYINPUT30), .A3(new_n602), .A4(new_n547), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n505), .A2(G179), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n594), .A2(new_n597), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n731), .A2(new_n732), .A3(new_n552), .A4(new_n667), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n728), .A2(new_n730), .A3(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n734), .A2(KEYINPUT31), .A3(new_n687), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(KEYINPUT31), .B1(new_n734), .B2(new_n687), .ZN(new_n737));
  OAI21_X1  g0537(.A(KEYINPUT96), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n734), .A2(new_n687), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT31), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT96), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n741), .A2(new_n742), .A3(new_n735), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n724), .A2(new_n738), .A3(new_n743), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n744), .A2(G330), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n687), .B1(new_n677), .B2(new_n679), .ZN(new_n746));
  OR2_X1    g0546(.A1(new_n746), .A2(KEYINPUT29), .ZN(new_n747));
  INV_X1    g0547(.A(new_n679), .ZN(new_n748));
  AOI22_X1  g0548(.A1(new_n633), .A2(new_n668), .B1(new_n563), .B2(new_n558), .ZN(new_n749));
  AND3_X1   g0549(.A1(new_n749), .A2(new_n604), .A3(new_n610), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n504), .A2(new_n511), .A3(new_n561), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n748), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n662), .B1(new_n651), .B2(new_n610), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n663), .A2(new_n669), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n687), .B1(new_n752), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(KEYINPUT29), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n745), .B1(new_n747), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n722), .B1(new_n758), .B2(G1), .ZN(G364));
  NOR2_X1   g0559(.A1(new_n304), .A2(G20), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(G45), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n717), .A2(G1), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n694), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n693), .A2(G330), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G13), .A2(G33), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(G20), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n693), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n762), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n210), .A2(new_n252), .ZN(new_n771));
  XNOR2_X1  g0571(.A(G355), .B(KEYINPUT97), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n771), .A2(new_n772), .B1(G116), .B2(new_n210), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n244), .A2(G45), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n774), .B1(new_n217), .B2(G45), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n714), .A2(new_n252), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n773), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n218), .B1(G20), .B2(new_n386), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n767), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n770), .B1(new_n777), .B2(new_n780), .ZN(new_n781));
  OR2_X1    g0581(.A1(new_n781), .A2(KEYINPUT98), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n357), .A2(new_n431), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n207), .A2(new_n335), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n357), .A2(G200), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(G58), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n785), .A2(new_n202), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(G179), .A2(G200), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G190), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G20), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G97), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n207), .A2(G190), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(new_n786), .ZN(new_n795));
  OAI211_X1 g0595(.A(new_n793), .B(new_n252), .C1(new_n297), .C2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n783), .A2(new_n794), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI211_X1 g0598(.A(new_n789), .B(new_n796), .C1(G68), .C2(new_n798), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n333), .A2(new_n357), .A3(new_n784), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(G87), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n794), .A2(new_n790), .ZN(new_n803));
  INV_X1    g0603(.A(G159), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT32), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n333), .A2(new_n357), .A3(new_n794), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(G107), .ZN(new_n809));
  NAND4_X1  g0609(.A1(new_n799), .A2(new_n802), .A3(new_n806), .A4(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n803), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n808), .A2(G283), .B1(G329), .B2(new_n811), .ZN(new_n812));
  XOR2_X1   g0612(.A(new_n812), .B(KEYINPUT100), .Z(new_n813));
  NOR2_X1   g0613(.A1(KEYINPUT33), .A2(G317), .ZN(new_n814));
  AND2_X1   g0614(.A1(KEYINPUT33), .A2(G317), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n798), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(G311), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n816), .B1(new_n817), .B2(new_n795), .ZN(new_n818));
  INV_X1    g0618(.A(new_n787), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n818), .B1(G322), .B2(new_n819), .ZN(new_n820));
  XNOR2_X1  g0620(.A(KEYINPUT99), .B(G326), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n326), .B1(new_n785), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(G294), .B2(new_n792), .ZN(new_n823));
  INV_X1    g0623(.A(G303), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n820), .B(new_n823), .C1(new_n824), .C2(new_n800), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n810), .B1(new_n813), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(new_n778), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n781), .A2(KEYINPUT98), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n782), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n763), .A2(new_n764), .B1(new_n769), .B2(new_n829), .ZN(G396));
  INV_X1    g0630(.A(G132), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n252), .B1(new_n803), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n832), .B1(G58), .B2(new_n792), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n833), .B1(new_n295), .B2(new_n807), .ZN(new_n834));
  INV_X1    g0634(.A(new_n785), .ZN(new_n835));
  INV_X1    g0635(.A(new_n795), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n835), .A2(G137), .B1(new_n836), .B2(G159), .ZN(new_n837));
  INV_X1    g0637(.A(G143), .ZN(new_n838));
  INV_X1    g0638(.A(G150), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n837), .B1(new_n838), .B2(new_n787), .C1(new_n839), .C2(new_n797), .ZN(new_n840));
  XOR2_X1   g0640(.A(new_n840), .B(KEYINPUT34), .Z(new_n841));
  AOI211_X1 g0641(.A(new_n834), .B(new_n841), .C1(G50), .C2(new_n801), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n808), .A2(G87), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n797), .A2(KEYINPUT101), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n797), .A2(KEYINPUT101), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(G283), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n843), .B1(new_n376), .B2(new_n800), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n835), .A2(G303), .B1(new_n836), .B2(G116), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(new_n817), .B2(new_n803), .ZN(new_n850));
  INV_X1    g0650(.A(G294), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n793), .B(new_n326), .C1(new_n851), .C2(new_n787), .ZN(new_n852));
  NOR3_X1   g0652(.A1(new_n848), .A2(new_n850), .A3(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n778), .B1(new_n842), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n778), .A2(new_n765), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n762), .B1(new_n297), .B2(new_n855), .ZN(new_n856));
  OR2_X1    g0656(.A1(new_n388), .A2(new_n688), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT102), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n372), .A2(new_n687), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n384), .A2(new_n388), .A3(new_n859), .A4(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n384), .A2(new_n388), .A3(new_n860), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(KEYINPUT102), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n858), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n854), .B(new_n856), .C1(new_n865), .C2(new_n766), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n746), .B(new_n864), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n745), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(new_n762), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n867), .A2(new_n745), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n866), .B1(new_n869), .B2(new_n870), .ZN(G384));
  NAND2_X1  g0671(.A1(new_n413), .A2(new_n448), .ZN(new_n872));
  INV_X1    g0672(.A(new_n447), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n685), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT37), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n874), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT82), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n439), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n413), .A2(new_n438), .A3(KEYINPUT82), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n878), .A2(new_n882), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n404), .A2(new_n406), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT16), .B1(new_n884), .B2(new_n398), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n407), .A2(new_n287), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n448), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n447), .A2(new_n685), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n877), .B1(new_n443), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(KEYINPUT103), .B1(new_n883), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n398), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n404), .A2(new_n406), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n411), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n894), .A2(new_n407), .A3(new_n287), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n685), .B1(new_n895), .B2(new_n448), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n896), .B1(new_n444), .B2(new_n451), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n895), .A2(new_n448), .B1(new_n447), .B2(new_n685), .ZN(new_n898));
  OAI21_X1  g0698(.A(KEYINPUT37), .B1(new_n882), .B2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n449), .A2(KEYINPUT37), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n443), .A2(new_n900), .A3(new_n876), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT103), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n899), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n891), .A2(new_n897), .A3(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT38), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n891), .A2(new_n897), .A3(new_n903), .A4(KEYINPUT38), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n741), .A2(new_n735), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n910), .B1(new_n652), .B2(new_n688), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n309), .A2(new_n688), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n313), .A2(new_n320), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n913), .B1(new_n313), .B2(new_n320), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n865), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT105), .B1(new_n911), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n724), .A2(new_n741), .A3(new_n735), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n321), .A2(new_n912), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n313), .A2(new_n320), .A3(new_n913), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n864), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(KEYINPUT105), .A2(KEYINPUT40), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n918), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  AND2_X1   g0723(.A1(new_n917), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n918), .A2(new_n921), .ZN(new_n925));
  OAI21_X1  g0725(.A(KEYINPUT104), .B1(new_n878), .B2(new_n882), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT104), .ZN(new_n927));
  NAND4_X1  g0727(.A1(new_n443), .A2(new_n900), .A3(new_n927), .A4(new_n876), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n874), .A2(new_n876), .A3(new_n439), .ZN(new_n929));
  AOI22_X1  g0729(.A1(new_n926), .A2(new_n928), .B1(KEYINPUT37), .B2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n440), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT17), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n931), .B1(new_n882), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n876), .B1(new_n933), .B2(new_n654), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n905), .B1(new_n930), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n925), .B1(new_n935), .B2(new_n907), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT40), .ZN(new_n937));
  OAI22_X1  g0737(.A1(new_n909), .A2(new_n924), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n453), .A2(new_n918), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n938), .B(new_n939), .Z(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(G330), .ZN(new_n941));
  XOR2_X1   g0741(.A(new_n941), .B(KEYINPUT106), .Z(new_n942));
  NAND2_X1  g0742(.A1(new_n746), .A2(new_n865), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n388), .A2(new_n687), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n914), .A2(new_n915), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n945), .A2(new_n947), .A3(new_n908), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT39), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n949), .B1(new_n906), .B2(new_n907), .ZN(new_n950));
  AND3_X1   g0750(.A1(new_n935), .A2(new_n949), .A3(new_n907), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n320), .A2(new_n687), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  OAI221_X1 g0754(.A(new_n948), .B1(new_n654), .B2(new_n875), .C1(new_n952), .C2(new_n954), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n453), .B(new_n757), .C1(new_n746), .C2(KEYINPUT29), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(new_n659), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n955), .B(new_n957), .Z(new_n958));
  OR2_X1    g0758(.A1(new_n942), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n942), .A2(new_n958), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n959), .B(new_n960), .C1(new_n206), .C2(new_n760), .ZN(new_n961));
  OAI211_X1 g0761(.A(G116), .B(new_n219), .C1(new_n577), .C2(KEYINPUT35), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n962), .B1(KEYINPUT35), .B2(new_n577), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT36), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n217), .B(G77), .C1(new_n788), .C2(new_n295), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(G50), .B2(new_n295), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n206), .A2(G13), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n964), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n961), .A2(new_n968), .ZN(G367));
  NAND2_X1  g0769(.A1(new_n669), .A2(new_n679), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n621), .A2(new_n687), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n748), .B2(new_n971), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n973), .A2(KEYINPUT107), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(KEYINPUT107), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n977), .A2(KEYINPUT43), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT110), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT109), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n604), .B(new_n610), .C1(new_n585), .C2(new_n688), .ZN(new_n983));
  OR3_X1    g0783(.A1(new_n708), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n982), .B1(new_n708), .B2(new_n983), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(KEYINPUT42), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT42), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n984), .A2(new_n985), .A3(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n610), .B1(new_n983), .B2(new_n561), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n688), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n987), .A2(new_n989), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n979), .B1(new_n981), .B2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n706), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n607), .A2(new_n609), .A3(new_n687), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n983), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n981), .A2(new_n992), .A3(new_n979), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n994), .A2(new_n995), .A3(new_n997), .A4(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n998), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n997), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n1000), .A2(new_n993), .B1(new_n706), .B2(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n717), .B(KEYINPUT41), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n710), .A2(new_n1001), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT45), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n710), .A2(new_n1001), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT44), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1006), .B(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1005), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n995), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n703), .B1(new_n691), .B2(new_n687), .ZN(new_n1011));
  AND3_X1   g0811(.A1(new_n1011), .A2(new_n694), .A3(new_n708), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n694), .B1(new_n1011), .B2(new_n708), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1005), .A2(new_n706), .A3(new_n1008), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n1010), .A2(new_n758), .A3(new_n1015), .A4(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1003), .B1(new_n1017), .B2(new_n758), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n761), .A2(G1), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n999), .B(new_n1002), .C1(new_n1018), .C2(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n776), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n240), .A2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n779), .B1(new_n210), .B2(new_n367), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n770), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(G137), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n787), .A2(new_n839), .B1(new_n803), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n792), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n1027), .A2(new_n295), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1029), .B(new_n252), .C1(new_n838), .C2(new_n785), .ZN(new_n1030));
  AOI211_X1 g0830(.A(new_n1026), .B(new_n1030), .C1(G50), .C2(new_n836), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(G58), .A2(new_n801), .B1(new_n808), .B2(G77), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1031), .B(new_n1032), .C1(new_n804), .C2(new_n846), .ZN(new_n1033));
  INV_X1    g0833(.A(G317), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n795), .A2(new_n847), .B1(new_n803), .B2(new_n1034), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n326), .B1(new_n785), .B2(new_n817), .C1(new_n1027), .C2(new_n376), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n1035), .B(new_n1036), .C1(G303), .C2(new_n819), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n846), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n1038), .A2(G294), .B1(G97), .B2(new_n808), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT46), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n801), .A2(G116), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1037), .B(new_n1039), .C1(new_n1040), .C2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1041), .A2(new_n1040), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT111), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1033), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT47), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  AND2_X1   g0847(.A1(new_n1047), .A2(new_n778), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1024), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n977), .B2(new_n768), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1020), .A2(new_n1051), .ZN(G387));
  INV_X1    g0852(.A(new_n719), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n771), .A2(new_n1053), .B1(G107), .B2(new_n210), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n236), .A2(G45), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n343), .A2(G50), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT50), .ZN(new_n1057));
  AOI211_X1 g0857(.A(G45), .B(new_n719), .C1(G68), .C2(G77), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1021), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1054), .B1(new_n1055), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n801), .A2(G77), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(new_n567), .B2(new_n807), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n785), .A2(new_n804), .B1(new_n787), .B2(new_n202), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n797), .A2(new_n343), .B1(new_n795), .B2(new_n295), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n252), .B1(new_n803), .B2(new_n839), .C1(new_n1027), .C2(new_n367), .ZN(new_n1065));
  NOR4_X1   g0865(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n326), .B1(new_n803), .B2(new_n821), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n835), .A2(G322), .B1(new_n836), .B2(G303), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n1034), .B2(new_n787), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(G311), .B2(new_n1038), .ZN(new_n1070));
  OR2_X1    g0870(.A1(new_n1070), .A2(KEYINPUT48), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1070), .A2(KEYINPUT48), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n801), .A2(G294), .B1(G283), .B2(new_n792), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT49), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n1067), .B(new_n1076), .C1(G116), .C2(new_n808), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1066), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n778), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n770), .B1(new_n780), .B2(new_n1060), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(new_n703), .B2(new_n767), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(new_n1015), .B2(new_n1019), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1015), .A2(new_n758), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(new_n718), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1015), .A2(new_n758), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1083), .B1(new_n1085), .B2(new_n1086), .ZN(G393));
  NAND2_X1  g0887(.A1(new_n1016), .A2(KEYINPUT112), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT112), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n1005), .A2(new_n706), .A3(new_n1008), .A4(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1088), .A2(new_n1010), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1019), .ZN(new_n1092));
  OR2_X1    g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n779), .B1(new_n567), .B2(new_n210), .C1(new_n1021), .C2(new_n247), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n770), .A2(new_n1094), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n252), .B1(new_n803), .B2(new_n838), .C1(new_n343), .C2(new_n795), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(G77), .B2(new_n792), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1097), .B(new_n843), .C1(new_n202), .C2(new_n846), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n785), .A2(new_n839), .B1(new_n787), .B2(new_n804), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT51), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1100), .B1(new_n295), .B2(new_n800), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n801), .A2(G283), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT52), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n785), .A2(new_n1034), .B1(new_n787), .B2(new_n817), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n1102), .B1(new_n1103), .B2(new_n1104), .C1(new_n846), .C2(new_n824), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n326), .B1(new_n795), .B2(new_n851), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(G322), .B2(new_n811), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n792), .A2(G116), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1104), .A2(new_n1103), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n809), .A2(new_n1107), .A3(new_n1108), .A4(new_n1109), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n1098), .A2(new_n1101), .B1(new_n1105), .B2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1095), .B1(new_n1111), .B2(new_n778), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n997), .B2(new_n768), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1091), .A2(new_n1084), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1017), .A2(new_n718), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1093), .B(new_n1113), .C1(new_n1115), .C2(new_n1116), .ZN(G390));
  INV_X1    g0917(.A(KEYINPUT116), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT114), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n744), .A2(G330), .A3(new_n921), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  XOR2_X1   g0921(.A(new_n953), .B(KEYINPUT113), .Z(new_n1122));
  INV_X1    g0922(.A(new_n944), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n863), .A2(new_n861), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1123), .B1(new_n756), .B2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1122), .B1(new_n1126), .B2(new_n946), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1127), .B1(new_n907), .B2(new_n935), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1123), .B1(new_n746), .B2(new_n865), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n954), .B1(new_n1129), .B2(new_n946), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n1121), .B(new_n1128), .C1(new_n952), .C2(new_n1130), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n918), .A2(G330), .A3(new_n865), .A4(new_n947), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n908), .A2(KEYINPUT39), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n935), .A2(new_n949), .A3(new_n907), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1130), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1128), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1132), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1119), .B1(new_n1131), .B2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n744), .A2(G330), .A3(new_n865), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(new_n946), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n1132), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n945), .ZN(new_n1142));
  AND2_X1   g0942(.A1(new_n1120), .A2(new_n1126), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n865), .A2(G330), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n946), .B1(new_n911), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1142), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n939), .A2(G330), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1148), .A2(new_n659), .A3(new_n956), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1147), .A2(new_n1150), .A3(KEYINPUT115), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT115), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n1141), .A2(new_n945), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1152), .B1(new_n1153), .B2(new_n1149), .ZN(new_n1154));
  AND2_X1   g0954(.A1(new_n1151), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1135), .A2(new_n1136), .A3(new_n1120), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1128), .B1(new_n952), .B2(new_n1130), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n1156), .B(KEYINPUT114), .C1(new_n1132), .C2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1138), .A2(new_n1155), .A3(new_n1158), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1131), .A2(new_n1137), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1153), .A2(new_n1149), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n717), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1118), .B1(new_n1159), .B2(new_n1162), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1156), .B(new_n1019), .C1(new_n1132), .C2(new_n1157), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n762), .B1(new_n343), .B2(new_n855), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n1038), .A2(G107), .B1(G68), .B2(new_n808), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n819), .A2(G116), .B1(new_n792), .B2(G77), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n1167), .B(KEYINPUT117), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n795), .A2(new_n567), .B1(new_n803), .B2(new_n851), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n252), .B(new_n1169), .C1(G283), .C2(new_n835), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1166), .A2(new_n1168), .A3(new_n802), .A4(new_n1170), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n1171), .A2(KEYINPUT118), .ZN(new_n1172));
  INV_X1    g0972(.A(G128), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(KEYINPUT54), .B(G143), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n785), .A2(new_n1173), .B1(new_n795), .B2(new_n1174), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n252), .B1(new_n787), .B2(new_n831), .C1(new_n1027), .C2(new_n804), .ZN(new_n1176));
  AOI211_X1 g0976(.A(new_n1175), .B(new_n1176), .C1(G125), .C2(new_n811), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n800), .A2(new_n839), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1178), .B(KEYINPUT53), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n1038), .A2(G137), .B1(G50), .B2(new_n808), .ZN(new_n1180));
  AND3_X1   g0980(.A1(new_n1177), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1171), .A2(KEYINPUT118), .ZN(new_n1182));
  NOR3_X1   g0982(.A1(new_n1172), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n1165), .B1(new_n1080), .B2(new_n1183), .C1(new_n1184), .C2(new_n766), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1164), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1186), .A2(KEYINPUT119), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT119), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1164), .A2(new_n1188), .A3(new_n1185), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1187), .A2(new_n1189), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1163), .A2(new_n1190), .ZN(new_n1191));
  AND3_X1   g0991(.A1(new_n1159), .A2(new_n1162), .A3(new_n1118), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1191), .A2(new_n1193), .ZN(G378));
  OAI211_X1 g0994(.A(new_n1156), .B(new_n1161), .C1(new_n1132), .C2(new_n1157), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(new_n1150), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n361), .B(new_n1197), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n347), .A2(new_n685), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(new_n1199), .B(KEYINPUT120), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n1198), .B(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(new_n938), .B2(G330), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n935), .A2(new_n907), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n925), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n937), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n906), .A2(new_n907), .B1(new_n917), .B2(new_n923), .ZN(new_n1207));
  OAI211_X1 g1007(.A(G330), .B(new_n1202), .C1(new_n1206), .C2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n955), .B1(new_n1203), .B2(new_n1209), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n1184), .A2(new_n953), .B1(new_n451), .B2(new_n685), .ZN(new_n1211));
  OAI21_X1  g1011(.A(G330), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(new_n1201), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1211), .A2(new_n1213), .A3(new_n948), .A4(new_n1208), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1210), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT57), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n1196), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1216), .B1(new_n1196), .B2(new_n1215), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n718), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n326), .A2(new_n476), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n1220), .B(new_n1028), .C1(new_n642), .C2(new_n836), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(G116), .A2(new_n835), .B1(new_n819), .B2(G107), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(G97), .A2(new_n798), .B1(new_n811), .B2(G283), .ZN(new_n1223));
  AND2_X1   g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n807), .A2(new_n788), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  AND4_X1   g1026(.A1(new_n1061), .A2(new_n1221), .A3(new_n1224), .A4(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(KEYINPUT58), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n1220), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1229));
  AND2_X1   g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n787), .A2(new_n1173), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n797), .A2(new_n831), .B1(new_n795), .B2(new_n1025), .ZN(new_n1232));
  AOI211_X1 g1032(.A(new_n1231), .B(new_n1232), .C1(G125), .C2(new_n835), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n1233), .B1(new_n839), .B2(new_n1027), .C1(new_n800), .C2(new_n1174), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1234), .A2(KEYINPUT59), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1234), .A2(KEYINPUT59), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n808), .A2(G159), .ZN(new_n1237));
  AOI211_X1 g1037(.A(G33), .B(G41), .C1(new_n811), .C2(G124), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1236), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n1230), .B1(KEYINPUT58), .B2(new_n1227), .C1(new_n1235), .C2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(new_n778), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n762), .B1(new_n202), .B2(new_n855), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1241), .B(new_n1242), .C1(new_n1202), .C2(new_n766), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(new_n1215), .B2(new_n1019), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1219), .A2(new_n1245), .ZN(G375));
  INV_X1    g1046(.A(new_n1003), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1153), .A2(new_n1149), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1155), .A2(new_n1247), .A3(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n762), .B1(new_n295), .B2(new_n855), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(new_n1250), .B(KEYINPUT121), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n785), .A2(new_n831), .ZN(new_n1252));
  XNOR2_X1  g1052(.A(new_n1252), .B(KEYINPUT122), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1226), .B1(new_n846), .B2(new_n1174), .ZN(new_n1254));
  AOI211_X1 g1054(.A(new_n1253), .B(new_n1254), .C1(G159), .C2(new_n801), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n252), .B1(new_n787), .B2(new_n1025), .ZN(new_n1256));
  OAI22_X1  g1056(.A1(new_n795), .A2(new_n839), .B1(new_n803), .B2(new_n1173), .ZN(new_n1257));
  AOI211_X1 g1057(.A(new_n1256), .B(new_n1257), .C1(G50), .C2(new_n792), .ZN(new_n1258));
  OAI22_X1  g1058(.A1(new_n785), .A2(new_n851), .B1(new_n795), .B2(new_n376), .ZN(new_n1259));
  OAI221_X1 g1059(.A(new_n326), .B1(new_n787), .B2(new_n847), .C1(new_n1027), .C2(new_n367), .ZN(new_n1260));
  AOI211_X1 g1060(.A(new_n1259), .B(new_n1260), .C1(G303), .C2(new_n811), .ZN(new_n1261));
  OAI22_X1  g1061(.A1(new_n297), .A2(new_n807), .B1(new_n800), .B2(new_n567), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1262), .B1(new_n1038), .B2(G116), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n1255), .A2(new_n1258), .B1(new_n1261), .B2(new_n1263), .ZN(new_n1264));
  OAI221_X1 g1064(.A(new_n1251), .B1(new_n1080), .B2(new_n1264), .C1(new_n947), .C2(new_n766), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1265), .B1(new_n1153), .B2(new_n1092), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1249), .A2(new_n1267), .ZN(G381));
  OAI21_X1  g1068(.A(new_n1113), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1116), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1269), .B1(new_n1270), .B2(new_n1114), .ZN(new_n1271));
  INV_X1    g1071(.A(G384), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  OR2_X1    g1073(.A1(G393), .A2(G396), .ZN(new_n1274));
  NOR4_X1   g1074(.A1(new_n1273), .A2(G387), .A3(G381), .A4(new_n1274), .ZN(new_n1275));
  XNOR2_X1  g1075(.A(new_n1275), .B(KEYINPUT123), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1245), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1196), .A2(new_n1215), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(KEYINPUT57), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1196), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1277), .B1(new_n1281), .B2(new_n718), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1186), .B1(new_n1159), .B2(new_n1162), .ZN(new_n1283));
  AND2_X1   g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1276), .A2(new_n1284), .ZN(G407));
  INV_X1    g1085(.A(G213), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1286), .A2(G343), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1284), .A2(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(G407), .A2(G213), .A3(new_n1288), .ZN(G409));
  OAI21_X1  g1089(.A(new_n1245), .B1(new_n1278), .B2(new_n1003), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(new_n1283), .ZN(new_n1291));
  NOR3_X1   g1091(.A1(new_n1192), .A2(new_n1163), .A3(new_n1190), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1291), .B1(G375), .B2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1287), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT60), .ZN(new_n1295));
  XNOR2_X1  g1095(.A(new_n1248), .B(new_n1295), .ZN(new_n1296));
  NOR3_X1   g1096(.A1(new_n1296), .A2(new_n717), .A3(new_n1161), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1272), .B1(new_n1297), .B2(new_n1266), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n718), .B1(new_n1153), .B2(new_n1149), .ZN(new_n1299));
  OAI211_X1 g1099(.A(G384), .B(new_n1267), .C1(new_n1296), .C2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1298), .A2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1293), .A2(new_n1294), .A3(new_n1302), .ZN(new_n1303));
  XNOR2_X1  g1103(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT61), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT62), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1293), .A2(new_n1307), .A3(new_n1294), .A4(new_n1302), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1301), .A2(G2897), .A3(new_n1287), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1287), .A2(G2897), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1298), .A2(new_n1300), .A3(new_n1310), .ZN(new_n1311));
  AND2_X1   g1111(.A1(new_n1309), .A2(new_n1311), .ZN(new_n1312));
  AOI22_X1  g1112(.A1(new_n1282), .A2(G378), .B1(new_n1283), .B2(new_n1290), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1312), .B1(new_n1313), .B2(new_n1287), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1305), .A2(new_n1306), .A3(new_n1308), .A4(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(G393), .A2(G396), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(G387), .A2(new_n1271), .ZN(new_n1317));
  AOI21_X1  g1117(.A(G390), .B1(new_n1020), .B2(new_n1051), .ZN(new_n1318));
  OAI211_X1 g1118(.A(new_n1274), .B(new_n1316), .C1(new_n1317), .C2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1274), .A2(new_n1316), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT124), .ZN(new_n1321));
  NAND4_X1  g1121(.A1(G390), .A2(new_n1321), .A3(new_n1020), .A4(new_n1051), .ZN(new_n1322));
  AOI21_X1  g1122(.A(KEYINPUT124), .B1(G387), .B2(new_n1271), .ZN(new_n1323));
  OAI211_X1 g1123(.A(new_n1320), .B(new_n1322), .C1(new_n1323), .C2(new_n1317), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1319), .B1(new_n1324), .B2(KEYINPUT125), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT125), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(G390), .A2(new_n1020), .A3(new_n1051), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1327), .B1(new_n1318), .B2(KEYINPUT124), .ZN(new_n1328));
  AND2_X1   g1128(.A1(new_n1322), .A2(new_n1320), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1326), .B1(new_n1328), .B2(new_n1329), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1325), .A2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1315), .A2(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1309), .A2(new_n1311), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1333), .B1(new_n1294), .B2(new_n1293), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT63), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n1303), .B1(new_n1334), .B2(new_n1335), .ZN(new_n1336));
  NOR2_X1   g1136(.A1(new_n1331), .A2(KEYINPUT61), .ZN(new_n1337));
  OR2_X1    g1137(.A1(new_n1303), .A2(new_n1335), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1336), .A2(new_n1337), .A3(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1332), .A2(new_n1339), .ZN(G405));
  NAND2_X1  g1140(.A1(new_n1282), .A2(G378), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(G375), .A2(new_n1283), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1341), .A2(new_n1342), .ZN(new_n1343));
  OR2_X1    g1143(.A1(new_n1343), .A2(KEYINPUT127), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1343), .A2(KEYINPUT127), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1344), .A2(new_n1345), .ZN(new_n1346));
  OAI21_X1  g1146(.A(new_n1301), .B1(new_n1325), .B2(new_n1330), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1324), .A2(KEYINPUT125), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1328), .A2(new_n1329), .A3(new_n1326), .ZN(new_n1349));
  NAND4_X1  g1149(.A1(new_n1348), .A2(new_n1349), .A3(new_n1319), .A4(new_n1302), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1346), .A2(new_n1347), .A3(new_n1350), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1347), .A2(new_n1350), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1352), .A2(new_n1345), .A3(new_n1344), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1351), .A2(new_n1353), .ZN(G402));
endmodule


