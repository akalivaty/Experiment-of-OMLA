
module locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, 
        G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, 
        G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, 
        G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39, 
        G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584;

  INV_X1 U297 ( .A(G953), .ZN(n574) );
  NOR2_X2 U298 ( .A1(n584), .A2(n583), .ZN(n458) );
  AND2_X2 U299 ( .A1(n325), .A2(n324), .ZN(n427) );
  XNOR2_X2 U300 ( .A(n399), .B(n336), .ZN(n570) );
  XNOR2_X2 U301 ( .A(n384), .B(G128), .ZN(n399) );
  AND2_X2 U302 ( .A1(n299), .A2(n304), .ZN(n551) );
  NAND2_X1 U303 ( .A1(n296), .A2(n295), .ZN(n299) );
  AND2_X1 U304 ( .A1(n331), .A2(KEYINPUT44), .ZN(n327) );
  XNOR2_X1 U305 ( .A(n415), .B(KEYINPUT32), .ZN(n582) );
  NOR2_X1 U306 ( .A1(n446), .A2(n417), .ZN(n418) );
  AND2_X1 U307 ( .A1(n409), .A2(n408), .ZN(n411) );
  XNOR2_X1 U308 ( .A(n444), .B(KEYINPUT1), .ZN(n501) );
  XNOR2_X1 U309 ( .A(n543), .B(n542), .ZN(n544) );
  NAND2_X1 U310 ( .A1(n300), .A2(KEYINPUT2), .ZN(n295) );
  XNOR2_X1 U311 ( .A(n333), .B(n332), .ZN(n450) );
  NOR2_X2 U312 ( .A1(n555), .A2(n546), .ZN(n547) );
  XNOR2_X2 U313 ( .A(KEYINPUT0), .B(n352), .ZN(n409) );
  XNOR2_X1 U314 ( .A(n570), .B(n337), .ZN(n377) );
  INV_X1 U315 ( .A(G101), .ZN(n337) );
  NOR2_X1 U316 ( .A1(n581), .A2(KEYINPUT44), .ZN(n329) );
  NOR2_X1 U317 ( .A1(n432), .A2(n407), .ZN(n502) );
  INV_X1 U318 ( .A(KEYINPUT47), .ZN(n287) );
  INV_X1 U319 ( .A(KEYINPUT4), .ZN(n336) );
  XNOR2_X1 U320 ( .A(n292), .B(n291), .ZN(n395) );
  INV_X1 U321 ( .A(KEYINPUT8), .ZN(n291) );
  XOR2_X1 U322 ( .A(G125), .B(KEYINPUT10), .Z(n569) );
  XNOR2_X1 U323 ( .A(n311), .B(G131), .ZN(n387) );
  INV_X1 U324 ( .A(G146), .ZN(n311) );
  XOR2_X1 U325 ( .A(G137), .B(G140), .Z(n357) );
  XNOR2_X1 U326 ( .A(n387), .B(G134), .ZN(n371) );
  XNOR2_X1 U327 ( .A(n315), .B(KEYINPUT48), .ZN(n464) );
  AND2_X1 U328 ( .A1(n318), .A2(n281), .ZN(n317) );
  AND2_X1 U329 ( .A1(n432), .A2(n293), .ZN(n445) );
  AND2_X1 U330 ( .A1(n496), .A2(n276), .ZN(n293) );
  XNOR2_X1 U331 ( .A(n356), .B(n355), .ZN(n444) );
  INV_X1 U332 ( .A(G469), .ZN(n355) );
  NOR2_X1 U333 ( .A1(G902), .A2(n539), .ZN(n356) );
  XNOR2_X1 U334 ( .A(n340), .B(n313), .ZN(n372) );
  XNOR2_X1 U335 ( .A(n314), .B(G116), .ZN(n313) );
  INV_X1 U336 ( .A(G113), .ZN(n314) );
  XNOR2_X1 U337 ( .A(G110), .B(G128), .ZN(n358) );
  XNOR2_X1 U338 ( .A(n377), .B(n339), .ZN(n353) );
  INV_X1 U339 ( .A(n562), .ZN(n339) );
  XNOR2_X1 U340 ( .A(n422), .B(n421), .ZN(n524) );
  NAND2_X1 U341 ( .A1(n330), .A2(n329), .ZN(n324) );
  XNOR2_X1 U342 ( .A(n319), .B(KEYINPUT39), .ZN(n465) );
  NOR2_X1 U343 ( .A1(n524), .A2(n423), .ZN(n309) );
  XNOR2_X1 U344 ( .A(n378), .B(G472), .ZN(n500) );
  XNOR2_X1 U345 ( .A(n411), .B(n410), .ZN(n416) );
  INV_X1 U346 ( .A(KEYINPUT22), .ZN(n410) );
  XNOR2_X1 U347 ( .A(n372), .B(n335), .ZN(n563) );
  XNOR2_X1 U348 ( .A(KEYINPUT16), .B(G122), .ZN(n335) );
  NOR2_X1 U349 ( .A1(n282), .A2(n285), .ZN(n281) );
  NOR2_X1 U350 ( .A1(n485), .A2(n286), .ZN(n285) );
  NAND2_X1 U351 ( .A1(n288), .A2(n287), .ZN(n286) );
  NAND2_X1 U352 ( .A1(G237), .A2(G234), .ZN(n348) );
  XOR2_X1 U353 ( .A(n451), .B(KEYINPUT38), .Z(n511) );
  NAND2_X1 U354 ( .A1(n501), .A2(n502), .ZN(n419) );
  OR2_X1 U355 ( .A1(G902), .A2(G237), .ZN(n347) );
  XNOR2_X1 U356 ( .A(n312), .B(n371), .ZN(n376) );
  XNOR2_X1 U357 ( .A(n375), .B(n372), .ZN(n312) );
  XNOR2_X1 U358 ( .A(G104), .B(G110), .ZN(n338) );
  INV_X1 U359 ( .A(n573), .ZN(n298) );
  NOR2_X1 U360 ( .A1(G953), .A2(G237), .ZN(n388) );
  OR2_X1 U361 ( .A1(n559), .A2(n303), .ZN(n304) );
  AND2_X1 U362 ( .A1(n320), .A2(n440), .ZN(n452) );
  AND2_X1 U363 ( .A1(n441), .A2(n276), .ZN(n320) );
  INV_X1 U364 ( .A(KEYINPUT19), .ZN(n332) );
  XNOR2_X1 U365 ( .A(n368), .B(n294), .ZN(n432) );
  INV_X1 U366 ( .A(KEYINPUT25), .ZN(n294) );
  XNOR2_X1 U367 ( .A(n290), .B(n362), .ZN(n363) );
  XNOR2_X1 U368 ( .A(n353), .B(n310), .ZN(n539) );
  XNOR2_X1 U369 ( .A(n571), .B(n354), .ZN(n310) );
  XNOR2_X1 U370 ( .A(n353), .B(n334), .ZN(n532) );
  XNOR2_X1 U371 ( .A(n563), .B(n345), .ZN(n334) );
  XOR2_X1 U372 ( .A(G146), .B(G125), .Z(n343) );
  NAND2_X1 U373 ( .A1(n308), .A2(n307), .ZN(n306) );
  INV_X1 U374 ( .A(n443), .ZN(n307) );
  XNOR2_X1 U375 ( .A(n309), .B(KEYINPUT34), .ZN(n308) );
  OR2_X1 U376 ( .A1(n416), .A2(n321), .ZN(n415) );
  NAND2_X1 U377 ( .A1(n414), .A2(n322), .ZN(n321) );
  INV_X1 U378 ( .A(n433), .ZN(n322) );
  OR2_X1 U379 ( .A1(n450), .A2(n456), .ZN(n485) );
  INV_X1 U380 ( .A(G143), .ZN(n384) );
  AND2_X1 U381 ( .A1(G210), .A2(n347), .ZN(n275) );
  OR2_X1 U382 ( .A1(n431), .A2(n430), .ZN(n276) );
  AND2_X1 U383 ( .A1(n494), .A2(KEYINPUT2), .ZN(n277) );
  AND2_X1 U384 ( .A1(n301), .A2(n302), .ZN(n278) );
  AND2_X1 U385 ( .A1(n289), .A2(n284), .ZN(n279) );
  XNOR2_X1 U386 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n280) );
  INV_X1 U387 ( .A(KEYINPUT2), .ZN(n305) );
  NAND2_X1 U388 ( .A1(n283), .A2(n279), .ZN(n282) );
  NAND2_X1 U389 ( .A1(n485), .A2(KEYINPUT47), .ZN(n283) );
  NAND2_X1 U390 ( .A1(n515), .A2(KEYINPUT47), .ZN(n284) );
  INV_X1 U391 ( .A(n515), .ZN(n288) );
  INV_X1 U392 ( .A(n484), .ZN(n289) );
  NAND2_X1 U393 ( .A1(n395), .A2(G221), .ZN(n290) );
  NAND2_X1 U394 ( .A1(n574), .A2(G234), .ZN(n292) );
  NAND2_X1 U395 ( .A1(n559), .A2(n305), .ZN(n301) );
  NAND2_X1 U396 ( .A1(n573), .A2(n305), .ZN(n302) );
  NAND2_X1 U397 ( .A1(n298), .A2(n297), .ZN(n296) );
  NOR2_X2 U398 ( .A1(n559), .A2(n468), .ZN(n297) );
  NAND2_X1 U399 ( .A1(n278), .A2(n304), .ZN(n528) );
  INV_X1 U400 ( .A(n468), .ZN(n300) );
  NAND2_X1 U401 ( .A1(n467), .A2(n494), .ZN(n573) );
  XNOR2_X2 U402 ( .A(n427), .B(KEYINPUT45), .ZN(n559) );
  NAND2_X1 U403 ( .A1(n467), .A2(n277), .ZN(n303) );
  XNOR2_X2 U404 ( .A(n306), .B(KEYINPUT35), .ZN(n581) );
  NOR2_X2 U405 ( .A1(n495), .A2(n464), .ZN(n467) );
  NOR2_X2 U406 ( .A1(n555), .A2(n535), .ZN(n536) );
  NAND2_X1 U407 ( .A1(n317), .A2(n316), .ZN(n315) );
  XNOR2_X1 U408 ( .A(n458), .B(KEYINPUT46), .ZN(n316) );
  INV_X1 U409 ( .A(n492), .ZN(n318) );
  NAND2_X1 U410 ( .A1(n452), .A2(n511), .ZN(n319) );
  OR2_X1 U411 ( .A1(n416), .A2(n433), .ZN(n323) );
  NOR2_X1 U412 ( .A1(n323), .A2(n501), .ZN(n412) );
  NOR2_X1 U413 ( .A1(n327), .A2(n326), .ZN(n325) );
  NAND2_X1 U414 ( .A1(n328), .A2(n426), .ZN(n326) );
  NAND2_X1 U415 ( .A1(n581), .A2(KEYINPUT44), .ZN(n328) );
  INV_X1 U416 ( .A(n331), .ZN(n330) );
  NAND2_X1 U417 ( .A1(n582), .A2(n481), .ZN(n331) );
  NOR2_X1 U418 ( .A1(n460), .A2(n333), .ZN(n461) );
  NAND2_X1 U419 ( .A1(n451), .A2(n510), .ZN(n333) );
  NOR2_X1 U420 ( .A1(n472), .A2(n555), .ZN(n474) );
  XNOR2_X1 U421 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U422 ( .A(n532), .B(n280), .ZN(n533) );
  NOR2_X2 U423 ( .A1(n450), .A2(n351), .ZN(n352) );
  INV_X1 U424 ( .A(KEYINPUT33), .ZN(n421) );
  XNOR2_X1 U425 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U426 ( .A(n469), .B(KEYINPUT62), .ZN(n470) );
  INV_X1 U427 ( .A(n501), .ZN(n463) );
  XNOR2_X1 U428 ( .A(n545), .B(n544), .ZN(n546) );
  INV_X1 U429 ( .A(KEYINPUT63), .ZN(n473) );
  NOR2_X1 U430 ( .A1(G952), .A2(n574), .ZN(n555) );
  XNOR2_X1 U431 ( .A(G902), .B(KEYINPUT15), .ZN(n468) );
  XNOR2_X1 U432 ( .A(n338), .B(G107), .ZN(n562) );
  XNOR2_X1 U433 ( .A(KEYINPUT3), .B(G119), .ZN(n340) );
  XOR2_X1 U434 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n342) );
  NAND2_X1 U435 ( .A1(G224), .A2(n574), .ZN(n341) );
  XNOR2_X1 U436 ( .A(n342), .B(n341), .ZN(n344) );
  NAND2_X1 U437 ( .A1(n468), .A2(n532), .ZN(n346) );
  XNOR2_X2 U438 ( .A(n346), .B(n275), .ZN(n451) );
  NAND2_X1 U439 ( .A1(G214), .A2(n347), .ZN(n510) );
  XNOR2_X1 U440 ( .A(n348), .B(KEYINPUT14), .ZN(n349) );
  NAND2_X1 U441 ( .A1(G952), .A2(n349), .ZN(n523) );
  NOR2_X1 U442 ( .A1(G953), .A2(n523), .ZN(n431) );
  INV_X1 U443 ( .A(G898), .ZN(n558) );
  NAND2_X1 U444 ( .A1(G953), .A2(n558), .ZN(n565) );
  NAND2_X1 U445 ( .A1(G902), .A2(n349), .ZN(n428) );
  NOR2_X1 U446 ( .A1(n565), .A2(n428), .ZN(n350) );
  NOR2_X1 U447 ( .A1(n431), .A2(n350), .ZN(n351) );
  INV_X1 U448 ( .A(n409), .ZN(n423) );
  XNOR2_X1 U449 ( .A(n357), .B(n371), .ZN(n571) );
  AND2_X1 U450 ( .A1(G227), .A2(n574), .ZN(n354) );
  XNOR2_X1 U451 ( .A(n357), .B(n569), .ZN(n361) );
  XOR2_X1 U452 ( .A(G146), .B(G119), .Z(n359) );
  XNOR2_X1 U453 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U454 ( .A(n361), .B(n360), .ZN(n364) );
  XOR2_X1 U455 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n362) );
  XNOR2_X1 U456 ( .A(n364), .B(n363), .ZN(n553) );
  NOR2_X1 U457 ( .A1(n553), .A2(G902), .ZN(n367) );
  NAND2_X1 U458 ( .A1(G234), .A2(n468), .ZN(n365) );
  XNOR2_X1 U459 ( .A(KEYINPUT20), .B(n365), .ZN(n369) );
  NAND2_X1 U460 ( .A1(n369), .A2(G217), .ZN(n366) );
  XNOR2_X1 U461 ( .A(n367), .B(n366), .ZN(n368) );
  NAND2_X1 U462 ( .A1(n369), .A2(G221), .ZN(n370) );
  XOR2_X1 U463 ( .A(KEYINPUT21), .B(n370), .Z(n496) );
  INV_X1 U464 ( .A(n496), .ZN(n407) );
  NAND2_X1 U465 ( .A1(n444), .A2(n502), .ZN(n438) );
  NOR2_X1 U466 ( .A1(n423), .A2(n438), .ZN(n379) );
  XOR2_X1 U467 ( .A(G137), .B(KEYINPUT5), .Z(n374) );
  NAND2_X1 U468 ( .A1(n388), .A2(G210), .ZN(n373) );
  XNOR2_X1 U469 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U470 ( .A(n377), .B(n376), .ZN(n469) );
  NOR2_X1 U471 ( .A1(n469), .A2(G902), .ZN(n378) );
  NAND2_X1 U472 ( .A1(n379), .A2(n500), .ZN(n477) );
  NOR2_X1 U473 ( .A1(n500), .A2(n419), .ZN(n507) );
  NAND2_X1 U474 ( .A1(n409), .A2(n507), .ZN(n380) );
  XOR2_X1 U475 ( .A(KEYINPUT31), .B(n380), .Z(n489) );
  NAND2_X1 U476 ( .A1(n477), .A2(n489), .ZN(n406) );
  XOR2_X1 U477 ( .A(KEYINPUT11), .B(G140), .Z(n382) );
  XNOR2_X1 U478 ( .A(G113), .B(G122), .ZN(n381) );
  XNOR2_X1 U479 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U480 ( .A(n383), .B(n569), .Z(n386) );
  XNOR2_X1 U481 ( .A(G104), .B(G143), .ZN(n385) );
  XNOR2_X1 U482 ( .A(n386), .B(n385), .ZN(n392) );
  XOR2_X1 U483 ( .A(n387), .B(KEYINPUT12), .Z(n390) );
  NAND2_X1 U484 ( .A1(G214), .A2(n388), .ZN(n389) );
  XNOR2_X1 U485 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U486 ( .A(n392), .B(n391), .ZN(n543) );
  NOR2_X1 U487 ( .A1(G902), .A2(n543), .ZN(n394) );
  XNOR2_X1 U488 ( .A(KEYINPUT13), .B(G475), .ZN(n393) );
  XNOR2_X1 U489 ( .A(n394), .B(n393), .ZN(n424) );
  INV_X1 U490 ( .A(n424), .ZN(n405) );
  XOR2_X1 U491 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n397) );
  NAND2_X1 U492 ( .A1(G217), .A2(n395), .ZN(n396) );
  XNOR2_X1 U493 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U494 ( .A(n398), .B(G116), .Z(n401) );
  XNOR2_X1 U495 ( .A(G107), .B(n399), .ZN(n400) );
  XNOR2_X1 U496 ( .A(n401), .B(n400), .ZN(n403) );
  XOR2_X1 U497 ( .A(G122), .B(G134), .Z(n402) );
  XNOR2_X1 U498 ( .A(n403), .B(n402), .ZN(n549) );
  NOR2_X1 U499 ( .A1(n549), .A2(G902), .ZN(n404) );
  XOR2_X1 U500 ( .A(n404), .B(G478), .Z(n425) );
  NOR2_X1 U501 ( .A1(n405), .A2(n425), .ZN(n453) );
  NAND2_X1 U502 ( .A1(n405), .A2(n425), .ZN(n490) );
  INV_X1 U503 ( .A(n490), .ZN(n466) );
  NOR2_X1 U504 ( .A1(n453), .A2(n466), .ZN(n515) );
  NAND2_X1 U505 ( .A1(n406), .A2(n288), .ZN(n413) );
  XNOR2_X1 U506 ( .A(KEYINPUT6), .B(n500), .ZN(n433) );
  OR2_X1 U507 ( .A1(n425), .A2(n424), .ZN(n513) );
  NOR2_X1 U508 ( .A1(n513), .A2(n407), .ZN(n408) );
  INV_X1 U509 ( .A(n432), .ZN(n497) );
  NAND2_X1 U510 ( .A1(n412), .A2(n497), .ZN(n475) );
  AND2_X1 U511 ( .A1(n413), .A2(n475), .ZN(n426) );
  NOR2_X1 U512 ( .A1(n497), .A2(n463), .ZN(n414) );
  INV_X1 U513 ( .A(n500), .ZN(n446) );
  OR2_X1 U514 ( .A1(n501), .A2(n416), .ZN(n417) );
  NAND2_X1 U515 ( .A1(n432), .A2(n418), .ZN(n481) );
  INV_X1 U516 ( .A(n419), .ZN(n420) );
  NAND2_X1 U517 ( .A1(n420), .A2(n433), .ZN(n422) );
  NAND2_X1 U518 ( .A1(n425), .A2(n424), .ZN(n443) );
  INV_X1 U519 ( .A(n453), .ZN(n487) );
  OR2_X1 U520 ( .A1(n574), .A2(n428), .ZN(n429) );
  NOR2_X1 U521 ( .A1(G900), .A2(n429), .ZN(n430) );
  NAND2_X1 U522 ( .A1(n433), .A2(n445), .ZN(n434) );
  NOR2_X1 U523 ( .A1(n487), .A2(n434), .ZN(n459) );
  NAND2_X1 U524 ( .A1(n459), .A2(n510), .ZN(n435) );
  NOR2_X1 U525 ( .A1(n501), .A2(n435), .ZN(n436) );
  XNOR2_X1 U526 ( .A(n436), .B(KEYINPUT43), .ZN(n437) );
  NOR2_X1 U527 ( .A1(n451), .A2(n437), .ZN(n495) );
  INV_X1 U528 ( .A(n438), .ZN(n441) );
  NAND2_X1 U529 ( .A1(n446), .A2(n510), .ZN(n439) );
  XOR2_X1 U530 ( .A(KEYINPUT30), .B(n439), .Z(n440) );
  NAND2_X1 U531 ( .A1(n451), .A2(n452), .ZN(n442) );
  NOR2_X1 U532 ( .A1(n443), .A2(n442), .ZN(n484) );
  INV_X1 U533 ( .A(n444), .ZN(n449) );
  AND2_X1 U534 ( .A1(n446), .A2(n445), .ZN(n447) );
  XOR2_X1 U535 ( .A(KEYINPUT28), .B(n447), .Z(n448) );
  OR2_X1 U536 ( .A1(n449), .A2(n448), .ZN(n456) );
  AND2_X1 U537 ( .A1(n465), .A2(n453), .ZN(n454) );
  XNOR2_X1 U538 ( .A(n454), .B(KEYINPUT40), .ZN(n584) );
  NAND2_X1 U539 ( .A1(n511), .A2(n510), .ZN(n514) );
  NOR2_X1 U540 ( .A1(n513), .A2(n514), .ZN(n455) );
  XNOR2_X1 U541 ( .A(KEYINPUT41), .B(n455), .ZN(n525) );
  NOR2_X1 U542 ( .A1(n525), .A2(n456), .ZN(n457) );
  XNOR2_X1 U543 ( .A(KEYINPUT42), .B(n457), .ZN(n583) );
  INV_X1 U544 ( .A(n459), .ZN(n460) );
  XOR2_X1 U545 ( .A(KEYINPUT36), .B(n461), .Z(n462) );
  NOR2_X1 U546 ( .A1(n463), .A2(n462), .ZN(n492) );
  NAND2_X1 U547 ( .A1(n466), .A2(n465), .ZN(n494) );
  NAND2_X1 U548 ( .A1(n551), .A2(G472), .ZN(n471) );
  XNOR2_X1 U549 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U550 ( .A(n474), .B(n473), .ZN(G57) );
  XNOR2_X1 U551 ( .A(G101), .B(n475), .ZN(G3) );
  NOR2_X1 U552 ( .A1(n487), .A2(n477), .ZN(n476) );
  XOR2_X1 U553 ( .A(G104), .B(n476), .Z(G6) );
  NOR2_X1 U554 ( .A1(n490), .A2(n477), .ZN(n479) );
  XNOR2_X1 U555 ( .A(KEYINPUT26), .B(KEYINPUT27), .ZN(n478) );
  XNOR2_X1 U556 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U557 ( .A(G107), .B(n480), .ZN(G9) );
  XNOR2_X1 U558 ( .A(G110), .B(n481), .ZN(G12) );
  NOR2_X1 U559 ( .A1(n490), .A2(n485), .ZN(n483) );
  XNOR2_X1 U560 ( .A(G128), .B(KEYINPUT29), .ZN(n482) );
  XNOR2_X1 U561 ( .A(n483), .B(n482), .ZN(G30) );
  XOR2_X1 U562 ( .A(G143), .B(n484), .Z(G45) );
  NOR2_X1 U563 ( .A1(n487), .A2(n485), .ZN(n486) );
  XOR2_X1 U564 ( .A(G146), .B(n486), .Z(G48) );
  NOR2_X1 U565 ( .A1(n487), .A2(n489), .ZN(n488) );
  XOR2_X1 U566 ( .A(G113), .B(n488), .Z(G15) );
  NOR2_X1 U567 ( .A1(n490), .A2(n489), .ZN(n491) );
  XOR2_X1 U568 ( .A(G116), .B(n491), .Z(G18) );
  XNOR2_X1 U569 ( .A(G125), .B(n492), .ZN(n493) );
  XNOR2_X1 U570 ( .A(n493), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U571 ( .A(G134), .B(n494), .ZN(G36) );
  XOR2_X1 U572 ( .A(G140), .B(n495), .Z(G42) );
  NOR2_X1 U573 ( .A1(n497), .A2(n496), .ZN(n498) );
  XNOR2_X1 U574 ( .A(n498), .B(KEYINPUT49), .ZN(n499) );
  NAND2_X1 U575 ( .A1(n500), .A2(n499), .ZN(n505) );
  NOR2_X1 U576 ( .A1(n502), .A2(n501), .ZN(n503) );
  XNOR2_X1 U577 ( .A(n503), .B(KEYINPUT50), .ZN(n504) );
  NOR2_X1 U578 ( .A1(n505), .A2(n504), .ZN(n506) );
  NOR2_X1 U579 ( .A1(n507), .A2(n506), .ZN(n508) );
  XOR2_X1 U580 ( .A(KEYINPUT51), .B(n508), .Z(n509) );
  NOR2_X1 U581 ( .A1(n525), .A2(n509), .ZN(n520) );
  NOR2_X1 U582 ( .A1(n511), .A2(n510), .ZN(n512) );
  NOR2_X1 U583 ( .A1(n513), .A2(n512), .ZN(n517) );
  NOR2_X1 U584 ( .A1(n515), .A2(n514), .ZN(n516) );
  NOR2_X1 U585 ( .A1(n517), .A2(n516), .ZN(n518) );
  NOR2_X1 U586 ( .A1(n518), .A2(n524), .ZN(n519) );
  NOR2_X1 U587 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U588 ( .A(n521), .B(KEYINPUT52), .ZN(n522) );
  NOR2_X1 U589 ( .A1(n523), .A2(n522), .ZN(n527) );
  NOR2_X1 U590 ( .A1(n525), .A2(n524), .ZN(n526) );
  NOR2_X1 U591 ( .A1(n527), .A2(n526), .ZN(n529) );
  NAND2_X1 U592 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U593 ( .A1(n530), .A2(G953), .ZN(n531) );
  XNOR2_X1 U594 ( .A(n531), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U595 ( .A1(n551), .A2(G210), .ZN(n534) );
  XNOR2_X1 U596 ( .A(KEYINPUT56), .B(n536), .ZN(G51) );
  XOR2_X1 U597 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n538) );
  NAND2_X1 U598 ( .A1(n551), .A2(G469), .ZN(n537) );
  XNOR2_X1 U599 ( .A(n538), .B(n537), .ZN(n540) );
  XNOR2_X1 U600 ( .A(n540), .B(n539), .ZN(n541) );
  NOR2_X1 U601 ( .A1(n555), .A2(n541), .ZN(G54) );
  NAND2_X1 U602 ( .A1(n551), .A2(G475), .ZN(n545) );
  INV_X1 U603 ( .A(KEYINPUT59), .ZN(n542) );
  XNOR2_X1 U604 ( .A(KEYINPUT60), .B(n547), .ZN(G60) );
  NAND2_X1 U605 ( .A1(G478), .A2(n551), .ZN(n548) );
  XNOR2_X1 U606 ( .A(n549), .B(n548), .ZN(n550) );
  NOR2_X1 U607 ( .A1(n555), .A2(n550), .ZN(G63) );
  NAND2_X1 U608 ( .A1(G217), .A2(n551), .ZN(n552) );
  XNOR2_X1 U609 ( .A(n553), .B(n552), .ZN(n554) );
  NOR2_X1 U610 ( .A1(n555), .A2(n554), .ZN(G66) );
  NAND2_X1 U611 ( .A1(G953), .A2(G224), .ZN(n556) );
  XOR2_X1 U612 ( .A(KEYINPUT61), .B(n556), .Z(n557) );
  NOR2_X1 U613 ( .A1(n558), .A2(n557), .ZN(n561) );
  NOR2_X1 U614 ( .A1(G953), .A2(n559), .ZN(n560) );
  NOR2_X1 U615 ( .A1(n561), .A2(n560), .ZN(n568) );
  XNOR2_X1 U616 ( .A(n562), .B(G101), .ZN(n564) );
  XNOR2_X1 U617 ( .A(n564), .B(n563), .ZN(n566) );
  NAND2_X1 U618 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U619 ( .A(n568), .B(n567), .ZN(G69) );
  XNOR2_X1 U620 ( .A(n570), .B(n569), .ZN(n572) );
  XNOR2_X1 U621 ( .A(n572), .B(n571), .ZN(n576) );
  XNOR2_X1 U622 ( .A(n573), .B(n576), .ZN(n575) );
  NAND2_X1 U623 ( .A1(n575), .A2(n574), .ZN(n580) );
  XNOR2_X1 U624 ( .A(G227), .B(n576), .ZN(n577) );
  NAND2_X1 U625 ( .A1(n577), .A2(G900), .ZN(n578) );
  NAND2_X1 U626 ( .A1(n578), .A2(G953), .ZN(n579) );
  NAND2_X1 U627 ( .A1(n580), .A2(n579), .ZN(G72) );
  XOR2_X1 U628 ( .A(n581), .B(G122), .Z(G24) );
  XNOR2_X1 U629 ( .A(n582), .B(G119), .ZN(G21) );
  XOR2_X1 U630 ( .A(G137), .B(n583), .Z(G39) );
  XOR2_X1 U631 ( .A(n584), .B(G131), .Z(G33) );
endmodule

