//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 1 1 0 0 0 1 1 1 0 0 1 0 0 0 0 1 1 0 1 1 0 0 0 1 0 0 1 0 0 0 0 0 1 1 0 0 1 1 1 1 1 0 0 0 1 1 1 0 0 0 1 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n779, new_n780, new_n781, new_n782, new_n783, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n792, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n822, new_n823, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n874, new_n875, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n984, new_n985, new_n986, new_n987;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(KEYINPUT91), .A2(G8gat), .ZN(new_n205));
  OAI211_X1 g004(.A(new_n204), .B(new_n205), .C1(G1gat), .C2(new_n202), .ZN(new_n206));
  NOR2_X1   g005(.A1(KEYINPUT91), .A2(G8gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n206), .B(new_n207), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT87), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT14), .ZN(new_n212));
  INV_X1    g011(.A(G29gat), .ZN(new_n213));
  INV_X1    g012(.A(G36gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n210), .B1(new_n211), .B2(new_n215), .ZN(new_n216));
  NOR3_X1   g015(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT87), .ZN(new_n218));
  AOI22_X1  g017(.A1(new_n216), .A2(new_n218), .B1(G29gat), .B2(G36gat), .ZN(new_n219));
  XNOR2_X1  g018(.A(G43gat), .B(G50gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT15), .ZN(new_n221));
  XOR2_X1   g020(.A(G43gat), .B(G50gat), .Z(new_n222));
  INV_X1    g021(.A(KEYINPUT15), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(G29gat), .A2(G36gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT89), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n225), .B(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n224), .A2(new_n221), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n215), .A2(KEYINPUT88), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT88), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n217), .A2(new_n230), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n210), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  OAI22_X1  g031(.A1(new_n219), .A2(new_n221), .B1(new_n228), .B2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT90), .ZN(new_n234));
  AND3_X1   g033(.A1(new_n233), .A2(new_n234), .A3(KEYINPUT17), .ZN(new_n235));
  AOI21_X1  g034(.A(KEYINPUT17), .B1(new_n233), .B2(new_n234), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n208), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n233), .ZN(new_n238));
  OR2_X1    g037(.A1(new_n208), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(G229gat), .A2(G233gat), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n237), .A2(KEYINPUT18), .A3(new_n239), .A4(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n208), .B(new_n238), .ZN(new_n242));
  XOR2_X1   g041(.A(new_n240), .B(KEYINPUT13), .Z(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n241), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n237), .A2(new_n239), .A3(new_n240), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT18), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT92), .ZN(new_n250));
  XNOR2_X1  g049(.A(G113gat), .B(G141gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(KEYINPUT86), .B(G197gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(KEYINPUT11), .B(G169gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n255), .B(KEYINPUT12), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n246), .B(new_n249), .C1(new_n250), .C2(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n241), .A2(new_n244), .A3(new_n250), .ZN(new_n258));
  INV_X1    g057(.A(new_n256), .ZN(new_n259));
  INV_X1    g058(.A(new_n249), .ZN(new_n260));
  OAI211_X1 g059(.A(new_n258), .B(new_n259), .C1(new_n260), .C2(new_n245), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n257), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  AND2_X1   g062(.A1(KEYINPUT76), .A2(G155gat), .ZN(new_n264));
  NOR2_X1   g063(.A1(KEYINPUT76), .A2(G155gat), .ZN(new_n265));
  OAI21_X1  g064(.A(G162gat), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT2), .ZN(new_n267));
  INV_X1    g066(.A(G141gat), .ZN(new_n268));
  INV_X1    g067(.A(G148gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(G162gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(G155gat), .ZN(new_n272));
  INV_X1    g071(.A(G155gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(G162gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(G141gat), .A2(G148gat), .ZN(new_n275));
  AND4_X1   g074(.A1(new_n270), .A2(new_n272), .A3(new_n274), .A4(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT2), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n270), .A2(new_n277), .A3(new_n275), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n272), .A2(new_n274), .ZN(new_n279));
  AOI22_X1  g078(.A1(new_n267), .A2(new_n276), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT3), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT29), .ZN(new_n283));
  XOR2_X1   g082(.A(G211gat), .B(G218gat), .Z(new_n284));
  OR2_X1    g083(.A1(G197gat), .A2(G204gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(G197gat), .A2(G204gat), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT22), .ZN(new_n287));
  NAND2_X1  g086(.A1(G211gat), .A2(G218gat), .ZN(new_n288));
  AOI22_X1  g087(.A1(new_n285), .A2(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT70), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n284), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n285), .A2(new_n286), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n288), .A2(new_n287), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n284), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n294), .A2(KEYINPUT70), .A3(new_n295), .ZN(new_n296));
  AOI22_X1  g095(.A1(new_n282), .A2(new_n283), .B1(new_n291), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n296), .A2(new_n291), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n281), .B1(new_n299), .B2(KEYINPUT29), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n278), .A2(new_n279), .ZN(new_n301));
  XNOR2_X1  g100(.A(KEYINPUT76), .B(G155gat), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n277), .B1(new_n302), .B2(G162gat), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n270), .A2(new_n272), .A3(new_n274), .A4(new_n275), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n301), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n300), .A2(new_n305), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n298), .A2(new_n306), .A3(G228gat), .A4(G233gat), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT80), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n294), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n289), .A2(KEYINPUT80), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n309), .A2(new_n310), .A3(new_n284), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n295), .A2(new_n294), .A3(new_n308), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n311), .A2(new_n283), .A3(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n280), .B1(new_n313), .B2(new_n281), .ZN(new_n314));
  INV_X1    g113(.A(G228gat), .ZN(new_n315));
  INV_X1    g114(.A(G233gat), .ZN(new_n316));
  OAI22_X1  g115(.A1(new_n314), .A2(new_n297), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n307), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(G22gat), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(G78gat), .B(G106gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(KEYINPUT31), .B(G50gat), .ZN(new_n322));
  XOR2_X1   g121(.A(new_n321), .B(new_n322), .Z(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(G22gat), .B1(new_n307), .B2(new_n317), .ZN(new_n325));
  NOR3_X1   g124(.A1(new_n320), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n319), .A2(KEYINPUT81), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n323), .B1(new_n318), .B2(new_n327), .ZN(new_n328));
  OAI211_X1 g127(.A(new_n307), .B(new_n317), .C1(KEYINPUT81), .C2(new_n319), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT82), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n328), .A2(KEYINPUT82), .A3(new_n329), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n326), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(G225gat), .A2(G233gat), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT1), .ZN(new_n336));
  AND2_X1   g135(.A1(G113gat), .A2(G120gat), .ZN(new_n337));
  NOR2_X1   g136(.A1(G113gat), .A2(G120gat), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  AND2_X1   g138(.A1(G127gat), .A2(G134gat), .ZN(new_n340));
  NOR2_X1   g139(.A1(G127gat), .A2(G134gat), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT66), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n336), .B(new_n339), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(G113gat), .ZN(new_n345));
  INV_X1    g144(.A(G120gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(G113gat), .A2(G120gat), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n347), .A2(new_n336), .A3(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n347), .A2(new_n343), .A3(new_n348), .ZN(new_n350));
  XNOR2_X1  g149(.A(G127gat), .B(G134gat), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n344), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n353), .B1(new_n305), .B2(KEYINPUT3), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n335), .B1(new_n354), .B2(new_n282), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT5), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT4), .ZN(new_n359));
  AND2_X1   g158(.A1(new_n344), .A2(new_n352), .ZN(new_n360));
  OAI21_X1  g159(.A(KEYINPUT77), .B1(new_n360), .B2(new_n305), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT77), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n280), .A2(new_n353), .A3(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n359), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n280), .A2(new_n353), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(new_n359), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  NOR3_X1   g166(.A1(new_n364), .A2(KEYINPUT78), .A3(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT78), .ZN(new_n369));
  AND3_X1   g168(.A1(new_n280), .A2(new_n362), .A3(new_n353), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n362), .B1(new_n280), .B2(new_n353), .ZN(new_n371));
  OAI21_X1  g170(.A(KEYINPUT4), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n369), .B1(new_n372), .B2(new_n366), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n358), .B1(new_n368), .B2(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(G1gat), .B(G29gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n375), .B(KEYINPUT0), .ZN(new_n376));
  XNOR2_X1  g175(.A(G57gat), .B(G85gat), .ZN(new_n377));
  XOR2_X1   g176(.A(new_n376), .B(new_n377), .Z(new_n378));
  OAI211_X1 g177(.A(new_n361), .B(new_n363), .C1(new_n280), .C2(new_n353), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n356), .B1(new_n379), .B2(new_n335), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n361), .A2(new_n359), .A3(new_n363), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n381), .B(new_n355), .C1(new_n359), .C2(new_n365), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n374), .A2(new_n378), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT79), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT6), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n374), .A2(KEYINPUT79), .A3(new_n378), .A4(new_n383), .ZN(new_n388));
  AND3_X1   g187(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT85), .ZN(new_n390));
  INV_X1    g189(.A(new_n383), .ZN(new_n391));
  OAI21_X1  g190(.A(KEYINPUT78), .B1(new_n364), .B2(new_n367), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n372), .A2(new_n369), .A3(new_n366), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n357), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n390), .B1(new_n391), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n378), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n374), .A2(KEYINPUT85), .A3(new_n383), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n396), .B1(new_n391), .B2(new_n394), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  AOI22_X1  g199(.A1(new_n389), .A2(new_n398), .B1(KEYINPUT6), .B2(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(G8gat), .B(G36gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(G64gat), .B(G92gat), .ZN(new_n403));
  XOR2_X1   g202(.A(new_n402), .B(new_n403), .Z(new_n404));
  NOR2_X1   g203(.A1(G169gat), .A2(G176gat), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(KEYINPUT23), .ZN(new_n406));
  AND2_X1   g205(.A1(G169gat), .A2(G176gat), .ZN(new_n407));
  INV_X1    g206(.A(G169gat), .ZN(new_n408));
  INV_X1    g207(.A(G176gat), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT23), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n407), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(G183gat), .ZN(new_n413));
  INV_X1    g212(.A(G190gat), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT64), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n415), .B(new_n416), .C1(new_n417), .C2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(G183gat), .A2(G190gat), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT24), .ZN(new_n421));
  AND3_X1   g220(.A1(new_n420), .A2(new_n418), .A3(new_n421), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n406), .B(new_n412), .C1(new_n419), .C2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT25), .ZN(new_n424));
  INV_X1    g223(.A(new_n417), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n425), .A2(new_n415), .A3(new_n416), .ZN(new_n426));
  NAND2_X1  g225(.A1(G169gat), .A2(G176gat), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n411), .B1(G169gat), .B2(G176gat), .ZN(new_n428));
  AND4_X1   g227(.A1(KEYINPUT25), .A2(new_n406), .A3(new_n427), .A4(new_n428), .ZN(new_n429));
  AOI22_X1  g228(.A1(new_n423), .A2(new_n424), .B1(new_n426), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT26), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n410), .A2(new_n431), .A3(new_n427), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n405), .A2(KEYINPUT26), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n432), .A2(new_n420), .A3(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(KEYINPUT27), .B1(new_n413), .B2(KEYINPUT65), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT65), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT27), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n436), .A2(new_n437), .A3(G183gat), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n435), .A2(new_n438), .A3(new_n414), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT28), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  XNOR2_X1  g240(.A(KEYINPUT27), .B(G183gat), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n442), .A2(KEYINPUT28), .A3(new_n414), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n434), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(G226gat), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n445), .A2(new_n316), .ZN(new_n446));
  NOR3_X1   g245(.A1(new_n430), .A2(new_n444), .A3(new_n446), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n446), .A2(KEYINPUT29), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n429), .A2(new_n426), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n406), .A2(new_n427), .A3(new_n428), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n415), .A2(new_n416), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n418), .B1(new_n420), .B2(new_n421), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n417), .A2(new_n418), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n450), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n449), .B1(new_n455), .B2(KEYINPUT25), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n443), .ZN(new_n457));
  INV_X1    g256(.A(new_n434), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n448), .B1(new_n456), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n299), .B1(new_n447), .B2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT71), .ZN(new_n462));
  INV_X1    g261(.A(new_n448), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n463), .B1(new_n430), .B2(new_n444), .ZN(new_n464));
  INV_X1    g263(.A(new_n446), .ZN(new_n465));
  INV_X1    g264(.A(new_n452), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n466), .A2(new_n454), .A3(new_n415), .A4(new_n416), .ZN(new_n467));
  INV_X1    g266(.A(new_n450), .ZN(new_n468));
  AOI21_X1  g267(.A(KEYINPUT25), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AND2_X1   g268(.A1(new_n429), .A2(new_n426), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n459), .B(new_n465), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n299), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n464), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n461), .A2(new_n462), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n472), .B1(new_n464), .B2(new_n471), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT71), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT37), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n404), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n461), .A2(new_n473), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT38), .B1(new_n480), .B2(KEYINPUT37), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n477), .A2(new_n404), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n464), .A2(new_n472), .A3(new_n471), .ZN(new_n485));
  NOR3_X1   g284(.A1(new_n485), .A2(new_n475), .A3(KEYINPUT71), .ZN(new_n486));
  INV_X1    g285(.A(new_n476), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT72), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT72), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n474), .A2(new_n489), .A3(new_n476), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT37), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(new_n479), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n484), .B1(new_n493), .B2(KEYINPUT38), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n333), .B1(new_n401), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT84), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n392), .A2(new_n393), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n354), .A2(new_n282), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n334), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT39), .B1(new_n379), .B2(new_n335), .ZN(new_n500));
  OR2_X1    g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT39), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n396), .B1(new_n499), .B2(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n496), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT40), .ZN(new_n505));
  OR2_X1    g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n505), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n506), .A2(new_n507), .A3(new_n398), .ZN(new_n508));
  INV_X1    g307(.A(new_n404), .ZN(new_n509));
  AND3_X1   g308(.A1(new_n474), .A2(new_n489), .A3(new_n476), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n489), .B1(new_n474), .B2(new_n476), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT73), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n491), .A2(KEYINPUT73), .A3(new_n509), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT30), .ZN(new_n517));
  OAI21_X1  g316(.A(KEYINPUT74), .B1(new_n483), .B2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT74), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n477), .A2(new_n519), .A3(KEYINPUT30), .A4(new_n404), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n483), .A2(new_n517), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n516), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n495), .B1(new_n508), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n326), .ZN(new_n526));
  INV_X1    g325(.A(new_n332), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n526), .B1(new_n527), .B2(new_n330), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n528), .B(KEYINPUT83), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT75), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n530), .B1(new_n516), .B2(new_n521), .ZN(new_n531));
  AOI21_X1  g330(.A(KEYINPUT73), .B1(new_n491), .B2(new_n509), .ZN(new_n532));
  AOI211_X1 g331(.A(new_n513), .B(new_n404), .C1(new_n488), .C2(new_n490), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n530), .B(new_n521), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n522), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n386), .A2(new_n387), .A3(new_n399), .A4(new_n388), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n400), .A2(KEYINPUT6), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n534), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n529), .B1(new_n531), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(G227gat), .A2(G233gat), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n353), .B1(new_n430), .B2(new_n444), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  NOR3_X1   g342(.A1(new_n430), .A2(new_n444), .A3(new_n353), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n541), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT34), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n546), .B1(new_n541), .B2(KEYINPUT68), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n545), .B(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n430), .A2(new_n444), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(new_n360), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n551), .A2(G227gat), .A3(G233gat), .A4(new_n542), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(KEYINPUT32), .ZN(new_n553));
  XOR2_X1   g352(.A(G71gat), .B(G99gat), .Z(new_n554));
  XNOR2_X1  g353(.A(G15gat), .B(G43gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n554), .B(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT67), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT33), .ZN(new_n558));
  AND3_X1   g357(.A1(new_n552), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n557), .B1(new_n552), .B2(new_n558), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n553), .B(new_n556), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n556), .A2(KEYINPUT33), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n552), .A2(KEYINPUT32), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n549), .B1(new_n564), .B2(KEYINPUT69), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT69), .ZN(new_n566));
  AOI211_X1 g365(.A(new_n566), .B(new_n548), .C1(new_n561), .C2(new_n563), .ZN(new_n567));
  OAI21_X1  g366(.A(KEYINPUT36), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n564), .A2(new_n548), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n561), .A2(new_n549), .A3(new_n563), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n568), .B1(new_n572), .B2(KEYINPUT36), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n525), .A2(new_n540), .A3(new_n573), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n523), .A2(new_n571), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT35), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n528), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n401), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n528), .B1(new_n565), .B2(new_n567), .ZN(new_n580));
  NOR3_X1   g379(.A1(new_n539), .A2(new_n531), .A3(new_n580), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n579), .B1(new_n581), .B2(new_n576), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n263), .B1(new_n574), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT100), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT93), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(G57gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(G64gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(G71gat), .A2(G78gat), .ZN(new_n588));
  OR2_X1    g387(.A1(G71gat), .A2(G78gat), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT9), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n593));
  AND2_X1   g392(.A1(G57gat), .A2(G64gat), .ZN(new_n594));
  OAI211_X1 g393(.A(new_n588), .B(new_n589), .C1(new_n593), .C2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT21), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G127gat), .B(G155gat), .ZN(new_n599));
  XOR2_X1   g398(.A(new_n598), .B(new_n599), .Z(new_n600));
  OAI21_X1  g399(.A(new_n208), .B1(new_n597), .B2(new_n596), .ZN(new_n601));
  OR2_X1    g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(new_n601), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  XOR2_X1   g403(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT95), .ZN(new_n606));
  NAND2_X1  g405(.A1(G231gat), .A2(G233gat), .ZN(new_n607));
  XOR2_X1   g406(.A(new_n607), .B(KEYINPUT94), .Z(new_n608));
  XNOR2_X1  g407(.A(new_n606), .B(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G183gat), .B(G211gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n604), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n602), .A2(new_n603), .A3(new_n611), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(G190gat), .B(G218gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(KEYINPUT99), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(G85gat), .A2(G92gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(KEYINPUT7), .ZN(new_n621));
  NAND2_X1  g420(.A1(G99gat), .A2(G106gat), .ZN(new_n622));
  INV_X1    g421(.A(G85gat), .ZN(new_n623));
  INV_X1    g422(.A(G92gat), .ZN(new_n624));
  AOI22_X1  g423(.A1(KEYINPUT8), .A2(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT97), .ZN(new_n626));
  AND2_X1   g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n625), .A2(new_n626), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n621), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G99gat), .B(G106gat), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n629), .A2(KEYINPUT98), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n629), .A2(new_n631), .ZN(new_n633));
  OAI211_X1 g432(.A(new_n630), .B(new_n621), .C1(new_n627), .C2(new_n628), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT98), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  OAI211_X1 g435(.A(new_n632), .B(new_n636), .C1(new_n235), .C2(new_n236), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n632), .ZN(new_n638));
  AND2_X1   g437(.A1(G232gat), .A2(G233gat), .ZN(new_n639));
  AOI22_X1  g438(.A1(new_n638), .A2(new_n233), .B1(KEYINPUT41), .B2(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n619), .B1(new_n637), .B2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n639), .A2(KEYINPUT41), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(KEYINPUT96), .ZN(new_n644));
  XNOR2_X1  g443(.A(G134gat), .B(G162gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n637), .A2(new_n640), .A3(new_n619), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n642), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n646), .ZN(new_n649));
  INV_X1    g448(.A(new_n647), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n649), .B1(new_n650), .B2(new_n641), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n584), .B1(new_n616), .B2(new_n652), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n615), .A2(new_n651), .A3(KEYINPUT100), .A4(new_n648), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT10), .ZN(new_n655));
  INV_X1    g454(.A(new_n596), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n656), .A2(new_n633), .A3(new_n634), .ZN(new_n657));
  OAI211_X1 g456(.A(new_n655), .B(new_n657), .C1(new_n638), .C2(new_n656), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT101), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n596), .A2(new_n655), .ZN(new_n660));
  AND3_X1   g459(.A1(new_n638), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n659), .B1(new_n638), .B2(new_n660), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n658), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(G230gat), .A2(G233gat), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n657), .B1(new_n638), .B2(new_n656), .ZN(new_n666));
  INV_X1    g465(.A(new_n664), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(G120gat), .B(G148gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(G176gat), .B(G204gat), .ZN(new_n671));
  XOR2_X1   g470(.A(new_n670), .B(new_n671), .Z(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n665), .A2(new_n668), .A3(new_n672), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NAND4_X1  g476(.A1(new_n583), .A2(new_n653), .A3(new_n654), .A4(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n536), .A2(new_n537), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(KEYINPUT102), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n679), .A2(KEYINPUT102), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n678), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(KEYINPUT103), .B(G1gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(G1324gat));
  INV_X1    g486(.A(KEYINPUT42), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n678), .A2(new_n524), .ZN(new_n689));
  XOR2_X1   g488(.A(KEYINPUT16), .B(G8gat), .Z(new_n690));
  AOI21_X1  g489(.A(new_n688), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(G8gat), .B1(new_n678), .B2(new_n524), .ZN(new_n692));
  NOR2_X1   g491(.A1(KEYINPUT104), .A2(KEYINPUT42), .ZN(new_n693));
  MUX2_X1   g492(.A(KEYINPUT104), .B(new_n693), .S(new_n690), .Z(new_n694));
  AOI22_X1  g493(.A1(new_n691), .A2(new_n692), .B1(new_n689), .B2(new_n694), .ZN(G1325gat));
  OAI21_X1  g494(.A(G15gat), .B1(new_n678), .B2(new_n573), .ZN(new_n696));
  OR2_X1    g495(.A1(new_n571), .A2(G15gat), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n696), .B1(new_n678), .B2(new_n697), .ZN(G1326gat));
  INV_X1    g497(.A(new_n529), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n678), .A2(new_n699), .ZN(new_n700));
  XOR2_X1   g499(.A(KEYINPUT43), .B(G22gat), .Z(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(G1327gat));
  NAND2_X1  g501(.A1(new_n677), .A2(new_n616), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n703), .A2(new_n263), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n582), .A2(KEYINPUT106), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT106), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n516), .A2(new_n521), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(KEYINPUT75), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n564), .A2(KEYINPUT69), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n548), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n564), .A2(KEYINPUT69), .A3(new_n549), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n333), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n709), .A2(new_n713), .A3(new_n534), .A4(new_n538), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(KEYINPUT35), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n707), .B1(new_n715), .B2(new_n579), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n574), .B1(new_n706), .B2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n652), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n718), .A2(KEYINPUT44), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n718), .B1(new_n574), .B2(new_n582), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT44), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n705), .B1(new_n720), .B2(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n213), .B1(new_n725), .B2(new_n683), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n703), .A2(new_n718), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT105), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n583), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT45), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n683), .A2(new_n213), .ZN(new_n731));
  OR3_X1    g530(.A1(new_n729), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n730), .B1(new_n729), .B2(new_n731), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(KEYINPUT107), .B1(new_n726), .B2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n574), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n582), .A2(KEYINPUT106), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n715), .A2(new_n707), .A3(new_n579), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(new_n719), .ZN(new_n740));
  OAI22_X1  g539(.A1(new_n739), .A2(new_n740), .B1(new_n722), .B2(new_n721), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(new_n704), .ZN(new_n742));
  OAI21_X1  g541(.A(G29gat), .B1(new_n742), .B2(new_n684), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT107), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n743), .A2(new_n744), .A3(new_n733), .A4(new_n732), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n735), .A2(new_n745), .ZN(G1328gat));
  NOR3_X1   g545(.A1(new_n729), .A2(G36gat), .A3(new_n524), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT46), .ZN(new_n748));
  OAI21_X1  g547(.A(G36gat), .B1(new_n742), .B2(new_n524), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(G1329gat));
  INV_X1    g549(.A(G43gat), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n751), .B1(new_n729), .B2(new_n571), .ZN(new_n752));
  OR2_X1    g551(.A1(new_n573), .A2(new_n751), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n752), .B1(new_n742), .B2(new_n753), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g554(.A1(new_n737), .A2(new_n738), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n740), .B1(new_n756), .B2(new_n574), .ZN(new_n757));
  OAI211_X1 g556(.A(new_n333), .B(new_n704), .C1(new_n757), .C2(new_n723), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(KEYINPUT110), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT110), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n741), .A2(new_n760), .A3(new_n333), .A4(new_n704), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n759), .A2(G50gat), .A3(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(G50gat), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n529), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n729), .A2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT48), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n762), .A2(new_n767), .ZN(new_n768));
  XOR2_X1   g567(.A(KEYINPUT108), .B(KEYINPUT48), .Z(new_n769));
  AOI21_X1  g568(.A(new_n763), .B1(new_n725), .B2(new_n529), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n765), .B(KEYINPUT109), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n768), .A2(new_n772), .ZN(G1331gat));
  AND4_X1   g572(.A1(new_n263), .A2(new_n653), .A3(new_n654), .A4(new_n676), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n717), .A2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(new_n683), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g577(.A(KEYINPUT49), .B(G64gat), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n776), .A2(new_n523), .A3(new_n779), .ZN(new_n780));
  OAI22_X1  g579(.A1(new_n775), .A2(new_n524), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT111), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n782), .B(new_n783), .ZN(G1333gat));
  XNOR2_X1  g583(.A(new_n571), .B(KEYINPUT112), .ZN(new_n785));
  AOI21_X1  g584(.A(G71gat), .B1(new_n776), .B2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(G71gat), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n775), .A2(new_n787), .A3(new_n573), .ZN(new_n788));
  OR3_X1    g587(.A1(new_n786), .A2(new_n788), .A3(KEYINPUT50), .ZN(new_n789));
  OAI21_X1  g588(.A(KEYINPUT50), .B1(new_n786), .B2(new_n788), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(G1334gat));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n529), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n792), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g592(.A1(new_n262), .A2(new_n615), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(KEYINPUT113), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n676), .ZN(new_n796));
  XOR2_X1   g595(.A(new_n796), .B(KEYINPUT114), .Z(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n798), .B1(new_n720), .B2(new_n724), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(G85gat), .B1(new_n800), .B2(new_n684), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT51), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n795), .A2(new_n652), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n802), .B1(new_n739), .B2(new_n803), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n717), .A2(KEYINPUT51), .A3(new_n652), .A4(new_n795), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT115), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n739), .A2(new_n803), .ZN(new_n808));
  AOI21_X1  g607(.A(KEYINPUT115), .B1(new_n808), .B2(KEYINPUT51), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n683), .A2(new_n623), .A3(new_n676), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n801), .B1(new_n810), .B2(new_n811), .ZN(G1336gat));
  NAND3_X1  g611(.A1(new_n741), .A2(new_n523), .A3(new_n797), .ZN(new_n813));
  AOI21_X1  g612(.A(KEYINPUT52), .B1(new_n813), .B2(G92gat), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n524), .A2(G92gat), .A3(new_n677), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n814), .B1(new_n810), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n624), .B1(new_n799), .B2(new_n523), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n816), .B1(new_n804), .B2(new_n805), .ZN(new_n819));
  OAI21_X1  g618(.A(KEYINPUT52), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n817), .A2(new_n820), .ZN(G1337gat));
  OAI21_X1  g620(.A(G99gat), .B1(new_n800), .B2(new_n573), .ZN(new_n822));
  OR3_X1    g621(.A1(new_n677), .A2(new_n571), .A3(G99gat), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n822), .B1(new_n810), .B2(new_n823), .ZN(G1338gat));
  NAND3_X1  g623(.A1(new_n741), .A2(new_n333), .A3(new_n797), .ZN(new_n825));
  AOI21_X1  g624(.A(KEYINPUT53), .B1(new_n825), .B2(G106gat), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n677), .A2(new_n528), .A3(G106gat), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n826), .B1(new_n810), .B2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(G106gat), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n830), .B1(new_n799), .B2(new_n529), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n828), .B1(new_n804), .B2(new_n805), .ZN(new_n832));
  OAI21_X1  g631(.A(KEYINPUT53), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n829), .A2(new_n833), .ZN(G1339gat));
  NAND4_X1  g633(.A1(new_n653), .A2(new_n263), .A3(new_n677), .A4(new_n654), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT116), .ZN(new_n836));
  XNOR2_X1  g635(.A(new_n835), .B(new_n836), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n667), .B(new_n658), .C1(new_n661), .C2(new_n662), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n665), .A2(KEYINPUT54), .A3(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT54), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n663), .A2(new_n840), .A3(new_n664), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n839), .A2(KEYINPUT55), .A3(new_n673), .A4(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(KEYINPUT117), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n841), .A2(new_n673), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT117), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n845), .A2(new_n846), .A3(KEYINPUT55), .A4(new_n839), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n843), .A2(new_n847), .A3(new_n675), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT55), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n665), .A2(KEYINPUT54), .A3(new_n838), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n849), .B1(new_n850), .B2(new_n844), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n260), .A2(new_n245), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n237), .A2(new_n239), .ZN(new_n853));
  OAI22_X1  g652(.A1(new_n853), .A2(new_n240), .B1(new_n242), .B2(new_n243), .ZN(new_n854));
  AOI22_X1  g653(.A1(new_n852), .A2(new_n256), .B1(new_n255), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n851), .A2(new_n652), .A3(new_n855), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n848), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n855), .A2(new_n676), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n851), .A2(new_n262), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n858), .B1(new_n848), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n857), .B1(new_n860), .B2(new_n718), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n837), .B1(new_n861), .B2(new_n615), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n862), .A2(new_n699), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n863), .A2(new_n575), .A3(new_n683), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n864), .A2(new_n345), .A3(new_n263), .ZN(new_n865));
  AND3_X1   g664(.A1(new_n862), .A2(new_n524), .A3(new_n683), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(new_n713), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(new_n262), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n865), .B1(new_n869), .B2(new_n345), .ZN(G1340gat));
  NOR3_X1   g669(.A1(new_n864), .A2(new_n346), .A3(new_n677), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n868), .A2(new_n676), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n871), .B1(new_n872), .B2(new_n346), .ZN(G1341gat));
  OAI21_X1  g672(.A(G127gat), .B1(new_n864), .B2(new_n616), .ZN(new_n874));
  OR2_X1    g673(.A1(new_n616), .A2(G127gat), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n874), .B1(new_n867), .B2(new_n875), .ZN(G1342gat));
  NOR2_X1   g675(.A1(new_n718), .A2(G134gat), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  OR3_X1    g677(.A1(new_n867), .A2(KEYINPUT56), .A3(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(G134gat), .B1(new_n864), .B2(new_n718), .ZN(new_n880));
  OAI21_X1  g679(.A(KEYINPUT56), .B1(new_n867), .B2(new_n878), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(G1343gat));
  NAND2_X1  g681(.A1(new_n573), .A2(new_n333), .ZN(new_n883));
  XNOR2_X1  g682(.A(new_n883), .B(KEYINPUT118), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n866), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n885), .A2(new_n268), .A3(new_n262), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT57), .ZN(new_n887));
  AND3_X1   g686(.A1(new_n862), .A2(new_n887), .A3(new_n333), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n887), .B1(new_n862), .B2(new_n529), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n683), .A2(new_n524), .A3(new_n573), .ZN(new_n890));
  NOR4_X1   g689(.A1(new_n888), .A2(new_n889), .A3(new_n263), .A4(new_n890), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n886), .B1(new_n891), .B2(new_n268), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(KEYINPUT58), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT58), .ZN(new_n894));
  OAI211_X1 g693(.A(new_n886), .B(new_n894), .C1(new_n268), .C2(new_n891), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n893), .A2(new_n895), .ZN(G1344gat));
  NAND3_X1  g695(.A1(new_n885), .A2(new_n269), .A3(new_n676), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT59), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n890), .A2(new_n677), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n862), .A2(KEYINPUT57), .A3(new_n333), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT119), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n862), .A2(KEYINPUT119), .A3(KEYINPUT57), .A4(new_n333), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n835), .B1(new_n861), .B2(new_n615), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT120), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n699), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n860), .A2(new_n718), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n616), .B1(new_n908), .B2(new_n857), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n909), .A2(KEYINPUT120), .A3(new_n835), .ZN(new_n910));
  AOI21_X1  g709(.A(KEYINPUT57), .B1(new_n907), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n899), .B1(new_n904), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n898), .B1(new_n912), .B2(G148gat), .ZN(new_n913));
  NOR3_X1   g712(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n914));
  AOI211_X1 g713(.A(KEYINPUT59), .B(new_n269), .C1(new_n914), .C2(new_n676), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n897), .B1(new_n913), .B2(new_n915), .ZN(G1345gat));
  INV_X1    g715(.A(new_n914), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n302), .B1(new_n917), .B2(new_n616), .ZN(new_n918));
  INV_X1    g717(.A(new_n302), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n885), .A2(new_n919), .A3(new_n615), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n920), .ZN(G1346gat));
  NAND3_X1  g720(.A1(new_n885), .A2(new_n271), .A3(new_n652), .ZN(new_n922));
  OAI21_X1  g721(.A(KEYINPUT121), .B1(new_n917), .B2(new_n718), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(G162gat), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n917), .A2(KEYINPUT121), .A3(new_n718), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n922), .B1(new_n924), .B2(new_n925), .ZN(G1347gat));
  AND2_X1   g725(.A1(new_n862), .A2(new_n684), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n713), .A2(new_n523), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n928), .B(KEYINPUT122), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(G169gat), .B1(new_n930), .B2(new_n262), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n683), .A2(new_n524), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(new_n785), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n863), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n263), .A2(new_n408), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n931), .B1(new_n935), .B2(new_n936), .ZN(G1348gat));
  NAND2_X1  g736(.A1(new_n930), .A2(new_n676), .ZN(new_n938));
  AND3_X1   g737(.A1(new_n938), .A2(KEYINPUT123), .A3(new_n409), .ZN(new_n939));
  NAND4_X1  g738(.A1(new_n863), .A2(G176gat), .A3(new_n676), .A4(new_n934), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT124), .ZN(new_n941));
  AOI21_X1  g740(.A(KEYINPUT123), .B1(new_n938), .B2(new_n409), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n939), .A2(new_n941), .A3(new_n942), .ZN(G1349gat));
  NAND3_X1  g742(.A1(new_n863), .A2(new_n615), .A3(new_n934), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT125), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND4_X1  g745(.A1(new_n863), .A2(KEYINPUT125), .A3(new_n615), .A4(new_n934), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n946), .A2(new_n947), .A3(G183gat), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n930), .A2(new_n442), .A3(new_n615), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(KEYINPUT60), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT60), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n948), .A2(new_n949), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n951), .A2(new_n953), .ZN(G1350gat));
  NAND3_X1  g753(.A1(new_n930), .A2(new_n414), .A3(new_n652), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT126), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n955), .B(new_n956), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n935), .A2(new_n652), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(G190gat), .ZN(new_n959));
  XNOR2_X1  g758(.A(KEYINPUT127), .B(KEYINPUT61), .ZN(new_n960));
  OR2_X1    g759(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n959), .A2(new_n960), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n957), .A2(new_n961), .A3(new_n962), .ZN(G1351gat));
  NAND2_X1  g762(.A1(new_n932), .A2(new_n573), .ZN(new_n964));
  INV_X1    g763(.A(new_n964), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n262), .A2(G197gat), .ZN(new_n966));
  OAI211_X1 g765(.A(new_n965), .B(new_n966), .C1(new_n904), .C2(new_n911), .ZN(new_n967));
  INV_X1    g766(.A(new_n967), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n883), .A2(new_n524), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n927), .A2(new_n969), .ZN(new_n970));
  INV_X1    g769(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g770(.A(G197gat), .B1(new_n971), .B2(new_n262), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n968), .A2(new_n972), .ZN(G1352gat));
  NOR3_X1   g772(.A1(new_n970), .A2(G204gat), .A3(new_n677), .ZN(new_n974));
  XNOR2_X1  g773(.A(new_n974), .B(KEYINPUT62), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n965), .B1(new_n904), .B2(new_n911), .ZN(new_n976));
  OAI21_X1  g775(.A(G204gat), .B1(new_n976), .B2(new_n677), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n975), .A2(new_n977), .ZN(G1353gat));
  OR3_X1    g777(.A1(new_n970), .A2(G211gat), .A3(new_n616), .ZN(new_n979));
  OAI211_X1 g778(.A(new_n615), .B(new_n965), .C1(new_n904), .C2(new_n911), .ZN(new_n980));
  AND3_X1   g779(.A1(new_n980), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n981));
  AOI21_X1  g780(.A(KEYINPUT63), .B1(new_n980), .B2(G211gat), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n979), .B1(new_n981), .B2(new_n982), .ZN(G1354gat));
  INV_X1    g782(.A(G218gat), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n971), .A2(new_n984), .A3(new_n652), .ZN(new_n985));
  OAI211_X1 g784(.A(new_n652), .B(new_n965), .C1(new_n904), .C2(new_n911), .ZN(new_n986));
  INV_X1    g785(.A(new_n986), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n985), .B1(new_n987), .B2(new_n984), .ZN(G1355gat));
endmodule


