//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 1 0 1 0 0 1 1 0 0 0 0 1 0 1 0 0 1 1 0 1 1 0 1 1 0 0 0 1 1 0 0 1 0 0 1 0 0 1 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:54 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  XOR2_X1   g001(.A(new_n187), .B(KEYINPUT74), .Z(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT11), .ZN(new_n190));
  INV_X1    g004(.A(G134), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n190), .B1(new_n191), .B2(G137), .ZN(new_n192));
  INV_X1    g006(.A(G137), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n193), .A2(KEYINPUT11), .A3(G134), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n191), .A2(G137), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n192), .A2(new_n194), .A3(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G131), .ZN(new_n197));
  INV_X1    g011(.A(G131), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n192), .A2(new_n194), .A3(new_n198), .A4(new_n195), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G143), .ZN(new_n202));
  INV_X1    g016(.A(G143), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G146), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(KEYINPUT0), .A2(G128), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT64), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT0), .ZN(new_n208));
  INV_X1    g022(.A(G128), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n205), .A2(new_n206), .A3(new_n210), .A4(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT65), .ZN(new_n213));
  XNOR2_X1  g027(.A(G143), .B(G146), .ZN(new_n214));
  INV_X1    g028(.A(new_n206), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n212), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n211), .ZN(new_n218));
  NOR3_X1   g032(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n220), .A2(new_n213), .A3(new_n205), .A4(new_n206), .ZN(new_n221));
  AND3_X1   g035(.A1(new_n217), .A2(KEYINPUT70), .A3(new_n221), .ZN(new_n222));
  AOI21_X1  g036(.A(KEYINPUT70), .B1(new_n217), .B2(new_n221), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n200), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n193), .A2(G134), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(new_n195), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G131), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(KEYINPUT66), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n226), .A2(new_n229), .A3(G131), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n228), .A2(new_n199), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT71), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n228), .A2(KEYINPUT71), .A3(new_n230), .A4(new_n199), .ZN(new_n234));
  AND2_X1   g048(.A1(KEYINPUT67), .A2(G128), .ZN(new_n235));
  NOR2_X1   g049(.A1(KEYINPUT67), .A2(G128), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT1), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n238), .B1(G143), .B2(new_n201), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n205), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n202), .A2(new_n204), .A3(new_n238), .A4(G128), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n233), .A2(new_n234), .A3(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT69), .ZN(new_n244));
  NAND2_X1  g058(.A1(KEYINPUT2), .A2(G113), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(KEYINPUT68), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT68), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n247), .A2(KEYINPUT2), .A3(G113), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT2), .ZN(new_n250));
  INV_X1    g064(.A(G113), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G119), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G116), .ZN(new_n255));
  INV_X1    g069(.A(G116), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G119), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n253), .A2(new_n258), .ZN(new_n259));
  AOI22_X1  g073(.A1(new_n246), .A2(new_n248), .B1(new_n250), .B2(new_n251), .ZN(new_n260));
  INV_X1    g074(.A(new_n258), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n244), .B1(new_n259), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n253), .A2(new_n258), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n260), .A2(new_n261), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n264), .A2(KEYINPUT69), .A3(new_n265), .ZN(new_n266));
  AND2_X1   g080(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n224), .A2(new_n243), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(KEYINPUT72), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT72), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n224), .A2(new_n267), .A3(new_n243), .A4(new_n270), .ZN(new_n271));
  AND2_X1   g085(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n224), .A2(KEYINPUT30), .A3(new_n243), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n263), .A2(new_n266), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n217), .A2(new_n221), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(new_n200), .ZN(new_n276));
  AND2_X1   g090(.A1(new_n240), .A2(new_n241), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n276), .B1(new_n231), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT30), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n273), .A2(new_n274), .A3(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G237), .ZN(new_n282));
  INV_X1    g096(.A(G953), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n282), .A2(new_n283), .A3(G210), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n284), .B(KEYINPUT27), .ZN(new_n285));
  XNOR2_X1  g099(.A(KEYINPUT26), .B(G101), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n285), .B(new_n286), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n272), .A2(KEYINPUT73), .A3(new_n281), .A4(new_n287), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n281), .A2(new_n269), .A3(new_n271), .A4(new_n287), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT73), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AND3_X1   g105(.A1(new_n288), .A2(KEYINPUT31), .A3(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT28), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n268), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n278), .A2(new_n274), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n269), .A2(new_n271), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n295), .B1(new_n297), .B2(KEYINPUT28), .ZN(new_n298));
  OAI22_X1  g112(.A1(new_n298), .A2(new_n287), .B1(KEYINPUT31), .B2(new_n289), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n189), .B1(new_n292), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(KEYINPUT75), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT32), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n289), .A2(KEYINPUT31), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n297), .A2(KEYINPUT28), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n294), .ZN(new_n305));
  INV_X1    g119(.A(new_n287), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n303), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n288), .A2(KEYINPUT31), .A3(new_n291), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT75), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n309), .A2(new_n310), .A3(new_n189), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n301), .A2(new_n302), .A3(new_n311), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n188), .A2(new_n302), .ZN(new_n313));
  AOI21_X1  g127(.A(KEYINPUT76), .B1(new_n309), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT76), .ZN(new_n315));
  INV_X1    g129(.A(new_n313), .ZN(new_n316));
  AOI211_X1 g130(.A(new_n315), .B(new_n316), .C1(new_n307), .C2(new_n308), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n281), .A2(new_n269), .A3(new_n271), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(new_n306), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT29), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n322), .B1(new_n287), .B2(new_n298), .ZN(new_n323));
  INV_X1    g137(.A(G902), .ZN(new_n324));
  AND2_X1   g138(.A1(new_n224), .A2(new_n243), .ZN(new_n325));
  OAI211_X1 g139(.A(new_n269), .B(new_n271), .C1(new_n325), .C2(new_n267), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(KEYINPUT28), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(new_n294), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n287), .A2(KEYINPUT29), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n324), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(G472), .B1(new_n323), .B2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n312), .A2(new_n318), .A3(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G140), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n333), .A2(KEYINPUT78), .A3(G125), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(G125), .ZN(new_n335));
  INV_X1    g149(.A(G125), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(G140), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  OAI211_X1 g152(.A(KEYINPUT16), .B(new_n334), .C1(new_n338), .C2(KEYINPUT78), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT16), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n335), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G146), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n338), .A2(G146), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  XOR2_X1   g159(.A(KEYINPUT24), .B(G110), .Z(new_n346));
  NOR3_X1   g160(.A1(new_n235), .A2(new_n236), .A3(new_n254), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n209), .A2(G119), .ZN(new_n348));
  OAI21_X1  g162(.A(KEYINPUT77), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT67), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n209), .ZN(new_n351));
  NAND2_X1  g165(.A1(KEYINPUT67), .A2(G128), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n351), .A2(G119), .A3(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT77), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n353), .B(new_n354), .C1(G119), .C2(new_n209), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n346), .B1(new_n349), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n347), .A2(KEYINPUT23), .ZN(new_n357));
  INV_X1    g171(.A(G110), .ZN(new_n358));
  AOI21_X1  g172(.A(KEYINPUT23), .B1(new_n209), .B2(G119), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n359), .A2(new_n348), .ZN(new_n360));
  AND3_X1   g174(.A1(new_n357), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n343), .B(new_n345), .C1(new_n356), .C2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT79), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n201), .B1(new_n339), .B2(new_n341), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n365), .A2(new_n344), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n366), .B(KEYINPUT79), .C1(new_n361), .C2(new_n356), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n349), .A2(new_n355), .A3(new_n346), .ZN(new_n368));
  AND2_X1   g182(.A1(new_n357), .A2(new_n360), .ZN(new_n369));
  AND3_X1   g183(.A1(new_n339), .A2(new_n201), .A3(new_n341), .ZN(new_n370));
  OAI221_X1 g184(.A(new_n368), .B1(new_n369), .B2(new_n358), .C1(new_n370), .C2(new_n365), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n364), .A2(new_n367), .A3(new_n371), .ZN(new_n372));
  XNOR2_X1  g186(.A(KEYINPUT22), .B(G137), .ZN(new_n373));
  AND3_X1   g187(.A1(new_n283), .A2(G221), .A3(G234), .ZN(new_n374));
  XOR2_X1   g188(.A(new_n373), .B(new_n374), .Z(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n372), .A2(new_n376), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n364), .A2(new_n367), .A3(new_n371), .A4(new_n375), .ZN(new_n378));
  AND2_X1   g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G217), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n380), .B1(G234), .B2(new_n324), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n381), .A2(G902), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n377), .A2(new_n324), .A3(new_n378), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT25), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n377), .A2(KEYINPUT25), .A3(new_n324), .A4(new_n378), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n386), .A2(KEYINPUT80), .A3(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n381), .B1(new_n386), .B2(KEYINPUT80), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n383), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT20), .ZN(new_n392));
  XNOR2_X1  g206(.A(G113), .B(G122), .ZN(new_n393));
  INV_X1    g207(.A(G104), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n393), .B(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n282), .A2(new_n283), .A3(G214), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n396), .B(G143), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT18), .ZN(new_n398));
  OR3_X1    g212(.A1(new_n397), .A2(new_n398), .A3(new_n198), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n334), .B1(new_n338), .B2(KEYINPUT78), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n345), .B1(new_n400), .B2(new_n201), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n397), .B1(new_n398), .B2(new_n198), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n399), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n339), .A2(new_n201), .A3(new_n341), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n343), .A2(new_n404), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n397), .A2(new_n198), .ZN(new_n406));
  AOI22_X1  g220(.A1(new_n405), .A2(KEYINPUT88), .B1(KEYINPUT17), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT88), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n343), .A2(new_n408), .A3(new_n404), .ZN(new_n409));
  AOI21_X1  g223(.A(KEYINPUT89), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(KEYINPUT88), .B1(new_n370), .B2(new_n365), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n406), .A2(KEYINPUT17), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n411), .A2(new_n409), .A3(KEYINPUT89), .A4(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n397), .B(new_n198), .ZN(new_n414));
  OR2_X1    g228(.A1(new_n414), .A2(KEYINPUT17), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n395), .B(new_n403), .C1(new_n410), .C2(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(KEYINPUT19), .B1(new_n335), .B2(new_n337), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n418), .B1(new_n400), .B2(KEYINPUT19), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n414), .B(new_n343), .C1(G146), .C2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n403), .ZN(new_n421));
  INV_X1    g235(.A(new_n395), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n417), .A2(new_n423), .ZN(new_n424));
  NOR2_X1   g238(.A1(G475), .A2(G902), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n392), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n425), .ZN(new_n427));
  AOI211_X1 g241(.A(KEYINPUT20), .B(new_n427), .C1(new_n417), .C2(new_n423), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n403), .B1(new_n410), .B2(new_n416), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n422), .ZN(new_n430));
  AOI21_X1  g244(.A(G902), .B1(new_n430), .B2(new_n417), .ZN(new_n431));
  INV_X1    g245(.A(G475), .ZN(new_n432));
  OAI22_X1  g246(.A1(new_n426), .A2(new_n428), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  XNOR2_X1  g248(.A(G110), .B(G122), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT85), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n256), .A2(G119), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT5), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n251), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n255), .A2(new_n257), .A3(KEYINPUT5), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n265), .A2(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(KEYINPUT3), .B1(new_n394), .B2(G107), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT3), .ZN(new_n445));
  INV_X1    g259(.A(G107), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n445), .A2(new_n446), .A3(G104), .ZN(new_n447));
  INV_X1    g261(.A(G101), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n394), .A2(G107), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n444), .A2(new_n447), .A3(new_n448), .A4(new_n449), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n394), .A2(G107), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n446), .A2(G104), .ZN(new_n452));
  OAI21_X1  g266(.A(G101), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n437), .B1(new_n443), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n454), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n456), .A2(KEYINPUT85), .A3(new_n265), .A4(new_n442), .ZN(new_n457));
  AND2_X1   g271(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n444), .A2(new_n447), .A3(new_n449), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(G101), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n460), .A2(KEYINPUT4), .A3(new_n450), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT4), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n459), .A2(new_n462), .A3(G101), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n464), .B1(new_n263), .B2(new_n266), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n436), .B1(new_n458), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n455), .A2(new_n457), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n435), .B(new_n467), .C1(new_n267), .C2(new_n464), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n466), .A2(new_n468), .A3(KEYINPUT6), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT6), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n470), .B(new_n436), .C1(new_n458), .C2(new_n465), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n275), .A2(G125), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n242), .A2(new_n336), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(KEYINPUT86), .B(G224), .ZN(new_n475));
  OR2_X1    g289(.A1(new_n475), .A2(G953), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n474), .B(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n469), .A2(new_n471), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n476), .A2(KEYINPUT7), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n474), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n472), .A2(new_n473), .A3(new_n479), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n454), .A2(new_n265), .A3(new_n442), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n435), .B(KEYINPUT8), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT87), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n441), .A2(new_n485), .ZN(new_n486));
  AND2_X1   g300(.A1(new_n486), .A2(new_n440), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n261), .A2(KEYINPUT87), .A3(KEYINPUT5), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n259), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n483), .B(new_n484), .C1(new_n489), .C2(new_n454), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n481), .A2(new_n482), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(G902), .B1(new_n491), .B2(new_n468), .ZN(new_n492));
  OAI21_X1  g306(.A(G210), .B1(G237), .B2(G902), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n478), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n493), .B1(new_n478), .B2(new_n492), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(G952), .ZN(new_n498));
  AOI211_X1 g312(.A(G953), .B(new_n498), .C1(G234), .C2(G237), .ZN(new_n499));
  NAND2_X1  g313(.A1(G234), .A2(G237), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n500), .A2(G902), .A3(G953), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n501), .B(KEYINPUT93), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(KEYINPUT21), .B(G898), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n499), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(G214), .B1(G237), .B2(G902), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  NOR3_X1   g321(.A1(new_n497), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(G478), .ZN(new_n509));
  OR2_X1    g323(.A1(new_n509), .A2(KEYINPUT15), .ZN(new_n510));
  XNOR2_X1  g324(.A(KEYINPUT9), .B(G234), .ZN(new_n511));
  NOR3_X1   g325(.A1(new_n511), .A2(new_n380), .A3(G953), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n351), .A2(G143), .A3(new_n352), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n203), .A2(G128), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT13), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n203), .A2(KEYINPUT13), .A3(G128), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n513), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(G122), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(G116), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n256), .A2(G122), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(G107), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n520), .A2(new_n521), .A3(new_n446), .ZN(new_n524));
  AOI22_X1  g338(.A1(new_n518), .A2(G134), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n513), .A2(new_n191), .A3(new_n514), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n519), .A2(G116), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT14), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n520), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n529), .A2(new_n530), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n531), .B1(KEYINPUT90), .B2(new_n532), .ZN(new_n533));
  OR2_X1    g347(.A1(new_n532), .A2(KEYINPUT90), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n446), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n191), .B1(new_n513), .B2(new_n514), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n524), .B1(new_n526), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n528), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT91), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n528), .B(KEYINPUT91), .C1(new_n535), .C2(new_n537), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n512), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n512), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n544), .B1(new_n538), .B2(new_n539), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(G902), .B1(new_n543), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT92), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AOI211_X1 g363(.A(KEYINPUT92), .B(G902), .C1(new_n543), .C2(new_n546), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n510), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  OR2_X1    g365(.A1(new_n550), .A2(new_n510), .ZN(new_n552));
  AND2_X1   g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(G221), .B1(new_n511), .B2(G902), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n283), .A2(G227), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n556), .B(KEYINPUT81), .ZN(new_n557));
  XNOR2_X1  g371(.A(G110), .B(G140), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n557), .B(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n200), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n277), .A2(new_n454), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT82), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n241), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n214), .A2(KEYINPUT82), .A3(new_n238), .A4(G128), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n205), .B1(new_n239), .B2(new_n209), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n456), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n561), .B1(new_n562), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n569), .B1(KEYINPUT83), .B2(KEYINPUT12), .ZN(new_n570));
  XOR2_X1   g384(.A(KEYINPUT83), .B(KEYINPUT12), .Z(new_n571));
  OAI21_X1  g385(.A(new_n570), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  AND2_X1   g386(.A1(new_n461), .A2(new_n463), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n573), .B1(new_n222), .B2(new_n223), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT10), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n575), .B1(new_n240), .B2(new_n241), .ZN(new_n576));
  AOI22_X1  g390(.A1(new_n568), .A2(new_n575), .B1(new_n456), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n574), .A2(new_n577), .A3(new_n561), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n560), .B1(new_n572), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n574), .A2(new_n577), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n200), .ZN(new_n581));
  AND3_X1   g395(.A1(new_n581), .A2(new_n578), .A3(new_n560), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(G469), .B1(new_n583), .B2(G902), .ZN(new_n584));
  INV_X1    g398(.A(G469), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT84), .ZN(new_n586));
  AND3_X1   g400(.A1(new_n578), .A2(new_n586), .A3(new_n560), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n586), .B1(new_n578), .B2(new_n560), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n569), .A2(new_n571), .ZN(new_n589));
  NOR2_X1   g403(.A1(KEYINPUT83), .A2(KEYINPUT12), .ZN(new_n590));
  AOI211_X1 g404(.A(new_n590), .B(new_n561), .C1(new_n562), .C2(new_n568), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NOR3_X1   g406(.A1(new_n587), .A2(new_n588), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n560), .B1(new_n581), .B2(new_n578), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n585), .B(new_n324), .C1(new_n593), .C2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n555), .B1(new_n584), .B2(new_n595), .ZN(new_n596));
  AND4_X1   g410(.A1(new_n434), .A2(new_n508), .A3(new_n553), .A4(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n332), .A2(new_n391), .A3(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(G101), .ZN(G3));
  INV_X1    g413(.A(G472), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n600), .B1(new_n309), .B2(new_n324), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(KEYINPUT94), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT94), .ZN(new_n603));
  AOI21_X1  g417(.A(G902), .B1(new_n307), .B2(new_n308), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n603), .B1(new_n604), .B2(new_n600), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  AND2_X1   g420(.A1(new_n301), .A2(new_n311), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n584), .A2(new_n595), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n554), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n608), .A2(new_n390), .A3(new_n610), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n544), .A2(KEYINPUT98), .ZN(new_n612));
  OR2_X1    g426(.A1(new_n538), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n538), .A2(new_n612), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n613), .A2(KEYINPUT33), .A3(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(KEYINPUT96), .B(KEYINPUT33), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n617), .B1(new_n542), .B2(new_n545), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT97), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI211_X1 g434(.A(KEYINPUT97), .B(new_n617), .C1(new_n542), .C2(new_n545), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n616), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n509), .A2(G902), .ZN(new_n623));
  INV_X1    g437(.A(new_n547), .ZN(new_n624));
  AOI22_X1  g438(.A1(new_n622), .A2(new_n623), .B1(new_n509), .B2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n431), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(G475), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n424), .A2(new_n425), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(KEYINPUT20), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n424), .A2(new_n392), .A3(new_n425), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n625), .B1(new_n627), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n478), .A2(new_n492), .ZN(new_n633));
  INV_X1    g447(.A(new_n493), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n635), .A2(KEYINPUT95), .A3(new_n494), .ZN(new_n636));
  INV_X1    g450(.A(new_n505), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT95), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n507), .B1(new_n496), .B2(new_n638), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n636), .A2(new_n637), .A3(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n611), .A2(new_n632), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT34), .B(G104), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G6));
  NOR2_X1   g457(.A1(new_n553), .A2(new_n433), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n611), .A2(new_n640), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT35), .B(G107), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G9));
  NOR2_X1   g461(.A1(new_n376), .A2(KEYINPUT36), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(KEYINPUT99), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n372), .B(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n382), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n651), .B1(new_n388), .B2(new_n389), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n606), .A2(new_n597), .A3(new_n607), .A4(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT37), .B(G110), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G12));
  AND2_X1   g469(.A1(new_n636), .A2(new_n639), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n656), .A2(new_n596), .A3(new_n652), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n551), .A2(new_n552), .ZN(new_n658));
  XNOR2_X1  g472(.A(KEYINPUT100), .B(G900), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n503), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n499), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n434), .A2(new_n658), .A3(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n657), .A2(new_n663), .ZN(new_n664));
  AND3_X1   g478(.A1(new_n301), .A2(new_n302), .A3(new_n311), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n313), .B1(new_n292), .B2(new_n299), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n315), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n309), .A2(KEYINPUT76), .A3(new_n313), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n667), .A2(new_n668), .A3(new_n331), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n664), .B1(new_n665), .B2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G128), .ZN(G30));
  XOR2_X1   g485(.A(new_n497), .B(KEYINPUT38), .Z(new_n672));
  NAND2_X1  g486(.A1(new_n658), .A2(new_n433), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n672), .A2(new_n506), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n662), .B(KEYINPUT39), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n596), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n677), .A2(KEYINPUT40), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n677), .A2(KEYINPUT40), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n675), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n288), .A2(new_n291), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n326), .A2(new_n306), .ZN(new_n682));
  AOI21_X1  g496(.A(KEYINPUT101), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n288), .A2(KEYINPUT101), .A3(new_n291), .A4(new_n682), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n324), .ZN(new_n685));
  OAI21_X1  g499(.A(G472), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n686), .A2(new_n667), .A3(new_n668), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(new_n312), .ZN(new_n689));
  INV_X1    g503(.A(new_n652), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n680), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G143), .ZN(G45));
  NAND2_X1  g506(.A1(new_n620), .A2(new_n621), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n693), .A2(new_n615), .A3(new_n623), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n624), .A2(new_n509), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n433), .A2(new_n696), .A3(new_n662), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n657), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n698), .B1(new_n665), .B2(new_n669), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G146), .ZN(G48));
  NAND2_X1  g514(.A1(new_n578), .A2(new_n560), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n592), .B1(new_n701), .B2(KEYINPUT84), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n578), .A2(new_n586), .A3(new_n560), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n594), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  OAI21_X1  g518(.A(G469), .B1(new_n704), .B2(G902), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n705), .A2(new_n554), .A3(new_n595), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n390), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n707), .A2(new_n632), .A3(new_n640), .ZN(new_n708));
  AND3_X1   g522(.A1(new_n667), .A2(new_n668), .A3(new_n331), .ZN(new_n709));
  AOI211_X1 g523(.A(KEYINPUT102), .B(new_n708), .C1(new_n709), .C2(new_n312), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT102), .ZN(new_n711));
  INV_X1    g525(.A(new_n708), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n711), .B1(new_n332), .B2(new_n712), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  XOR2_X1   g528(.A(KEYINPUT41), .B(G113), .Z(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G15));
  AND3_X1   g530(.A1(new_n644), .A2(new_n707), .A3(new_n640), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n717), .B1(new_n665), .B2(new_n669), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G116), .ZN(G18));
  INV_X1    g533(.A(new_n706), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n656), .A2(new_n720), .A3(new_n637), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n434), .A2(new_n553), .A3(new_n652), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n723), .B1(new_n665), .B2(new_n669), .ZN(new_n724));
  XOR2_X1   g538(.A(KEYINPUT103), .B(G119), .Z(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G21));
  NOR2_X1   g540(.A1(new_n721), .A2(new_n673), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n295), .B1(new_n326), .B2(KEYINPUT28), .ZN(new_n728));
  OAI22_X1  g542(.A1(new_n728), .A2(new_n287), .B1(KEYINPUT31), .B2(new_n289), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n188), .B1(new_n730), .B2(new_n308), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n601), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n727), .A2(new_n391), .A3(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G122), .ZN(G24));
  OAI21_X1  g548(.A(new_n189), .B1(new_n292), .B2(new_n729), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n735), .B(new_n652), .C1(new_n604), .C2(new_n600), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n656), .A2(new_n720), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n736), .A2(new_n737), .A3(new_n697), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(new_n336), .ZN(G27));
  INV_X1    g553(.A(KEYINPUT42), .ZN(new_n740));
  INV_X1    g554(.A(new_n697), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n495), .A2(new_n496), .A3(new_n507), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n610), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n332), .A2(new_n391), .A3(new_n741), .A4(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n596), .A2(KEYINPUT42), .A3(new_n742), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n746), .A2(new_n697), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT104), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n666), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n309), .A2(KEYINPUT104), .A3(new_n313), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n188), .B1(new_n307), .B2(new_n308), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n331), .B1(KEYINPUT32), .B2(new_n752), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n747), .B(new_n391), .C1(new_n751), .C2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(KEYINPUT105), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n300), .A2(new_n302), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n756), .A2(new_n749), .A3(new_n331), .A4(new_n750), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT105), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n757), .A2(new_n758), .A3(new_n391), .A4(new_n747), .ZN(new_n759));
  AOI22_X1  g573(.A1(new_n740), .A2(new_n745), .B1(new_n755), .B2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(new_n198), .ZN(G33));
  INV_X1    g575(.A(new_n663), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n332), .A2(new_n391), .A3(new_n762), .A4(new_n744), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G134), .ZN(G36));
  AOI21_X1  g578(.A(new_n690), .B1(new_n606), .B2(new_n607), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n433), .B(KEYINPUT107), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT43), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n625), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n767), .B1(new_n433), .B2(new_n625), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(KEYINPUT44), .B1(new_n765), .B2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n583), .A2(KEYINPUT45), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT45), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n775), .B1(new_n579), .B2(new_n582), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n774), .A2(new_n776), .A3(G469), .ZN(new_n777));
  NAND2_X1  g591(.A1(G469), .A2(G902), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT46), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n777), .A2(KEYINPUT46), .A3(new_n778), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n781), .A2(new_n595), .A3(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n783), .A2(new_n554), .A3(new_n676), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT106), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n783), .A2(KEYINPUT106), .A3(new_n554), .A4(new_n676), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n786), .A2(new_n742), .A3(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n765), .A2(KEYINPUT44), .A3(new_n771), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n773), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G137), .ZN(G39));
  NAND2_X1  g606(.A1(new_n783), .A2(new_n554), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT47), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n783), .A2(KEYINPUT47), .A3(new_n554), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n665), .A2(new_n669), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n697), .A2(new_n391), .A3(new_n743), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G140), .ZN(G42));
  NAND2_X1  g615(.A1(new_n498), .A2(new_n283), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT115), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n732), .A2(new_n391), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n672), .A2(new_n506), .A3(new_n706), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n771), .A2(new_n805), .A3(new_n499), .A4(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT50), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n661), .B1(new_n769), .B2(new_n770), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n810), .A2(KEYINPUT50), .A3(new_n805), .A4(new_n806), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(new_n736), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n743), .A2(new_n706), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n810), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  NOR4_X1   g629(.A1(new_n390), .A2(new_n743), .A3(new_n706), .A4(new_n661), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n433), .A2(new_n696), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n688), .A2(new_n816), .A3(new_n312), .A4(new_n817), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n705), .A2(new_n595), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT112), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n554), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n822), .B1(new_n821), .B2(new_n820), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n795), .A2(new_n796), .A3(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n824), .A2(new_n805), .A3(new_n742), .A4(new_n810), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n812), .A2(new_n819), .A3(KEYINPUT51), .A4(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT113), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n826), .B(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n812), .A2(new_n819), .A3(new_n825), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT51), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n737), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n810), .A2(new_n832), .A3(new_n805), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n688), .A2(new_n816), .A3(new_n312), .A4(new_n632), .ZN(new_n834));
  AND4_X1   g648(.A1(G952), .A2(new_n833), .A3(new_n283), .A4(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n757), .A2(new_n391), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n810), .A2(new_n837), .A3(new_n814), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(KEYINPUT48), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT48), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n810), .A2(new_n837), .A3(new_n840), .A4(new_n814), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT114), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n835), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n843), .B1(new_n835), .B2(new_n842), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n831), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n803), .B1(new_n828), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n718), .A2(new_n724), .A3(new_n733), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n332), .A2(new_n711), .A3(new_n712), .ZN(new_n849));
  OAI21_X1  g663(.A(KEYINPUT102), .B1(new_n798), .B2(new_n708), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n745), .A2(new_n740), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n755), .A2(new_n759), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n598), .A2(new_n653), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n610), .A2(new_n390), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n606), .A2(new_n607), .A3(new_n508), .A4(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n644), .A2(KEYINPUT109), .ZN(new_n858));
  INV_X1    g672(.A(new_n632), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT109), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n860), .B1(new_n553), .B2(new_n433), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n858), .A2(new_n859), .A3(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n857), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n855), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n744), .A2(new_n652), .ZN(new_n865));
  INV_X1    g679(.A(new_n662), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n658), .A2(new_n433), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n867), .B1(new_n665), .B2(new_n669), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n732), .A2(new_n741), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n865), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AND4_X1   g684(.A1(new_n332), .A2(new_n391), .A3(new_n762), .A4(new_n744), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n851), .A2(new_n854), .A3(new_n864), .A4(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n636), .A2(new_n639), .ZN(new_n874));
  NOR4_X1   g688(.A1(new_n673), .A2(new_n610), .A3(new_n874), .A4(new_n866), .ZN(new_n875));
  OAI211_X1 g689(.A(new_n690), .B(new_n875), .C1(new_n665), .C2(new_n687), .ZN(new_n876));
  INV_X1    g690(.A(new_n738), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n876), .A2(new_n670), .A3(new_n699), .A4(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT52), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n738), .B1(new_n332), .B2(new_n664), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n881), .A2(KEYINPUT52), .A3(new_n699), .A4(new_n876), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(KEYINPUT53), .B1(new_n873), .B2(new_n883), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n851), .A2(new_n864), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT53), .ZN(new_n886));
  AOI22_X1  g700(.A1(new_n332), .A2(new_n867), .B1(new_n741), .B2(new_n732), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n763), .B1(new_n887), .B2(new_n865), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n760), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n885), .A2(new_n886), .A3(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n880), .A2(KEYINPUT110), .A3(new_n882), .ZN(new_n891));
  OR3_X1    g705(.A1(new_n878), .A2(KEYINPUT110), .A3(new_n879), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n884), .B(KEYINPUT54), .C1(new_n890), .C2(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n886), .B1(new_n873), .B2(new_n883), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT54), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT111), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n897), .B1(new_n714), .B2(new_n848), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n850), .A2(new_n849), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n718), .A2(new_n724), .A3(new_n733), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n899), .A2(KEYINPUT111), .A3(new_n900), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n855), .A2(new_n863), .A3(new_n886), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n889), .A2(new_n898), .A3(new_n901), .A4(new_n902), .ZN(new_n903));
  OAI211_X1 g717(.A(new_n895), .B(new_n896), .C1(new_n893), .C2(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n847), .A2(new_n894), .A3(new_n904), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n828), .A2(new_n846), .A3(new_n803), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n802), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n820), .A2(KEYINPUT49), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n672), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n909), .B1(KEYINPUT49), .B2(new_n820), .ZN(new_n910));
  INV_X1    g724(.A(new_n766), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n391), .A2(new_n554), .A3(new_n506), .A4(new_n696), .ZN(new_n912));
  NOR4_X1   g726(.A1(new_n910), .A2(new_n689), .A3(new_n911), .A4(new_n912), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT108), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n907), .A2(new_n914), .ZN(G75));
  NOR2_X1   g729(.A1(new_n283), .A2(G952), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT117), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(new_n895), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n903), .A2(new_n893), .ZN(new_n920));
  OAI211_X1 g734(.A(G210), .B(G902), .C1(new_n919), .C2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT56), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n469), .A2(new_n471), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT116), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n477), .B(KEYINPUT55), .Z(new_n926));
  XOR2_X1   g740(.A(new_n925), .B(new_n926), .Z(new_n927));
  NAND2_X1  g741(.A1(new_n923), .A2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(new_n927), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n921), .A2(new_n922), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n918), .B1(new_n928), .B2(new_n930), .ZN(G51));
  XOR2_X1   g745(.A(new_n778), .B(KEYINPUT57), .Z(new_n932));
  INV_X1    g746(.A(new_n904), .ZN(new_n933));
  AND4_X1   g747(.A1(new_n889), .A2(new_n898), .A3(new_n901), .A4(new_n902), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n891), .A2(new_n892), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n896), .B1(new_n936), .B2(new_n895), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n932), .B1(new_n933), .B2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(new_n704), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n936), .A2(new_n895), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n777), .B(KEYINPUT118), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n941), .A2(G902), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n916), .B1(new_n940), .B2(new_n943), .ZN(G54));
  AND2_X1   g758(.A1(KEYINPUT58), .A2(G475), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n941), .A2(G902), .A3(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n946), .A2(new_n417), .A3(new_n423), .ZN(new_n947));
  INV_X1    g761(.A(new_n916), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n941), .A2(G902), .A3(new_n424), .A4(new_n945), .ZN(new_n949));
  AND3_X1   g763(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(G60));
  NAND2_X1  g764(.A1(new_n894), .A2(new_n904), .ZN(new_n951));
  NAND2_X1  g765(.A1(G478), .A2(G902), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT59), .Z(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n622), .B1(new_n951), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n622), .A2(new_n954), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n941), .A2(KEYINPUT54), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n956), .B1(new_n957), .B2(new_n904), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n955), .A2(new_n958), .A3(new_n918), .ZN(G63));
  XNOR2_X1  g773(.A(KEYINPUT119), .B(KEYINPUT60), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n380), .A2(new_n324), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n960), .B(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n941), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n379), .B(KEYINPUT120), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n650), .B(new_n962), .C1(new_n919), .C2(new_n920), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n965), .A2(KEYINPUT61), .A3(new_n917), .A4(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n962), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n968), .B1(new_n936), .B2(new_n895), .ZN(new_n969));
  INV_X1    g783(.A(new_n964), .ZN(new_n970));
  OAI211_X1 g784(.A(new_n966), .B(new_n917), .C1(new_n969), .C2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT61), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n967), .A2(new_n973), .ZN(G66));
  OAI21_X1  g788(.A(G953), .B1(new_n475), .B2(new_n504), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n975), .B1(new_n885), .B2(G953), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n925), .B1(G898), .B2(new_n283), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n976), .B(new_n977), .ZN(G69));
  AOI21_X1  g792(.A(new_n283), .B1(G227), .B2(G900), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n273), .A2(new_n280), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(new_n419), .ZN(new_n981));
  NAND2_X1  g795(.A1(G900), .A2(G953), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n670), .A2(new_n699), .A3(new_n877), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(KEYINPUT121), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT121), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n881), .A2(new_n985), .A3(new_n699), .ZN(new_n986));
  AND2_X1   g800(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n673), .A2(new_n874), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n837), .A2(new_n786), .A3(new_n787), .A4(new_n988), .ZN(new_n989));
  AND3_X1   g803(.A1(new_n800), .A2(new_n989), .A3(new_n763), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n987), .A2(new_n990), .A3(new_n854), .A4(new_n791), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n981), .B(new_n982), .C1(new_n991), .C2(G953), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n979), .B1(new_n992), .B2(KEYINPUT125), .ZN(new_n993));
  INV_X1    g807(.A(new_n790), .ZN(new_n994));
  NOR3_X1   g808(.A1(new_n994), .A2(new_n772), .A3(new_n788), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT123), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n390), .B1(new_n709), .B2(new_n312), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(new_n744), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n858), .A2(new_n859), .A3(new_n861), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n999), .A2(new_n676), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n996), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1000), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n1002), .A2(KEYINPUT123), .A3(new_n997), .A4(new_n744), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g818(.A(KEYINPUT124), .B1(new_n995), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(KEYINPUT124), .ZN(new_n1006));
  NAND4_X1  g820(.A1(new_n791), .A2(new_n1006), .A3(new_n1001), .A4(new_n1003), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g822(.A(KEYINPUT62), .ZN(new_n1009));
  NAND4_X1  g823(.A1(new_n984), .A2(new_n986), .A3(new_n1009), .A4(new_n691), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1010), .A2(new_n800), .ZN(new_n1011));
  INV_X1    g825(.A(new_n1011), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n984), .A2(new_n691), .A3(new_n986), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1013), .A2(KEYINPUT62), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n1014), .A2(KEYINPUT122), .ZN(new_n1015));
  INV_X1    g829(.A(KEYINPUT122), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1016), .B1(new_n1013), .B2(KEYINPUT62), .ZN(new_n1017));
  OAI211_X1 g831(.A(new_n1008), .B(new_n1012), .C1(new_n1015), .C2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n981), .B1(new_n1018), .B2(new_n283), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n981), .A2(new_n982), .ZN(new_n1020));
  AND4_X1   g834(.A1(new_n854), .A2(new_n987), .A3(new_n990), .A4(new_n791), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1020), .B1(new_n1021), .B2(new_n283), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n993), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g837(.A(new_n979), .ZN(new_n1024));
  INV_X1    g838(.A(KEYINPUT125), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n1024), .B1(new_n1022), .B2(new_n1025), .ZN(new_n1026));
  OR2_X1    g840(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n1011), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1028));
  AOI21_X1  g842(.A(G953), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  OAI211_X1 g843(.A(new_n1026), .B(new_n992), .C1(new_n1029), .C2(new_n981), .ZN(new_n1030));
  AND2_X1   g844(.A1(new_n1023), .A2(new_n1030), .ZN(G72));
  NAND2_X1  g845(.A1(G472), .A2(G902), .ZN(new_n1032));
  XNOR2_X1  g846(.A(new_n1032), .B(KEYINPUT63), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n1033), .B1(new_n681), .B2(new_n320), .ZN(new_n1034));
  OAI211_X1 g848(.A(new_n884), .B(new_n1034), .C1(new_n890), .C2(new_n893), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1021), .A2(new_n885), .ZN(new_n1036));
  XNOR2_X1  g850(.A(new_n1033), .B(KEYINPUT126), .ZN(new_n1037));
  AND2_X1   g851(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g852(.A(new_n319), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1039), .A2(new_n306), .ZN(new_n1040));
  OAI211_X1 g854(.A(new_n948), .B(new_n1035), .C1(new_n1038), .C2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n851), .A2(new_n864), .ZN(new_n1042));
  OAI21_X1  g856(.A(new_n1037), .B1(new_n1018), .B2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g857(.A1(new_n1039), .A2(new_n306), .ZN(new_n1044));
  AOI21_X1  g858(.A(new_n1041), .B1(new_n1043), .B2(new_n1044), .ZN(G57));
endmodule


