//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 1 1 0 1 1 0 1 0 1 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 1 0 0 0 0 1 0 1 0 1 1 1 1 0 1 1 0 1 0 1 1 0 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:10 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1284, new_n1285,
    new_n1286, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1342, new_n1343, new_n1344;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(G13), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(KEYINPUT64), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g0016(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n219), .A2(new_n207), .ZN(new_n220));
  OAI21_X1  g0020(.A(G50), .B1(G58), .B2(G68), .ZN(new_n221));
  INV_X1    g0021(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT1), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G107), .A2(G264), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n228));
  AND4_X1   g0028(.A1(new_n225), .A2(new_n226), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT65), .B(G238), .ZN(new_n230));
  INV_X1    g0030(.A(G68), .ZN(new_n231));
  OR2_X1    g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n208), .B1(new_n229), .B2(new_n232), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n213), .B(new_n223), .C1(new_n224), .C2(new_n233), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n233), .A2(new_n224), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT66), .ZN(new_n236));
  NOR2_X1   g0036(.A1(new_n234), .A2(new_n236), .ZN(G361));
  XOR2_X1   g0037(.A(G250), .B(G257), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT67), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G238), .B(G244), .ZN(new_n242));
  INV_X1    g0042(.A(G232), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(KEYINPUT2), .B(G226), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n241), .B(new_n246), .ZN(G358));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n202), .A2(G68), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n231), .A2(G50), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(G58), .B(G77), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n250), .B(new_n255), .ZN(G351));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  AND3_X1   g0057(.A1(new_n216), .A2(new_n217), .A3(new_n257), .ZN(new_n258));
  NOR3_X1   g0058(.A1(new_n209), .A2(new_n207), .A3(G1), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n206), .A2(G20), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G50), .ZN(new_n263));
  OAI22_X1  g0063(.A1(new_n261), .A2(new_n263), .B1(G50), .B2(new_n260), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT68), .ZN(new_n265));
  XNOR2_X1  g0065(.A(new_n264), .B(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n203), .A2(G20), .ZN(new_n267));
  NOR2_X1   g0067(.A1(G20), .A2(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G150), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT8), .B(G58), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n207), .A2(G33), .ZN(new_n271));
  OAI211_X1 g0071(.A(new_n267), .B(new_n269), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n216), .A2(new_n217), .A3(new_n257), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n266), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G274), .ZN(new_n276));
  AND2_X1   g0076(.A1(G1), .A2(G13), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G33), .A2(G41), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G226), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n278), .A2(G1), .A3(G13), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n280), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n282), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT3), .ZN(new_n287));
  INV_X1    g0087(.A(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(KEYINPUT3), .A2(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G1698), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n291), .A2(G222), .A3(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n291), .A2(G223), .A3(G1698), .ZN(new_n294));
  INV_X1    g0094(.A(G77), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n293), .B(new_n294), .C1(new_n295), .C2(new_n291), .ZN(new_n296));
  AND2_X1   g0096(.A1(G33), .A2(G41), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n297), .B1(new_n216), .B2(new_n217), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n286), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G179), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n275), .B(new_n301), .C1(G169), .C2(new_n299), .ZN(new_n302));
  XNOR2_X1  g0102(.A(new_n275), .B(KEYINPUT9), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT10), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT69), .ZN(new_n305));
  INV_X1    g0105(.A(G200), .ZN(new_n306));
  OR3_X1    g0106(.A1(new_n299), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n305), .B1(new_n299), .B2(new_n306), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n307), .A2(new_n308), .B1(G190), .B2(new_n299), .ZN(new_n309));
  AND3_X1   g0109(.A1(new_n303), .A2(new_n304), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n304), .B1(new_n303), .B2(new_n309), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n302), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G169), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n218), .A2(new_n278), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n283), .A2(G1698), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n291), .B(new_n315), .C1(G223), .C2(G1698), .ZN(new_n316));
  NAND2_X1  g0116(.A1(G33), .A2(G87), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n314), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n282), .B1(new_n243), .B2(new_n285), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n313), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  NOR3_X1   g0122(.A1(new_n318), .A2(new_n300), .A3(new_n320), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT16), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n289), .A2(new_n207), .A3(new_n290), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT7), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n289), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n290), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n231), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(G58), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n331), .A2(new_n231), .ZN(new_n332));
  OAI21_X1  g0132(.A(G20), .B1(new_n332), .B2(new_n201), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n268), .A2(G159), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n325), .B1(new_n330), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(KEYINPUT75), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n328), .A2(new_n329), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n335), .B1(new_n338), .B2(G68), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n258), .B1(new_n339), .B2(KEYINPUT16), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT75), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n341), .B(new_n325), .C1(new_n330), .C2(new_n335), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n337), .A2(new_n340), .A3(new_n342), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n273), .A2(new_n259), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n270), .B1(new_n206), .B2(G20), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n344), .A2(new_n345), .B1(new_n259), .B2(new_n270), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n324), .B1(new_n343), .B2(new_n346), .ZN(new_n347));
  XNOR2_X1  g0147(.A(new_n347), .B(KEYINPUT18), .ZN(new_n348));
  INV_X1    g0148(.A(G190), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n319), .A2(new_n321), .A3(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n306), .B1(new_n318), .B2(new_n320), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n343), .A2(new_n346), .A3(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT76), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n343), .A2(KEYINPUT76), .A3(new_n346), .A4(new_n352), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n355), .A2(KEYINPUT17), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT17), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n343), .A2(new_n359), .A3(new_n346), .A4(new_n352), .ZN(new_n360));
  XNOR2_X1  g0160(.A(new_n360), .B(KEYINPUT77), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n348), .B1(new_n358), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n259), .A2(new_n231), .ZN(new_n363));
  XOR2_X1   g0163(.A(new_n363), .B(KEYINPUT12), .Z(new_n364));
  INV_X1    g0164(.A(KEYINPUT11), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n268), .A2(G50), .B1(G20), .B2(new_n231), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n366), .B1(new_n295), .B2(new_n271), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n273), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n364), .B1(new_n365), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n367), .A2(KEYINPUT11), .A3(new_n273), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n344), .A2(G68), .A3(new_n262), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  AND2_X1   g0172(.A1(new_n284), .A2(new_n280), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n373), .A2(G238), .B1(new_n281), .B2(new_n279), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n283), .A2(new_n292), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n243), .A2(G1698), .ZN(new_n376));
  AND2_X1   g0176(.A1(KEYINPUT3), .A2(G33), .ZN(new_n377));
  NOR2_X1   g0177(.A1(KEYINPUT3), .A2(G33), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n375), .B(new_n376), .C1(new_n377), .C2(new_n378), .ZN(new_n379));
  AND3_X1   g0179(.A1(KEYINPUT70), .A2(G33), .A3(G97), .ZN(new_n380));
  AOI21_X1  g0180(.A(KEYINPUT70), .B1(G33), .B2(G97), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n298), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT13), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n374), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT71), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n314), .B1(new_n382), .B2(new_n379), .ZN(new_n389));
  INV_X1    g0189(.A(G238), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n282), .B1(new_n390), .B2(new_n285), .ZN(new_n391));
  OAI21_X1  g0191(.A(KEYINPUT13), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n374), .A2(new_n384), .A3(KEYINPUT71), .A4(new_n385), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n388), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT14), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n394), .A2(new_n395), .A3(G169), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n392), .A2(G179), .A3(new_n386), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(KEYINPUT74), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT74), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n392), .A2(new_n399), .A3(G179), .A4(new_n386), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n395), .B1(new_n394), .B2(G169), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n396), .B(new_n401), .C1(new_n402), .C2(KEYINPUT73), .ZN(new_n403));
  AND2_X1   g0203(.A1(new_n392), .A2(new_n393), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n313), .B1(new_n404), .B2(new_n388), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT73), .ZN(new_n406));
  NOR3_X1   g0206(.A1(new_n405), .A2(new_n406), .A3(new_n395), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n372), .B1(new_n403), .B2(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n392), .A2(G190), .A3(new_n386), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT72), .ZN(new_n410));
  XNOR2_X1  g0210(.A(new_n409), .B(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n394), .A2(G200), .ZN(new_n412));
  INV_X1    g0212(.A(new_n372), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n408), .A2(new_n414), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n377), .A2(new_n378), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n230), .A2(G1698), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n243), .A2(new_n292), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n416), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n298), .B1(G107), .B2(new_n291), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(G244), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n282), .B1(new_n422), .B2(new_n285), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(G200), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n424), .A2(G190), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n344), .A2(G77), .A3(new_n262), .ZN(new_n428));
  INV_X1    g0228(.A(new_n270), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n429), .A2(new_n268), .B1(G20), .B2(G77), .ZN(new_n430));
  XNOR2_X1  g0230(.A(KEYINPUT15), .B(G87), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n430), .B1(new_n271), .B2(new_n431), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n432), .A2(new_n273), .B1(new_n295), .B2(new_n259), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n426), .A2(new_n427), .A3(new_n428), .A4(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n425), .A2(new_n313), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n433), .A2(new_n428), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n424), .A2(new_n300), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  NOR4_X1   g0239(.A1(new_n312), .A2(new_n362), .A3(new_n415), .A4(new_n439), .ZN(new_n440));
  AND2_X1   g0240(.A1(KEYINPUT5), .A2(G41), .ZN(new_n441));
  NOR2_X1   g0241(.A1(KEYINPUT5), .A2(G41), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n206), .A2(G45), .ZN(new_n444));
  OAI211_X1 g0244(.A(G270), .B(new_n284), .C1(new_n443), .C2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(G45), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n446), .A2(G1), .ZN(new_n447));
  XNOR2_X1  g0247(.A(KEYINPUT5), .B(G41), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n279), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  AND2_X1   g0249(.A1(new_n445), .A2(new_n449), .ZN(new_n450));
  OAI211_X1 g0250(.A(G264), .B(G1698), .C1(new_n377), .C2(new_n378), .ZN(new_n451));
  OAI211_X1 g0251(.A(G257), .B(new_n292), .C1(new_n377), .C2(new_n378), .ZN(new_n452));
  INV_X1    g0252(.A(G303), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n451), .B(new_n452), .C1(new_n453), .C2(new_n291), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(new_n298), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n450), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n456), .A2(KEYINPUT21), .A3(G169), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n445), .A2(new_n449), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n458), .B1(new_n298), .B2(new_n454), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(G179), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g0261(.A(KEYINPUT78), .B1(new_n288), .B2(G1), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT78), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n463), .A2(new_n206), .A3(G33), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n258), .A2(G116), .A3(new_n260), .A4(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(G116), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n259), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(G20), .B1(G33), .B2(G283), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n288), .A2(G97), .ZN(new_n470));
  AOI22_X1  g0270(.A1(new_n469), .A2(new_n470), .B1(G20), .B2(new_n467), .ZN(new_n471));
  AND3_X1   g0271(.A1(new_n471), .A2(new_n273), .A3(KEYINPUT20), .ZN(new_n472));
  AOI21_X1  g0272(.A(KEYINPUT20), .B1(new_n471), .B2(new_n273), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n466), .B(new_n468), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT82), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n471), .A2(new_n273), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT20), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n471), .A2(new_n273), .A3(KEYINPUT20), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n481), .A2(KEYINPUT82), .A3(new_n466), .A4(new_n468), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n476), .A2(new_n482), .ZN(new_n483));
  AND3_X1   g0283(.A1(new_n461), .A2(KEYINPUT83), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(KEYINPUT83), .B1(new_n461), .B2(new_n483), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n459), .A2(new_n313), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(KEYINPUT84), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT21), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT84), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n483), .A2(new_n491), .A3(new_n487), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n489), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n483), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n456), .A2(G200), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n494), .B(new_n495), .C1(new_n349), .C2(new_n456), .ZN(new_n496));
  AND3_X1   g0296(.A1(new_n486), .A2(new_n493), .A3(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT87), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n258), .A2(new_n260), .A3(new_n465), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(KEYINPUT86), .A2(KEYINPUT25), .ZN(new_n501));
  INV_X1    g0301(.A(G107), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n502), .B1(KEYINPUT86), .B2(KEYINPUT25), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n501), .B1(new_n260), .B2(new_n503), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n259), .A2(KEYINPUT86), .A3(KEYINPUT25), .A4(new_n502), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n500), .A2(G107), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n207), .B(G87), .C1(new_n377), .C2(new_n378), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(KEYINPUT22), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT22), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n291), .A2(new_n510), .A3(new_n207), .A4(G87), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT23), .ZN(new_n514));
  OAI22_X1  g0314(.A1(new_n513), .A2(G20), .B1(new_n514), .B2(new_n502), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n514), .A2(new_n502), .A3(G20), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(KEYINPUT85), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT85), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n518), .A2(new_n514), .A3(new_n502), .A4(G20), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n515), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n512), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(KEYINPUT24), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT24), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n512), .A2(new_n523), .A3(new_n520), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n507), .B1(new_n525), .B2(new_n273), .ZN(new_n526));
  OAI211_X1 g0326(.A(G257), .B(G1698), .C1(new_n377), .C2(new_n378), .ZN(new_n527));
  OAI211_X1 g0327(.A(G250), .B(new_n292), .C1(new_n377), .C2(new_n378), .ZN(new_n528));
  NAND2_X1  g0328(.A1(G33), .A2(G294), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n448), .A2(new_n447), .B1(new_n277), .B2(new_n278), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n530), .A2(new_n298), .B1(new_n531), .B2(G264), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n449), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n313), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n534), .B1(G179), .B2(new_n533), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n498), .B1(new_n526), .B2(new_n535), .ZN(new_n536));
  AND3_X1   g0336(.A1(new_n512), .A2(new_n523), .A3(new_n520), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n523), .B1(new_n512), .B2(new_n520), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n273), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n506), .ZN(new_n540));
  AND3_X1   g0340(.A1(new_n532), .A2(new_n300), .A3(new_n449), .ZN(new_n541));
  AOI21_X1  g0341(.A(G169), .B1(new_n532), .B2(new_n449), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n540), .A2(KEYINPUT87), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n536), .A2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(G97), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n259), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n547), .B1(new_n499), .B2(new_n546), .ZN(new_n548));
  AOI21_X1  g0348(.A(KEYINPUT7), .B1(new_n416), .B2(new_n207), .ZN(new_n549));
  INV_X1    g0349(.A(new_n329), .ZN(new_n550));
  OAI21_X1  g0350(.A(G107), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT6), .ZN(new_n552));
  AND2_X1   g0352(.A1(G97), .A2(G107), .ZN(new_n553));
  NOR2_X1   g0353(.A1(G97), .A2(G107), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n502), .A2(KEYINPUT6), .A3(G97), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n557), .A2(G20), .B1(G77), .B2(new_n268), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n551), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n548), .B1(new_n559), .B2(new_n273), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n284), .B1(new_n443), .B2(new_n444), .ZN(new_n561));
  INV_X1    g0361(.A(G257), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n449), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  OAI211_X1 g0363(.A(G244), .B(new_n292), .C1(new_n377), .C2(new_n378), .ZN(new_n564));
  NOR2_X1   g0364(.A1(KEYINPUT79), .A2(KEYINPUT4), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n565), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n291), .A2(G244), .A3(new_n292), .A4(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(G33), .A2(G283), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n291), .A2(G250), .A3(G1698), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n566), .A2(new_n568), .A3(new_n569), .A4(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n563), .B1(new_n571), .B2(new_n298), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n572), .A2(G200), .ZN(new_n573));
  AOI211_X1 g0373(.A(G190), .B(new_n563), .C1(new_n298), .C2(new_n571), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n560), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(new_n560), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n571), .A2(new_n298), .ZN(new_n577));
  INV_X1    g0377(.A(new_n563), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n313), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n572), .A2(new_n300), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n576), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n533), .A2(G200), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n532), .A2(G190), .A3(new_n449), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n539), .A2(new_n506), .A3(new_n583), .A4(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n575), .A2(new_n582), .A3(new_n585), .ZN(new_n586));
  OAI211_X1 g0386(.A(G238), .B(new_n292), .C1(new_n377), .C2(new_n378), .ZN(new_n587));
  OAI211_X1 g0387(.A(G244), .B(G1698), .C1(new_n377), .C2(new_n378), .ZN(new_n588));
  NAND2_X1  g0388(.A1(G33), .A2(G116), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n298), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n284), .A2(G274), .A3(new_n447), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n444), .B(G250), .C1(new_n297), .C2(new_n214), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n591), .A2(new_n349), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n594), .B1(new_n590), .B2(new_n298), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n596), .B1(G200), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n500), .A2(G87), .ZN(new_n599));
  INV_X1    g0399(.A(G87), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n554), .A2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT19), .ZN(new_n602));
  NAND2_X1  g0402(.A1(G33), .A2(G97), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT70), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(KEYINPUT70), .A2(G33), .A3(G97), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n602), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n601), .B1(new_n607), .B2(G20), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n207), .B(G68), .C1(new_n377), .C2(new_n378), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n602), .B1(new_n271), .B2(new_n546), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n258), .B1(new_n608), .B2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n431), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n613), .A2(new_n260), .ZN(new_n614));
  NOR3_X1   g0414(.A1(new_n612), .A2(KEYINPUT81), .A3(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT81), .ZN(new_n616));
  INV_X1    g0416(.A(new_n601), .ZN(new_n617));
  OAI21_X1  g0417(.A(KEYINPUT19), .B1(new_n380), .B2(new_n381), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n617), .B1(new_n618), .B2(new_n207), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n609), .A2(new_n610), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n273), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n614), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n616), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n598), .B(new_n599), .C1(new_n615), .C2(new_n623), .ZN(new_n624));
  AOI211_X1 g0424(.A(new_n300), .B(new_n594), .C1(new_n298), .C2(new_n590), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n313), .B1(new_n591), .B2(new_n595), .ZN(new_n626));
  OAI21_X1  g0426(.A(KEYINPUT80), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n597), .A2(G179), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT80), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n628), .B(new_n629), .C1(new_n313), .C2(new_n597), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g0431(.A(KEYINPUT81), .B1(new_n612), .B2(new_n614), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n621), .A2(new_n616), .A3(new_n622), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n632), .A2(new_n633), .B1(new_n613), .B2(new_n500), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n624), .B1(new_n631), .B2(new_n634), .ZN(new_n635));
  NOR3_X1   g0435(.A1(new_n545), .A2(new_n586), .A3(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n440), .A2(new_n497), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g0437(.A(new_n637), .B(KEYINPUT88), .ZN(G372));
  NAND2_X1  g0438(.A1(new_n343), .A2(new_n346), .ZN(new_n639));
  OR2_X1    g0439(.A1(new_n322), .A2(new_n323), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(KEYINPUT18), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT18), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n347), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n414), .A2(new_n436), .A3(new_n437), .A4(new_n435), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(new_n408), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT77), .ZN(new_n648));
  XNOR2_X1  g0448(.A(new_n360), .B(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n357), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n645), .B1(new_n647), .B2(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n310), .A2(new_n311), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n302), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT90), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  OAI211_X1 g0455(.A(KEYINPUT90), .B(new_n302), .C1(new_n651), .C2(new_n652), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n627), .A2(new_n630), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n500), .A2(new_n613), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n659), .B1(new_n615), .B2(new_n623), .ZN(new_n660));
  AOI22_X1  g0460(.A1(new_n632), .A2(new_n633), .B1(G87), .B2(new_n500), .ZN(new_n661));
  AOI22_X1  g0461(.A1(new_n658), .A2(new_n660), .B1(new_n661), .B2(new_n598), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT89), .ZN(new_n663));
  AOI211_X1 g0463(.A(G179), .B(new_n563), .C1(new_n298), .C2(new_n571), .ZN(new_n664));
  AOI21_X1  g0464(.A(G169), .B1(new_n577), .B2(new_n578), .ZN(new_n665));
  NOR3_X1   g0465(.A1(new_n664), .A2(new_n665), .A3(new_n560), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n662), .A2(new_n663), .A3(KEYINPUT26), .A4(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n625), .A2(new_n626), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n660), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n670), .A2(new_n666), .A3(new_n624), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT26), .ZN(new_n672));
  AOI21_X1  g0472(.A(KEYINPUT89), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NOR3_X1   g0473(.A1(new_n635), .A2(new_n672), .A3(new_n582), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n667), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n670), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n540), .A2(new_n543), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n461), .A2(new_n483), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n492), .A2(new_n490), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n491), .B1(new_n483), .B2(new_n487), .ZN(new_n681));
  OAI211_X1 g0481(.A(new_n678), .B(new_n679), .C1(new_n680), .C2(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n624), .B1(new_n634), .B2(new_n668), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n586), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n677), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n440), .B1(new_n676), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n657), .A2(new_n687), .ZN(G369));
  NAND2_X1  g0488(.A1(new_n493), .A2(new_n679), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n690));
  OR2_X1    g0490(.A1(new_n690), .A2(KEYINPUT27), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(KEYINPUT27), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n691), .A2(G213), .A3(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(G343), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n494), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n689), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n486), .A2(new_n493), .A3(new_n496), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n697), .B1(new_n698), .B2(new_n696), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n699), .A2(G330), .ZN(new_n700));
  AND3_X1   g0500(.A1(new_n540), .A2(KEYINPUT87), .A3(new_n543), .ZN(new_n701));
  AOI21_X1  g0501(.A(KEYINPUT87), .B1(new_n540), .B2(new_n543), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n703), .A2(new_n585), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n526), .B2(new_n695), .ZN(new_n705));
  INV_X1    g0505(.A(new_n695), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n540), .A2(new_n543), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n700), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n540), .A2(new_n543), .A3(new_n695), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n706), .B1(new_n486), .B2(new_n493), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n704), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n709), .A2(new_n710), .A3(new_n712), .ZN(G399));
  NOR2_X1   g0513(.A1(new_n210), .A2(G41), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n601), .A2(G116), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n715), .A2(G1), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n717), .B1(new_n221), .B2(new_n715), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n718), .B(KEYINPUT28), .ZN(new_n719));
  OAI21_X1  g0519(.A(KEYINPUT26), .B1(new_n683), .B2(new_n582), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n660), .A2(new_n627), .A3(new_n630), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n721), .A2(new_n672), .A3(new_n666), .A4(new_n624), .ZN(new_n722));
  AND3_X1   g0522(.A1(new_n720), .A2(new_n670), .A3(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT83), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n679), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n461), .A2(KEYINPUT83), .A3(new_n483), .ZN(new_n726));
  OAI211_X1 g0526(.A(new_n725), .B(new_n726), .C1(new_n680), .C2(new_n681), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n684), .B1(new_n727), .B2(new_n545), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n723), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(KEYINPUT91), .B1(new_n729), .B2(new_n695), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT91), .ZN(new_n731));
  AOI211_X1 g0531(.A(new_n731), .B(new_n706), .C1(new_n723), .C2(new_n728), .ZN(new_n732));
  OAI21_X1  g0532(.A(KEYINPUT29), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n706), .B1(new_n675), .B2(new_n685), .ZN(new_n734));
  OR2_X1    g0534(.A1(new_n734), .A2(KEYINPUT29), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(G179), .B1(new_n450), .B2(new_n455), .ZN(new_n737));
  INV_X1    g0537(.A(new_n597), .ZN(new_n738));
  AND4_X1   g0538(.A1(new_n579), .A2(new_n737), .A3(new_n533), .A4(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n572), .A2(new_n625), .A3(new_n459), .A4(new_n532), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(KEYINPUT30), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT30), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n532), .A2(new_n455), .A3(new_n450), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(new_n628), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n743), .B1(new_n745), .B2(new_n572), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n740), .B1(new_n742), .B2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT31), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n695), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n747), .A2(new_n706), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(new_n748), .ZN(new_n752));
  INV_X1    g0552(.A(new_n586), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n703), .A2(new_n753), .A3(new_n662), .A4(new_n695), .ZN(new_n754));
  OAI211_X1 g0554(.A(new_n750), .B(new_n752), .C1(new_n754), .C2(new_n698), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G330), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n736), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n719), .B1(new_n758), .B2(G1), .ZN(G364));
  NOR2_X1   g0559(.A1(new_n699), .A2(G330), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n760), .B(KEYINPUT92), .ZN(new_n761));
  INV_X1    g0561(.A(new_n700), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n207), .A2(G13), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n763), .B(KEYINPUT93), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n446), .ZN(new_n765));
  NOR3_X1   g0565(.A1(new_n765), .A2(new_n206), .A3(new_n714), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n761), .A2(new_n762), .A3(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n219), .B1(G20), .B2(new_n313), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n207), .A2(G179), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n771), .A2(G190), .A3(G200), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n600), .ZN(new_n773));
  NOR2_X1   g0573(.A1(G190), .A2(G200), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n771), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(G159), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(KEYINPUT32), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n207), .A2(new_n300), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G200), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(G190), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n773), .B(new_n778), .C1(G68), .C2(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n779), .A2(new_n774), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n291), .B1(new_n783), .B2(new_n295), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n779), .A2(G190), .A3(new_n306), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n784), .B1(G58), .B2(new_n786), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n771), .A2(new_n349), .A3(G200), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n777), .A2(KEYINPUT32), .B1(G107), .B2(new_n789), .ZN(new_n790));
  NOR3_X1   g0590(.A1(new_n349), .A2(G179), .A3(G200), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n207), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n780), .A2(new_n349), .ZN(new_n794));
  AOI22_X1  g0594(.A1(G97), .A2(new_n793), .B1(new_n794), .B2(G50), .ZN(new_n795));
  NAND4_X1  g0595(.A1(new_n782), .A2(new_n787), .A3(new_n790), .A4(new_n795), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n786), .A2(G322), .B1(new_n776), .B2(G329), .ZN(new_n797));
  INV_X1    g0597(.A(new_n783), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n291), .B1(new_n798), .B2(G311), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n794), .A2(G326), .ZN(new_n801));
  XNOR2_X1  g0601(.A(KEYINPUT33), .B(G317), .ZN(new_n802));
  INV_X1    g0602(.A(new_n772), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n781), .A2(new_n802), .B1(new_n803), .B2(G303), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n793), .A2(G294), .B1(new_n789), .B2(G283), .ZN(new_n805));
  NAND4_X1  g0605(.A1(new_n800), .A2(new_n801), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n770), .B1(new_n796), .B2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(G13), .A2(G33), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(G20), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n769), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n255), .A2(new_n446), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n210), .A2(new_n291), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n815), .B1(new_n446), .B2(new_n222), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n813), .B1(new_n816), .B2(KEYINPUT94), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(KEYINPUT94), .B2(new_n816), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n210), .A2(new_n416), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n819), .A2(G355), .B1(new_n467), .B2(new_n210), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n812), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  NOR3_X1   g0621(.A1(new_n807), .A2(new_n821), .A3(new_n767), .ZN(new_n822));
  INV_X1    g0622(.A(new_n810), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n822), .B1(new_n699), .B2(new_n823), .ZN(new_n824));
  AND2_X1   g0624(.A1(new_n768), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(G396));
  NAND2_X1  g0626(.A1(new_n436), .A2(new_n706), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n434), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n438), .ZN(new_n829));
  OR2_X1    g0629(.A1(new_n438), .A2(new_n706), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n734), .B(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n766), .B1(new_n833), .B2(new_n756), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(new_n756), .B2(new_n833), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n769), .A2(new_n808), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n767), .B1(new_n295), .B2(new_n836), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n786), .A2(G143), .B1(new_n798), .B2(G159), .ZN(new_n838));
  INV_X1    g0638(.A(new_n781), .ZN(new_n839));
  INV_X1    g0639(.A(G150), .ZN(new_n840));
  INV_X1    g0640(.A(G137), .ZN(new_n841));
  INV_X1    g0641(.A(new_n794), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n838), .B1(new_n839), .B2(new_n840), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n843), .B(KEYINPUT34), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n202), .A2(new_n772), .B1(new_n788), .B2(new_n231), .ZN(new_n845));
  AND2_X1   g0645(.A1(new_n845), .A2(KEYINPUT96), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n845), .A2(KEYINPUT96), .ZN(new_n847));
  INV_X1    g0647(.A(G132), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n291), .B1(new_n775), .B2(new_n848), .C1(new_n792), .C2(new_n331), .ZN(new_n849));
  NOR3_X1   g0649(.A1(new_n846), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n416), .B1(new_n772), .B2(new_n502), .ZN(new_n851));
  XOR2_X1   g0651(.A(new_n851), .B(KEYINPUT95), .Z(new_n852));
  AOI22_X1  g0652(.A1(G116), .A2(new_n798), .B1(new_n776), .B2(G311), .ZN(new_n853));
  INV_X1    g0653(.A(G294), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n853), .B1(new_n854), .B2(new_n785), .ZN(new_n855));
  INV_X1    g0655(.A(G283), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n839), .A2(new_n856), .B1(new_n546), .B2(new_n792), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n842), .A2(new_n453), .B1(new_n788), .B2(new_n600), .ZN(new_n858));
  NOR3_X1   g0658(.A1(new_n855), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n844), .A2(new_n850), .B1(new_n852), .B2(new_n859), .ZN(new_n860));
  OAI221_X1 g0660(.A(new_n837), .B1(new_n770), .B2(new_n860), .C1(new_n832), .C2(new_n809), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n835), .A2(new_n861), .ZN(G384));
  OR2_X1    g0662(.A1(new_n557), .A2(KEYINPUT35), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n557), .A2(KEYINPUT35), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n863), .A2(G116), .A3(new_n220), .A4(new_n864), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n865), .B(KEYINPUT36), .ZN(new_n866));
  OAI21_X1  g0666(.A(G77), .B1(new_n331), .B2(new_n231), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n251), .B1(new_n867), .B2(new_n221), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n868), .A2(G1), .A3(new_n209), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n340), .A2(new_n336), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(new_n346), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(new_n640), .B2(new_n694), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n355), .A2(new_n356), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(KEYINPUT37), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT97), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n641), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n347), .A2(KEYINPUT97), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n693), .B1(new_n343), .B2(new_n346), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n878), .A2(KEYINPUT37), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n876), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n355), .A2(new_n356), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n874), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n645), .B1(new_n357), .B2(new_n649), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n871), .A2(new_n694), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n882), .B(KEYINPUT38), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(KEYINPUT100), .B1(new_n358), .B2(new_n361), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT100), .ZN(new_n887));
  AND2_X1   g0687(.A1(new_n360), .A2(new_n648), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n360), .A2(new_n648), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n357), .B(new_n887), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n886), .A2(new_n348), .A3(new_n890), .ZN(new_n891));
  AND3_X1   g0691(.A1(new_n876), .A2(new_n877), .A3(new_n879), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n355), .A2(new_n356), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n641), .A2(new_n353), .ZN(new_n894));
  OAI21_X1  g0694(.A(KEYINPUT37), .B1(new_n894), .B2(new_n878), .ZN(new_n895));
  AOI22_X1  g0695(.A1(new_n892), .A2(new_n893), .B1(new_n895), .B2(KEYINPUT99), .ZN(new_n896));
  OR2_X1    g0696(.A1(new_n895), .A2(KEYINPUT99), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n891), .A2(new_n878), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  XOR2_X1   g0698(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n899));
  OAI21_X1  g0699(.A(new_n885), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT40), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n372), .A2(new_n706), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n408), .A2(new_n414), .A3(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n406), .B1(new_n405), .B2(new_n395), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n402), .A2(KEYINPUT73), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n904), .A2(new_n905), .A3(new_n396), .A4(new_n401), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n372), .B(new_n706), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n903), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n747), .A2(KEYINPUT101), .A3(new_n749), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT101), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n741), .A2(KEYINPUT30), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n745), .A2(new_n743), .A3(new_n572), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n739), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n749), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n911), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n910), .A2(new_n916), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n917), .B(new_n752), .C1(new_n754), .C2(new_n698), .ZN(new_n918));
  AND3_X1   g0718(.A1(new_n909), .A2(new_n918), .A3(new_n832), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT102), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n901), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n909), .A2(new_n918), .A3(new_n832), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(KEYINPUT102), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n900), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT38), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n884), .B1(new_n650), .B2(new_n348), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n892), .A2(new_n893), .B1(KEYINPUT37), .B2(new_n873), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n922), .B1(new_n928), .B2(new_n885), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n924), .B1(KEYINPUT40), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n440), .A2(new_n918), .ZN(new_n931));
  OAI21_X1  g0731(.A(G330), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(new_n930), .B2(new_n931), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n645), .A2(new_n693), .ZN(new_n934));
  INV_X1    g0734(.A(new_n884), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n362), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT38), .B1(new_n936), .B2(new_n882), .ZN(new_n937));
  INV_X1    g0737(.A(new_n885), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AOI211_X1 g0739(.A(new_n706), .B(new_n831), .C1(new_n675), .C2(new_n685), .ZN(new_n940));
  INV_X1    g0740(.A(new_n830), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n909), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n934), .B1(new_n939), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n906), .A2(new_n372), .A3(new_n695), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n893), .A2(new_n877), .A3(new_n876), .A4(new_n879), .ZN(new_n946));
  AOI22_X1  g0746(.A1(new_n362), .A2(new_n935), .B1(new_n946), .B2(new_n874), .ZN(new_n947));
  AOI21_X1  g0747(.A(KEYINPUT39), .B1(new_n947), .B2(KEYINPUT38), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n898), .B2(new_n899), .ZN(new_n949));
  OAI21_X1  g0749(.A(KEYINPUT39), .B1(new_n937), .B2(new_n938), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n943), .B1(new_n945), .B2(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n733), .A2(new_n440), .A3(new_n735), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n657), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n952), .B(new_n954), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n933), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n764), .A2(G1), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n933), .B2(new_n955), .ZN(new_n958));
  OAI211_X1 g0758(.A(new_n866), .B(new_n869), .C1(new_n956), .C2(new_n958), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n959), .B(KEYINPUT103), .Z(G367));
  AND2_X1   g0760(.A1(new_n241), .A2(new_n814), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n811), .B1(new_n211), .B2(new_n431), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n839), .A2(new_n854), .B1(new_n788), .B2(new_n546), .ZN(new_n963));
  INV_X1    g0763(.A(G311), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n842), .A2(new_n964), .B1(new_n502), .B2(new_n792), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n416), .B1(new_n783), .B2(new_n856), .ZN(new_n967));
  INV_X1    g0767(.A(G317), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n785), .A2(new_n453), .B1(new_n775), .B2(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n772), .A2(new_n467), .ZN(new_n970));
  AOI211_X1 g0770(.A(new_n967), .B(new_n969), .C1(KEYINPUT46), .C2(new_n970), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n966), .B(new_n971), .C1(KEYINPUT46), .C2(new_n970), .ZN(new_n972));
  OAI22_X1  g0772(.A1(new_n772), .A2(new_n331), .B1(new_n775), .B2(new_n841), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT107), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n291), .B1(new_n785), .B2(new_n840), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n975), .B1(G50), .B2(new_n798), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n792), .A2(new_n231), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(G143), .B2(new_n794), .ZN(new_n978));
  AOI22_X1  g0778(.A1(new_n781), .A2(G159), .B1(new_n789), .B2(G77), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n976), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n972), .B1(new_n974), .B2(new_n980), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n981), .B(KEYINPUT47), .Z(new_n982));
  OAI221_X1 g0782(.A(new_n766), .B1(new_n961), .B2(new_n962), .C1(new_n982), .C2(new_n770), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n983), .B(KEYINPUT108), .Z(new_n984));
  NOR2_X1   g0784(.A1(new_n661), .A2(new_n695), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n677), .A2(new_n985), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n986), .B(KEYINPUT104), .C1(new_n683), .C2(new_n985), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(KEYINPUT104), .B2(new_n986), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n984), .B1(new_n823), .B2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n989), .A2(KEYINPUT43), .ZN(new_n992));
  INV_X1    g0792(.A(new_n709), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n575), .B(new_n582), .C1(new_n560), .C2(new_n695), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n666), .A2(new_n706), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n993), .A2(KEYINPUT106), .A3(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT105), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT106), .ZN(new_n999));
  INV_X1    g0799(.A(new_n996), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n999), .B1(new_n709), .B2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n997), .A2(new_n998), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n998), .B1(new_n997), .B2(new_n1001), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n992), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1004), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n992), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1006), .A2(new_n1007), .A3(new_n1002), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n704), .A2(new_n711), .A3(new_n996), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n1009), .A2(KEYINPUT42), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n582), .B1(new_n703), .B2(new_n994), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n1009), .A2(KEYINPUT42), .B1(new_n695), .B2(new_n1011), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n1010), .A2(new_n1012), .B1(KEYINPUT43), .B2(new_n989), .ZN(new_n1013));
  AND3_X1   g0813(.A1(new_n1005), .A2(new_n1008), .A3(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1013), .B1(new_n1005), .B2(new_n1008), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n765), .A2(new_n206), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n712), .A2(new_n710), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(new_n1000), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT44), .Z(new_n1020));
  NOR2_X1   g0820(.A1(new_n1018), .A2(new_n1000), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT45), .ZN(new_n1022));
  AND3_X1   g0822(.A1(new_n1020), .A2(new_n709), .A3(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n709), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n712), .B1(new_n708), .B2(new_n711), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(new_n700), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n757), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n714), .B(KEYINPUT41), .Z(new_n1029));
  OAI21_X1  g0829(.A(new_n1017), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n991), .B1(new_n1016), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(G387));
  INV_X1    g0832(.A(new_n1017), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1027), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(KEYINPUT109), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT109), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1027), .A2(new_n1036), .A3(new_n1033), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n705), .A2(new_n707), .A3(new_n810), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n819), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n1039), .A2(new_n716), .B1(G107), .B2(new_n211), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n246), .A2(G45), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n1041), .B(KEYINPUT110), .Z(new_n1042));
  INV_X1    g0842(.A(new_n716), .ZN(new_n1043));
  AOI211_X1 g0843(.A(G45), .B(new_n1043), .C1(G68), .C2(G77), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n270), .A2(G50), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT50), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n815), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1040), .B1(new_n1042), .B2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n766), .B1(new_n1048), .B2(new_n812), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n786), .A2(G317), .B1(new_n798), .B2(G303), .ZN(new_n1050));
  XOR2_X1   g0850(.A(KEYINPUT112), .B(G322), .Z(new_n1051));
  OAI221_X1 g0851(.A(new_n1050), .B1(new_n839), .B2(new_n964), .C1(new_n842), .C2(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT48), .ZN(new_n1053));
  OR2_X1    g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n793), .A2(G283), .B1(new_n803), .B2(G294), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT49), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n788), .A2(new_n467), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n291), .B(new_n1061), .C1(G326), .C2(new_n776), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1059), .A2(new_n1060), .A3(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n416), .B1(new_n776), .B2(G150), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n1064), .B1(new_n295), .B2(new_n772), .C1(new_n546), .C2(new_n788), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT111), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n792), .A2(new_n431), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(G159), .B2(new_n794), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n786), .A2(G50), .B1(new_n798), .B2(G68), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1068), .B(new_n1069), .C1(new_n270), .C2(new_n839), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1063), .B1(new_n1066), .B2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1049), .B1(new_n1071), .B2(new_n769), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n1035), .A2(new_n1037), .B1(new_n1038), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n758), .A2(new_n1027), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n714), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n758), .A2(new_n1027), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1073), .B1(new_n1075), .B2(new_n1076), .ZN(G393));
  INV_X1    g0877(.A(new_n1074), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n715), .B1(new_n1025), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n993), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT113), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1020), .A2(new_n709), .A3(new_n1022), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1023), .B1(new_n1024), .B2(KEYINPUT113), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1079), .B1(new_n1086), .B2(new_n1078), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1000), .A2(new_n810), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n811), .B1(new_n546), .B2(new_n211), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n250), .A2(new_n815), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n766), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(G317), .A2(new_n794), .B1(new_n786), .B2(G311), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT52), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n416), .B1(new_n783), .B2(new_n854), .C1(new_n775), .C2(new_n1051), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n839), .A2(new_n453), .B1(new_n788), .B2(new_n502), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n792), .A2(new_n467), .B1(new_n772), .B2(new_n856), .ZN(new_n1096));
  OR4_X1    g0896(.A1(new_n1093), .A2(new_n1094), .A3(new_n1095), .A4(new_n1096), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(G150), .A2(new_n794), .B1(new_n786), .B2(G159), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT114), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT51), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n416), .B1(new_n776), .B2(G143), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n1101), .B1(new_n231), .B2(new_n772), .C1(new_n600), .C2(new_n788), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT115), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n783), .A2(new_n270), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n792), .A2(new_n295), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n1104), .B(new_n1105), .C1(G50), .C2(new_n781), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1097), .B1(new_n1100), .B2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1091), .B1(new_n1108), .B2(new_n769), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n1086), .A2(new_n1033), .B1(new_n1088), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1087), .A2(new_n1110), .ZN(G390));
  NOR2_X1   g0911(.A1(new_n951), .A2(new_n809), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(KEYINPUT54), .B(G143), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n793), .A2(G159), .B1(new_n798), .B2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(new_n841), .B2(new_n839), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n803), .A2(G150), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(new_n1118), .B(KEYINPUT53), .ZN(new_n1119));
  INV_X1    g0919(.A(G125), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n291), .B1(new_n775), .B2(new_n1120), .C1(new_n785), .C2(new_n848), .ZN(new_n1121));
  INV_X1    g0921(.A(G128), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n842), .A2(new_n1122), .B1(new_n788), .B2(new_n202), .ZN(new_n1123));
  OR4_X1    g0923(.A1(new_n1117), .A2(new_n1119), .A3(new_n1121), .A4(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1105), .B1(G116), .B2(new_n786), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT118), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n502), .A2(new_n839), .B1(new_n842), .B2(new_n856), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n788), .A2(new_n231), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n416), .B1(new_n775), .B2(new_n854), .C1(new_n546), .C2(new_n783), .ZN(new_n1130));
  OR4_X1    g0930(.A1(new_n773), .A2(new_n1128), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n1125), .A2(KEYINPUT117), .B1(new_n1127), .B2(new_n1131), .ZN(new_n1132));
  AND2_X1   g0932(.A1(new_n1125), .A2(KEYINPUT117), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n769), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n836), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1134), .B(new_n766), .C1(new_n429), .C2(new_n1135), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1112), .A2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n720), .A2(new_n670), .A3(new_n722), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n703), .A2(new_n493), .A3(new_n486), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1138), .B1(new_n684), .B2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n731), .B1(new_n1140), .B2(new_n706), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n729), .A2(KEYINPUT91), .A3(new_n695), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1141), .A2(new_n1142), .A3(new_n830), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1143), .A2(new_n829), .A3(new_n909), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1144), .A2(new_n944), .A3(new_n900), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n941), .B1(new_n734), .B2(new_n832), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n909), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n944), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n949), .A2(new_n1148), .A3(new_n950), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n909), .A2(new_n755), .A3(G330), .A4(new_n832), .ZN(new_n1150));
  AND3_X1   g0950(.A1(new_n1145), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n497), .A2(new_n636), .A3(new_n695), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n910), .A2(new_n916), .B1(new_n751), .B2(new_n748), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n831), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1154), .A2(G330), .A3(new_n909), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(new_n1145), .B2(new_n1149), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1151), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1137), .B1(new_n1157), .B2(new_n1033), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n909), .B1(new_n1154), .B2(G330), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1150), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1143), .A2(new_n829), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1147), .B1(new_n756), .B2(new_n831), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(new_n1155), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1146), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n1161), .A2(new_n1162), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n440), .A2(G330), .A3(new_n918), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n953), .A2(new_n657), .A3(new_n1167), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n714), .B1(new_n1157), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1145), .A2(new_n1149), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1155), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1145), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1173), .A2(new_n1174), .A3(new_n1169), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1158), .B1(new_n1170), .B2(new_n1176), .ZN(G378));
  NAND2_X1  g0977(.A1(new_n275), .A2(new_n694), .ZN(new_n1178));
  XOR2_X1   g0978(.A(new_n1178), .B(KEYINPUT121), .Z(new_n1179));
  NAND2_X1  g0979(.A1(new_n312), .A2(new_n1179), .ZN(new_n1180));
  XOR2_X1   g0980(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1181));
  INV_X1    g0981(.A(new_n1179), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1182), .B(new_n302), .C1(new_n311), .C2(new_n310), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1180), .A2(new_n1181), .A3(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1181), .B1(new_n1180), .B2(new_n1183), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1154), .A2(new_n920), .A3(new_n909), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n923), .A2(new_n1188), .A3(KEYINPUT40), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n890), .A2(new_n348), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n887), .B1(new_n649), .B2(new_n357), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n878), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n896), .A2(new_n897), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n899), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n938), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1189), .A2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(G330), .B1(new_n929), .B2(KEYINPUT40), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1187), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(G330), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n919), .B1(new_n937), .B2(new_n938), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1200), .B1(new_n1201), .B2(new_n901), .ZN(new_n1202));
  OR2_X1    g1002(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1202), .A2(new_n924), .A3(new_n1203), .ZN(new_n1204));
  AND3_X1   g1004(.A1(new_n1199), .A2(new_n952), .A3(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n952), .B1(new_n1199), .B2(new_n1204), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1203), .A2(new_n808), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n766), .B1(new_n1135), .B2(G50), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n977), .B1(G116), .B2(new_n794), .ZN(new_n1210));
  XOR2_X1   g1010(.A(new_n1210), .B(KEYINPUT119), .Z(new_n1211));
  OR2_X1    g1011(.A1(new_n291), .A2(G41), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(new_n786), .B2(G107), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n613), .A2(new_n798), .B1(new_n776), .B2(G283), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n839), .A2(new_n546), .B1(new_n772), .B2(new_n295), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(G58), .B2(new_n789), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1211), .A2(new_n1213), .A3(new_n1214), .A4(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT58), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1212), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1220));
  AND2_X1   g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n1120), .A2(new_n842), .B1(new_n839), .B2(new_n848), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n786), .A2(G128), .B1(new_n798), .B2(G137), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1223), .B1(new_n772), .B2(new_n1113), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n1222), .B(new_n1224), .C1(G150), .C2(new_n793), .ZN(new_n1225));
  XOR2_X1   g1025(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n1226));
  NOR2_X1   g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n789), .A2(G159), .ZN(new_n1229));
  AOI211_X1 g1029(.A(G33), .B(G41), .C1(new_n776), .C2(G124), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1228), .A2(new_n1229), .A3(new_n1230), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1221), .B1(new_n1218), .B2(new_n1217), .C1(new_n1227), .C2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1209), .B1(new_n1232), .B2(new_n769), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n1207), .A2(new_n1033), .B1(new_n1208), .B2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1168), .B1(new_n1157), .B2(new_n1169), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n943), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n951), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1236), .B1(new_n1237), .B2(new_n944), .ZN(new_n1238));
  NOR3_X1   g1038(.A1(new_n1197), .A2(new_n1198), .A3(new_n1187), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1203), .B1(new_n1202), .B2(new_n924), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1238), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1199), .A2(new_n952), .A3(new_n1204), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1241), .A2(KEYINPUT57), .A3(new_n1242), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n714), .B1(new_n1235), .B2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1168), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1175), .A2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(KEYINPUT57), .B1(new_n1207), .B2(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1234), .B1(new_n1244), .B2(new_n1247), .ZN(G375));
  NAND2_X1  g1048(.A1(new_n1147), .A2(new_n808), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n766), .B1(new_n1135), .B2(G68), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n794), .A2(G294), .B1(new_n798), .B2(G107), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1251), .B1(new_n467), .B2(new_n839), .ZN(new_n1252));
  XNOR2_X1  g1052(.A(new_n1252), .B(KEYINPUT122), .ZN(new_n1253));
  OAI221_X1 g1053(.A(new_n416), .B1(new_n775), .B2(new_n453), .C1(new_n785), .C2(new_n856), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1067), .B1(G77), .B2(new_n789), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1255), .B1(new_n546), .B2(new_n772), .ZN(new_n1256));
  OR3_X1    g1056(.A1(new_n1253), .A2(new_n1254), .A3(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT123), .ZN(new_n1258));
  OR2_X1    g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  OAI22_X1  g1059(.A1(new_n842), .A2(new_n848), .B1(new_n202), .B2(new_n792), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(G159), .B2(new_n803), .ZN(new_n1261));
  OAI22_X1  g1061(.A1(new_n783), .A2(new_n840), .B1(new_n775), .B2(new_n1122), .ZN(new_n1262));
  AOI211_X1 g1062(.A(new_n416), .B(new_n1262), .C1(G137), .C2(new_n786), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n781), .A2(new_n1114), .B1(new_n789), .B2(G58), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1261), .A2(new_n1263), .A3(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1259), .A2(new_n1265), .A3(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1250), .B1(new_n1267), .B2(new_n769), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1249), .A2(new_n1268), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1269), .B1(new_n1166), .B2(new_n1017), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1169), .A2(new_n1029), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1270), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(G381));
  XNOR2_X1  g1074(.A(G375), .B(KEYINPUT124), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1276));
  OAI22_X1  g1076(.A1(new_n1276), .A2(new_n1017), .B1(new_n1112), .B2(new_n1136), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1169), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n715), .B1(new_n1276), .B2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1277), .B1(new_n1175), .B2(new_n1279), .ZN(new_n1280));
  OAI211_X1 g1080(.A(new_n1073), .B(new_n825), .C1(new_n1076), .C2(new_n1075), .ZN(new_n1281));
  NOR4_X1   g1081(.A1(G390), .A2(G384), .A3(G381), .A4(new_n1281), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1275), .A2(new_n1031), .A3(new_n1280), .A4(new_n1282), .ZN(G407));
  INV_X1    g1083(.A(G213), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1284), .A2(G343), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1275), .A2(new_n1280), .A3(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(G407), .A2(new_n1286), .A3(G213), .ZN(G409));
  INV_X1    g1087(.A(KEYINPUT61), .ZN(new_n1288));
  OAI211_X1 g1088(.A(G378), .B(new_n1234), .C1(new_n1244), .C2(new_n1247), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1290));
  NOR3_X1   g1090(.A1(new_n1235), .A2(new_n1290), .A3(new_n1029), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1208), .A2(new_n1233), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1292), .B1(new_n1290), .B2(new_n1017), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1280), .B1(new_n1291), .B2(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1285), .B1(new_n1289), .B2(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1166), .A2(new_n1168), .A3(KEYINPUT60), .ZN(new_n1296));
  AND2_X1   g1096(.A1(new_n1296), .A2(new_n714), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT60), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1272), .B1(new_n1169), .B2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1297), .A2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1270), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(G384), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1300), .A2(G384), .A3(new_n1301), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1285), .A2(G2897), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1306), .A2(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(G384), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1310));
  AOI211_X1 g1110(.A(new_n1303), .B(new_n1270), .C1(new_n1297), .C2(new_n1299), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(new_n1307), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1309), .A2(new_n1313), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1288), .B1(new_n1295), .B2(new_n1314), .ZN(new_n1315));
  AND2_X1   g1115(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1316));
  AOI211_X1 g1116(.A(new_n1285), .B(new_n1306), .C1(new_n1289), .C2(new_n1294), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1316), .B1(new_n1317), .B2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1295), .A2(new_n1312), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1321), .A2(new_n1318), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1315), .B1(new_n1320), .B2(new_n1322), .ZN(new_n1323));
  OR2_X1    g1123(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n825), .B1(new_n1324), .B2(new_n1073), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1281), .ZN(new_n1326));
  OAI211_X1 g1126(.A(new_n1087), .B(new_n1110), .C1(new_n1325), .C2(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(G393), .A2(G396), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(G390), .A2(new_n1281), .A3(new_n1328), .ZN(new_n1329));
  AND3_X1   g1129(.A1(new_n1327), .A2(new_n1329), .A3(new_n1031), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1031), .B1(new_n1327), .B2(new_n1329), .ZN(new_n1331));
  NOR2_X1   g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  XNOR2_X1  g1132(.A(new_n1317), .B(KEYINPUT63), .ZN(new_n1333));
  XNOR2_X1  g1133(.A(new_n1312), .B(new_n1308), .ZN(new_n1334));
  AND2_X1   g1134(.A1(new_n1289), .A2(new_n1294), .ZN(new_n1335));
  OAI211_X1 g1135(.A(new_n1334), .B(KEYINPUT125), .C1(new_n1335), .C2(new_n1285), .ZN(new_n1336));
  NOR3_X1   g1136(.A1(new_n1330), .A2(new_n1331), .A3(KEYINPUT61), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT125), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1338), .B1(new_n1295), .B2(new_n1314), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1336), .A2(new_n1337), .A3(new_n1339), .ZN(new_n1340));
  OAI22_X1  g1140(.A1(new_n1323), .A2(new_n1332), .B1(new_n1333), .B2(new_n1340), .ZN(G405));
  NAND2_X1  g1141(.A1(G375), .A2(new_n1280), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1342), .A2(new_n1289), .ZN(new_n1343));
  XNOR2_X1  g1143(.A(new_n1343), .B(new_n1306), .ZN(new_n1344));
  XNOR2_X1  g1144(.A(new_n1344), .B(new_n1332), .ZN(G402));
endmodule


