//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 0 1 1 0 0 1 1 1 0 1 0 0 0 0 1 0 0 0 1 1 1 0 0 1 0 0 0 1 0 0 1 0 1 1 0 1 1 0 0 0 1 0 1 0 0 1 0 0 0 1 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:45 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n599, new_n600, new_n601, new_n602, new_n603,
    new_n604, new_n605, new_n606, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n653, new_n654, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935;
  XNOR2_X1  g000(.A(G143), .B(G146), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT0), .B(G128), .ZN(new_n188));
  OR2_X1    g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n187), .A2(KEYINPUT0), .A3(G128), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(KEYINPUT67), .A3(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  AOI21_X1  g006(.A(KEYINPUT67), .B1(new_n189), .B2(new_n190), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G131), .ZN(new_n195));
  INV_X1    g009(.A(G134), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT64), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G134), .ZN(new_n199));
  INV_X1    g013(.A(G137), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n197), .A2(new_n199), .A3(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT11), .ZN(new_n202));
  AND3_X1   g016(.A1(new_n201), .A2(KEYINPUT65), .A3(new_n202), .ZN(new_n203));
  AOI21_X1  g017(.A(KEYINPUT65), .B1(new_n201), .B2(new_n202), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NOR3_X1   g019(.A1(new_n202), .A2(new_n196), .A3(G137), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n197), .A2(new_n199), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n206), .B1(new_n207), .B2(G137), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n195), .B1(new_n205), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n201), .A2(new_n202), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT65), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n201), .A2(KEYINPUT65), .A3(new_n202), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n212), .A2(new_n195), .A3(new_n208), .A4(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n194), .B1(new_n209), .B2(new_n215), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n201), .B1(G134), .B2(new_n200), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G131), .ZN(new_n218));
  OR2_X1    g032(.A1(new_n187), .A2(G128), .ZN(new_n219));
  INV_X1    g033(.A(G143), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(KEYINPUT1), .A3(G146), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT1), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n187), .A2(new_n222), .A3(G128), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n219), .A2(new_n221), .A3(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n214), .A2(new_n218), .A3(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n216), .A2(KEYINPUT30), .A3(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT30), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n189), .A2(new_n190), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n212), .A2(new_n208), .A3(new_n213), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G131), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n228), .B1(new_n230), .B2(new_n214), .ZN(new_n231));
  INV_X1    g045(.A(new_n225), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n227), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  XOR2_X1   g047(.A(KEYINPUT2), .B(G113), .Z(new_n234));
  XNOR2_X1  g048(.A(G116), .B(G119), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g050(.A(new_n236), .B(KEYINPUT66), .ZN(new_n237));
  OR2_X1    g051(.A1(new_n234), .A2(new_n235), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n226), .A2(new_n233), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n239), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n216), .A2(new_n241), .A3(new_n225), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT68), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G953), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(KEYINPUT69), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT69), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G953), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G237), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n249), .A2(G210), .A3(new_n250), .ZN(new_n251));
  XOR2_X1   g065(.A(KEYINPUT26), .B(G101), .Z(new_n252));
  XNOR2_X1  g066(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n253), .B(new_n254), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n226), .A2(new_n233), .A3(KEYINPUT68), .A4(new_n239), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n244), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT31), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n239), .B1(new_n231), .B2(new_n232), .ZN(new_n259));
  AND2_X1   g073(.A1(new_n242), .A2(KEYINPUT28), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n242), .A2(KEYINPUT28), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n259), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n255), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT71), .B(KEYINPUT31), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n244), .A2(new_n255), .A3(new_n256), .A4(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n258), .A2(new_n264), .A3(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(G472), .A2(G902), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT32), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n267), .A2(KEYINPUT32), .A3(new_n268), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n262), .A2(new_n255), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n244), .A2(new_n263), .A3(new_n256), .ZN(new_n274));
  AOI21_X1  g088(.A(KEYINPUT29), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G902), .ZN(new_n276));
  INV_X1    g090(.A(new_n216), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n239), .B1(new_n277), .B2(new_n232), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n278), .B1(new_n260), .B2(new_n261), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n255), .A2(KEYINPUT29), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n276), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(G472), .B1(new_n275), .B2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n271), .A2(new_n272), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(KEYINPUT72), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT72), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n271), .A2(new_n285), .A3(new_n272), .A4(new_n282), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(G119), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G128), .ZN(new_n289));
  INV_X1    g103(.A(G128), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(G119), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(KEYINPUT24), .B(G110), .ZN(new_n293));
  AND2_X1   g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  OR2_X1    g108(.A1(new_n294), .A2(KEYINPUT76), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(KEYINPUT76), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT23), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n291), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n290), .A2(KEYINPUT23), .A3(G119), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n298), .A2(new_n289), .A3(new_n299), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n295), .B(new_n296), .C1(G110), .C2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G140), .ZN(new_n302));
  OR2_X1    g116(.A1(new_n302), .A2(G125), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(G125), .ZN(new_n304));
  INV_X1    g118(.A(G146), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(KEYINPUT16), .B1(new_n302), .B2(G125), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT74), .B(G140), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G125), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(KEYINPUT75), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT75), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n308), .A2(new_n311), .A3(G125), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n310), .A2(new_n303), .A3(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n307), .B1(new_n313), .B2(KEYINPUT16), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n301), .B(new_n306), .C1(new_n314), .C2(new_n305), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n315), .B(KEYINPUT77), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n300), .A2(G110), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n314), .A2(new_n305), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n314), .A2(new_n305), .ZN(new_n320));
  OAI221_X1 g134(.A(new_n317), .B1(new_n292), .B2(new_n293), .C1(new_n319), .C2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n316), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n249), .A2(G221), .A3(G234), .ZN(new_n323));
  XOR2_X1   g137(.A(new_n323), .B(KEYINPUT22), .Z(new_n324));
  XNOR2_X1  g138(.A(new_n324), .B(new_n200), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n322), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n316), .A2(new_n321), .A3(new_n325), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT73), .B(G217), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n330), .B1(G234), .B2(new_n276), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n331), .A2(G902), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n327), .A2(new_n328), .A3(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n333), .B(KEYINPUT78), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n327), .A2(new_n328), .ZN(new_n335));
  OAI21_X1  g149(.A(KEYINPUT25), .B1(new_n335), .B2(G902), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT25), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n327), .A2(new_n328), .A3(new_n337), .A4(new_n276), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n336), .A2(new_n331), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n334), .A2(new_n339), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n340), .B(KEYINPUT79), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT80), .ZN(new_n342));
  AND3_X1   g156(.A1(new_n287), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n342), .B1(new_n287), .B2(new_n341), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g159(.A(KEYINPUT94), .B1(new_n319), .B2(new_n320), .ZN(new_n346));
  OR2_X1    g160(.A1(new_n314), .A2(new_n305), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT94), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n347), .A2(new_n348), .A3(new_n318), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n249), .A2(G214), .A3(new_n250), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n220), .A2(KEYINPUT92), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n220), .A2(KEYINPUT92), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n351), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n350), .A2(new_n353), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n195), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(KEYINPUT17), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n356), .A2(new_n195), .A3(new_n357), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  OR3_X1    g175(.A1(new_n361), .A2(KEYINPUT17), .A3(new_n358), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n346), .A2(new_n349), .A3(new_n359), .A4(new_n362), .ZN(new_n363));
  XNOR2_X1  g177(.A(G113), .B(G122), .ZN(new_n364));
  INV_X1    g178(.A(G104), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n364), .B(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n358), .A2(KEYINPUT18), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n313), .A2(G146), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n306), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT18), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n356), .B(new_n370), .C1(new_n351), .C2(new_n352), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n367), .A2(new_n360), .A3(new_n369), .A4(new_n371), .ZN(new_n372));
  AND3_X1   g186(.A1(new_n363), .A2(new_n366), .A3(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n366), .B1(new_n363), .B2(new_n372), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n276), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(KEYINPUT95), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT95), .ZN(new_n377));
  OAI211_X1 g191(.A(new_n377), .B(new_n276), .C1(new_n373), .C2(new_n374), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n376), .A2(G475), .A3(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n363), .A2(new_n366), .A3(new_n372), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n313), .A2(KEYINPUT19), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n303), .A2(new_n304), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n381), .B1(KEYINPUT19), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n383), .A2(G146), .ZN(new_n384));
  OAI22_X1  g198(.A1(new_n361), .A2(new_n358), .B1(new_n314), .B2(new_n305), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n372), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n366), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(KEYINPUT93), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT93), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n386), .A2(new_n390), .A3(new_n387), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n380), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G475), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n392), .A2(new_n393), .A3(new_n276), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT20), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n392), .A2(KEYINPUT20), .A3(new_n393), .A4(new_n276), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n379), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(G234), .A2(G237), .ZN(new_n399));
  AND3_X1   g213(.A1(new_n399), .A2(G952), .A3(new_n245), .ZN(new_n400));
  INV_X1    g214(.A(new_n249), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(G902), .A3(new_n399), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n402), .B(KEYINPUT99), .ZN(new_n403));
  XNOR2_X1  g217(.A(KEYINPUT21), .B(G898), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n400), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n220), .A2(G128), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT13), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(KEYINPUT96), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n290), .A2(G143), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT96), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n406), .A2(new_n411), .A3(new_n407), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n409), .A2(new_n410), .A3(new_n412), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n406), .A2(new_n407), .ZN(new_n414));
  OAI21_X1  g228(.A(G134), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n207), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n406), .A2(new_n410), .ZN(new_n417));
  INV_X1    g231(.A(G122), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(G116), .ZN(new_n419));
  INV_X1    g233(.A(G116), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(G122), .ZN(new_n421));
  AND2_X1   g235(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(G107), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AND2_X1   g238(.A1(new_n422), .A2(new_n423), .ZN(new_n425));
  OAI221_X1 g239(.A(new_n415), .B1(new_n416), .B2(new_n417), .C1(new_n424), .C2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT97), .ZN(new_n427));
  OR2_X1    g241(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  XOR2_X1   g242(.A(new_n207), .B(new_n417), .Z(new_n429));
  NAND2_X1  g243(.A1(new_n421), .A2(KEYINPUT14), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n419), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n421), .A2(KEYINPUT14), .ZN(new_n432));
  OAI21_X1  g246(.A(G107), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n425), .A2(new_n427), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n428), .A2(new_n429), .A3(new_n433), .A4(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n426), .A2(new_n435), .ZN(new_n436));
  XOR2_X1   g250(.A(KEYINPUT9), .B(G234), .Z(new_n437));
  NAND3_X1  g251(.A1(new_n437), .A2(new_n245), .A3(new_n329), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n436), .B(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n276), .ZN(new_n440));
  INV_X1    g254(.A(G478), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n441), .A2(KEYINPUT15), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n440), .B(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n443), .B(KEYINPUT98), .ZN(new_n444));
  NOR3_X1   g258(.A1(new_n398), .A2(new_n405), .A3(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(G214), .B1(G237), .B2(G902), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT91), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n228), .A2(G125), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n449), .B1(G125), .B2(new_n224), .ZN(new_n450));
  XNOR2_X1  g264(.A(KEYINPUT89), .B(G224), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n452), .A2(G953), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT7), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n450), .B(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n235), .A2(KEYINPUT5), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n288), .A2(G116), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n457), .B(G113), .C1(KEYINPUT5), .C2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n237), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(KEYINPUT3), .B1(new_n365), .B2(G107), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT3), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n462), .A2(new_n423), .A3(G104), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n461), .B(new_n463), .C1(G104), .C2(new_n423), .ZN(new_n464));
  OR2_X1    g278(.A1(new_n464), .A2(G101), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n423), .A2(G104), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n365), .A2(G107), .ZN(new_n467));
  OAI21_X1  g281(.A(G101), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n460), .A2(new_n470), .ZN(new_n471));
  XNOR2_X1  g285(.A(G110), .B(G122), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n472), .B(KEYINPUT88), .ZN(new_n473));
  XOR2_X1   g287(.A(new_n473), .B(KEYINPUT8), .Z(new_n474));
  OR2_X1    g288(.A1(new_n459), .A2(KEYINPUT87), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n459), .A2(KEYINPUT87), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n475), .A2(new_n237), .A3(new_n476), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n471), .B(new_n474), .C1(new_n470), .C2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n456), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(KEYINPUT90), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n464), .A2(G101), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n465), .A2(KEYINPUT4), .A3(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT4), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n464), .A2(new_n483), .A3(G101), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(KEYINPUT86), .B1(new_n241), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n485), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT86), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n487), .A2(new_n488), .A3(new_n239), .ZN(new_n489));
  INV_X1    g303(.A(new_n473), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n470), .A2(new_n475), .A3(new_n237), .A4(new_n476), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n486), .A2(new_n489), .A3(new_n490), .A4(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT90), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n456), .A2(new_n478), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n480), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n448), .B1(new_n495), .B2(new_n276), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(G210), .B1(G237), .B2(G902), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n486), .A2(new_n489), .A3(new_n491), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n473), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n500), .A2(KEYINPUT6), .A3(new_n492), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n450), .B(new_n453), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT6), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n499), .A2(new_n503), .A3(new_n473), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n501), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n494), .A2(new_n492), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n493), .B1(new_n456), .B2(new_n478), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n448), .B(new_n276), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n497), .A2(new_n498), .A3(new_n505), .A4(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n498), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n505), .A2(new_n508), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n510), .B1(new_n511), .B2(new_n496), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n447), .B1(new_n509), .B2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(G221), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n514), .B1(new_n437), .B2(new_n276), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT82), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n219), .A2(new_n221), .A3(new_n223), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n516), .B1(new_n469), .B2(new_n517), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n224), .A2(new_n465), .A3(KEYINPUT82), .A4(new_n468), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT10), .ZN(new_n521));
  AOI22_X1  g335(.A1(new_n520), .A2(new_n521), .B1(new_n487), .B2(new_n194), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n209), .A2(new_n215), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n470), .A2(KEYINPUT10), .A3(new_n224), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  AOI22_X1  g339(.A1(new_n518), .A2(new_n519), .B1(new_n517), .B2(new_n469), .ZN(new_n526));
  OR2_X1    g340(.A1(KEYINPUT83), .A2(KEYINPUT12), .ZN(new_n527));
  OR3_X1    g341(.A1(new_n526), .A2(new_n523), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(KEYINPUT83), .A2(KEYINPUT12), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n527), .B(new_n529), .C1(new_n526), .C2(new_n523), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n525), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n249), .A2(G227), .ZN(new_n532));
  XNOR2_X1  g346(.A(G110), .B(G140), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n532), .B(new_n533), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n534), .B(KEYINPUT81), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n531), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n520), .A2(new_n521), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n487), .A2(new_n194), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n537), .A2(new_n524), .A3(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n523), .A2(KEYINPUT84), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n540), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n542), .A2(new_n522), .A3(new_n524), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n541), .A2(new_n543), .A3(new_n534), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n536), .A2(KEYINPUT85), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(KEYINPUT85), .B1(new_n536), .B2(new_n544), .ZN(new_n546));
  OAI21_X1  g360(.A(G469), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(G469), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n548), .A2(new_n276), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n541), .A2(new_n543), .ZN(new_n550));
  INV_X1    g364(.A(new_n534), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n525), .A2(new_n528), .A3(new_n534), .A4(new_n530), .ZN(new_n553));
  AOI21_X1  g367(.A(G902), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n549), .B1(new_n554), .B2(new_n548), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n515), .B1(new_n547), .B2(new_n555), .ZN(new_n556));
  AND3_X1   g370(.A1(new_n445), .A2(new_n513), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n345), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n558), .B(G101), .ZN(G3));
  NAND2_X1  g373(.A1(new_n267), .A2(new_n276), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(G472), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(new_n269), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  AND3_X1   g377(.A1(new_n341), .A2(new_n556), .A3(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n405), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT100), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n509), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n509), .A2(new_n512), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n568), .B(new_n446), .C1(KEYINPUT100), .C2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n439), .A2(KEYINPUT101), .ZN(new_n571));
  XOR2_X1   g385(.A(new_n571), .B(KEYINPUT33), .Z(new_n572));
  NAND3_X1  g386(.A1(new_n572), .A2(G478), .A3(new_n276), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n440), .A2(new_n441), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n398), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n570), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n564), .A2(new_n565), .A3(new_n577), .ZN(new_n578));
  XOR2_X1   g392(.A(KEYINPUT34), .B(G104), .Z(new_n579));
  XNOR2_X1  g393(.A(new_n578), .B(new_n579), .ZN(G6));
  OAI21_X1  g394(.A(new_n446), .B1(new_n569), .B2(KEYINPUT100), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n581), .A2(new_n567), .ZN(new_n582));
  AND3_X1   g396(.A1(new_n379), .A2(new_n396), .A3(new_n397), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n583), .A2(new_n565), .A3(new_n444), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(KEYINPUT102), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT102), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n583), .A2(new_n586), .A3(new_n565), .A4(new_n444), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n564), .A2(new_n582), .A3(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n589), .B(KEYINPUT35), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(new_n423), .ZN(G9));
  NOR2_X1   g405(.A1(new_n326), .A2(KEYINPUT36), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n322), .B(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n332), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n339), .A2(new_n594), .ZN(new_n595));
  AND3_X1   g409(.A1(new_n557), .A2(new_n563), .A3(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(KEYINPUT37), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(G110), .ZN(G12));
  INV_X1    g412(.A(G900), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n403), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n400), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n583), .A2(new_n444), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n556), .A2(new_n595), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  AND4_X1   g419(.A1(new_n287), .A2(new_n603), .A3(new_n582), .A4(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(new_n290), .ZN(G30));
  INV_X1    g421(.A(KEYINPUT38), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n569), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n509), .A2(new_n512), .A3(KEYINPUT38), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n611), .A2(new_n447), .ZN(new_n612));
  INV_X1    g426(.A(new_n595), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n263), .B1(new_n244), .B2(new_n256), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n278), .A2(new_n242), .A3(new_n263), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n276), .ZN(new_n616));
  OAI21_X1  g430(.A(G472), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n271), .A2(new_n272), .A3(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n612), .A2(new_n613), .A3(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n602), .B(KEYINPUT39), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n556), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(KEYINPUT40), .ZN(new_n623));
  AND2_X1   g437(.A1(new_n398), .A2(new_n444), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT40), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n556), .A2(new_n625), .A3(new_n621), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n623), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(KEYINPUT103), .B1(new_n620), .B2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT103), .ZN(new_n630));
  NOR3_X1   g444(.A1(new_n619), .A2(new_n627), .A3(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(G143), .ZN(G45));
  NAND3_X1  g447(.A1(new_n398), .A2(new_n575), .A3(new_n602), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n287), .A2(new_n582), .A3(new_n605), .A4(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(KEYINPUT104), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n604), .B1(new_n284), .B2(new_n286), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT104), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n638), .A2(new_n639), .A3(new_n582), .A4(new_n635), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(G146), .ZN(G48));
  OR2_X1    g456(.A1(new_n554), .A2(new_n548), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n554), .A2(new_n548), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n515), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n648), .A2(new_n405), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n577), .A2(new_n287), .A3(new_n341), .A4(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(KEYINPUT41), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G113), .ZN(G15));
  NOR2_X1   g466(.A1(new_n570), .A2(new_n648), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n588), .A2(new_n287), .A3(new_n341), .A4(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G116), .ZN(G18));
  NAND4_X1  g469(.A1(new_n653), .A2(new_n287), .A3(new_n445), .A4(new_n595), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G119), .ZN(G21));
  AND2_X1   g471(.A1(new_n582), .A2(new_n624), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n334), .A2(new_n339), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n561), .A2(KEYINPUT106), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT106), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n560), .A2(new_n661), .A3(G472), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n279), .A2(new_n263), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n258), .A2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT105), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n258), .A2(KEYINPUT105), .A3(new_n664), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n667), .A2(new_n266), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n268), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n663), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n658), .A2(new_n659), .A3(new_n649), .A4(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G122), .ZN(G24));
  AOI21_X1  g487(.A(new_n661), .B1(new_n560), .B2(G472), .ZN(new_n674));
  INV_X1    g488(.A(G472), .ZN(new_n675));
  AOI211_X1 g489(.A(KEYINPUT106), .B(new_n675), .C1(new_n267), .C2(new_n276), .ZN(new_n676));
  OAI211_X1 g490(.A(new_n670), .B(new_n595), .C1(new_n674), .C2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT107), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n663), .A2(KEYINPUT107), .A3(new_n595), .A4(new_n670), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n634), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n653), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT108), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n681), .A2(KEYINPUT108), .A3(new_n653), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G125), .ZN(G27));
  NOR2_X1   g501(.A1(new_n569), .A2(new_n447), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n536), .A2(KEYINPUT109), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT109), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n531), .A2(new_n690), .A3(new_n535), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n689), .A2(G469), .A3(new_n544), .A4(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n555), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n647), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT110), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n693), .A2(KEYINPUT110), .A3(new_n647), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n635), .A2(new_n688), .A3(new_n696), .A4(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n283), .A2(new_n659), .ZN(new_n699));
  OAI21_X1  g513(.A(KEYINPUT42), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n696), .A2(new_n697), .ZN(new_n701));
  INV_X1    g515(.A(new_n688), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n634), .A2(KEYINPUT42), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n703), .A2(new_n287), .A3(new_n341), .A4(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n700), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(new_n195), .ZN(G33));
  NAND4_X1  g521(.A1(new_n703), .A2(new_n287), .A3(new_n341), .A4(new_n603), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G134), .ZN(G36));
  NOR3_X1   g523(.A1(new_n545), .A2(new_n546), .A3(KEYINPUT45), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n689), .A2(KEYINPUT45), .A3(new_n544), .A4(new_n691), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(G469), .ZN(new_n712));
  OAI22_X1  g526(.A1(new_n710), .A2(new_n712), .B1(new_n548), .B2(new_n276), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT46), .ZN(new_n714));
  AOI22_X1  g528(.A1(new_n713), .A2(new_n714), .B1(new_n548), .B2(new_n554), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n715), .B1(new_n714), .B2(new_n713), .ZN(new_n716));
  AND3_X1   g530(.A1(new_n716), .A2(new_n647), .A3(new_n621), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT43), .ZN(new_n718));
  INV_X1    g532(.A(new_n575), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n718), .B1(new_n719), .B2(new_n398), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n583), .A2(KEYINPUT43), .A3(new_n575), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n722), .A2(new_n562), .A3(new_n595), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT44), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n722), .A2(KEYINPUT44), .A3(new_n562), .A4(new_n595), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n717), .A2(new_n725), .A3(new_n688), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G137), .ZN(G39));
  NAND2_X1  g542(.A1(new_n716), .A2(new_n647), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT111), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n730), .A2(KEYINPUT47), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  AND2_X1   g547(.A1(new_n730), .A2(KEYINPUT47), .ZN(new_n734));
  OAI211_X1 g548(.A(new_n716), .B(new_n647), .C1(new_n731), .C2(new_n734), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n287), .A2(new_n341), .A3(new_n634), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n733), .A2(new_n688), .A3(new_n735), .A4(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(KEYINPUT112), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(new_n302), .ZN(G42));
  AOI21_X1  g553(.A(new_n601), .B1(new_n720), .B2(new_n721), .ZN(new_n740));
  AND3_X1   g554(.A1(new_n740), .A2(new_n659), .A3(new_n671), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n733), .A2(new_n735), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n646), .A2(new_n515), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n702), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT117), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n745), .B1(new_n648), .B2(new_n446), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n646), .A2(KEYINPUT117), .A3(new_n447), .A4(new_n647), .ZN(new_n747));
  AND3_X1   g561(.A1(new_n746), .A2(new_n611), .A3(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT118), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT50), .ZN(new_n750));
  AND3_X1   g564(.A1(new_n748), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n741), .B1(new_n744), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n679), .A2(new_n680), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n702), .A2(new_n648), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n753), .A2(new_n754), .A3(new_n740), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n618), .A2(new_n601), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n754), .A2(new_n341), .A3(new_n756), .ZN(new_n757));
  NOR3_X1   g571(.A1(new_n757), .A2(new_n398), .A3(new_n575), .ZN(new_n758));
  AOI22_X1  g572(.A1(new_n741), .A2(new_n748), .B1(new_n749), .B2(new_n750), .ZN(new_n759));
  NAND2_X1  g573(.A1(KEYINPUT118), .A2(KEYINPUT50), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n758), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n752), .A2(new_n755), .A3(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT51), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  AND4_X1   g578(.A1(new_n283), .A2(new_n740), .A3(new_n659), .A4(new_n754), .ZN(new_n765));
  XOR2_X1   g579(.A(new_n765), .B(KEYINPUT48), .Z(new_n766));
  INV_X1    g580(.A(G952), .ZN(new_n767));
  AOI211_X1 g581(.A(new_n767), .B(G953), .C1(new_n741), .C2(new_n653), .ZN(new_n768));
  OAI211_X1 g582(.A(new_n766), .B(new_n768), .C1(new_n576), .C2(new_n757), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT119), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n762), .A2(new_n763), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n764), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n596), .B1(new_n345), .B2(new_n557), .ZN(new_n774));
  AND3_X1   g588(.A1(new_n700), .A2(new_n705), .A3(new_n708), .ZN(new_n775));
  AOI211_X1 g589(.A(new_n634), .B(new_n701), .C1(new_n679), .C2(new_n680), .ZN(new_n776));
  INV_X1    g590(.A(new_n443), .ZN(new_n777));
  AND4_X1   g591(.A1(new_n583), .A2(new_n638), .A3(new_n777), .A4(new_n602), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n688), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n576), .B1(new_n398), .B2(new_n777), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n564), .A2(new_n513), .A3(new_n565), .A4(new_n780), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n774), .A2(new_n775), .A3(new_n779), .A4(new_n781), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n606), .B1(new_n637), .B2(new_n640), .ZN(new_n783));
  INV_X1    g597(.A(new_n694), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n602), .B(KEYINPUT115), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n595), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n658), .A2(new_n618), .A3(new_n784), .A4(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(KEYINPUT108), .B1(new_n681), .B2(new_n653), .ZN(new_n788));
  AND4_X1   g602(.A1(KEYINPUT108), .A2(new_n753), .A3(new_n635), .A4(new_n653), .ZN(new_n789));
  OAI211_X1 g603(.A(new_n783), .B(new_n787), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n686), .A2(KEYINPUT52), .A3(new_n783), .A4(new_n787), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n782), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n672), .A2(new_n654), .A3(new_n650), .A4(new_n656), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(KEYINPUT114), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(KEYINPUT53), .ZN(new_n798));
  XNOR2_X1  g612(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n794), .A2(new_n796), .A3(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n798), .A2(KEYINPUT54), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n797), .A2(new_n800), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT53), .ZN(new_n804));
  OR2_X1    g618(.A1(new_n795), .A2(new_n804), .ZN(new_n805));
  AOI211_X1 g619(.A(new_n782), .B(new_n805), .C1(new_n792), .C2(new_n793), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n803), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n773), .A2(new_n802), .A3(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n769), .A2(new_n770), .ZN(new_n811));
  OAI22_X1  g625(.A1(new_n810), .A2(new_n811), .B1(G952), .B2(G953), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n719), .A2(new_n398), .A3(new_n447), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n813), .A2(new_n659), .A3(new_n647), .ZN(new_n814));
  XOR2_X1   g628(.A(new_n814), .B(KEYINPUT113), .Z(new_n815));
  INV_X1    g629(.A(KEYINPUT49), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n618), .B1(new_n816), .B2(new_n646), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n645), .A2(KEYINPUT49), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n815), .A2(new_n611), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n812), .A2(new_n819), .ZN(G75));
  AOI21_X1  g634(.A(new_n799), .B1(new_n794), .B2(new_n796), .ZN(new_n821));
  OAI211_X1 g635(.A(G210), .B(G902), .C1(new_n821), .C2(new_n806), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT56), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n501), .A2(new_n504), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(new_n502), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(KEYINPUT120), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(KEYINPUT55), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n822), .A2(KEYINPUT121), .A3(new_n823), .A4(new_n827), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n249), .A2(G952), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(KEYINPUT122), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n822), .A2(new_n823), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT121), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(new_n827), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n822), .A2(KEYINPUT121), .A3(new_n823), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n832), .B1(new_n836), .B2(new_n837), .ZN(G51));
  XNOR2_X1  g652(.A(new_n549), .B(KEYINPUT57), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n808), .B1(new_n803), .B2(new_n807), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n821), .A2(new_n806), .A3(KEYINPUT54), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n839), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n552), .A2(new_n553), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n821), .A2(new_n806), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n845), .A2(new_n276), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n710), .A2(new_n712), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n829), .B1(new_n844), .B2(new_n848), .ZN(G54));
  INV_X1    g663(.A(new_n392), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n803), .A2(new_n807), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n851), .A2(KEYINPUT58), .A3(G902), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n850), .B1(new_n852), .B2(new_n393), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n846), .A2(KEYINPUT58), .A3(G475), .A4(new_n392), .ZN(new_n854));
  INV_X1    g668(.A(new_n829), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(G60));
  NAND2_X1  g670(.A1(new_n809), .A2(new_n802), .ZN(new_n857));
  NAND2_X1  g671(.A1(G478), .A2(G902), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n858), .B(KEYINPUT59), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n572), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n572), .A2(new_n859), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n851), .A2(KEYINPUT54), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n861), .B1(new_n862), .B2(new_n809), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n860), .A2(new_n863), .A3(new_n830), .ZN(G63));
  INV_X1    g678(.A(KEYINPUT61), .ZN(new_n865));
  NAND2_X1  g679(.A1(G217), .A2(G902), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(KEYINPUT60), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  XOR2_X1   g682(.A(new_n593), .B(KEYINPUT123), .Z(new_n869));
  OAI211_X1 g683(.A(new_n868), .B(new_n869), .C1(new_n821), .C2(new_n806), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n867), .B1(new_n803), .B2(new_n807), .ZN(new_n871));
  INV_X1    g685(.A(new_n335), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n865), .B1(new_n873), .B2(new_n830), .ZN(new_n874));
  OAI21_X1  g688(.A(KEYINPUT124), .B1(new_n871), .B2(new_n872), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n870), .A2(KEYINPUT61), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT124), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n877), .B(new_n335), .C1(new_n845), .C2(new_n867), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n875), .A2(new_n876), .A3(new_n831), .A4(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n874), .A2(new_n879), .ZN(G66));
  OAI21_X1  g694(.A(G953), .B1(new_n452), .B2(new_n404), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n774), .A2(new_n781), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n796), .A2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n881), .B1(new_n884), .B2(new_n401), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n824), .B1(G898), .B2(new_n249), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT125), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n885), .B(new_n887), .ZN(G69));
  AND2_X1   g702(.A1(new_n226), .A2(new_n233), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n889), .B(new_n383), .Z(new_n890));
  NOR2_X1   g704(.A1(new_n249), .A2(new_n599), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT126), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n775), .A2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n708), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n706), .A2(new_n895), .A3(KEYINPUT126), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n727), .B(new_n737), .C1(new_n894), .C2(new_n896), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n717), .A2(new_n283), .A3(new_n659), .A4(new_n658), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n686), .A2(new_n783), .A3(new_n898), .ZN(new_n899));
  OR2_X1    g713(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n890), .B(new_n892), .C1(new_n900), .C2(new_n401), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT127), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n737), .A2(new_n727), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n632), .A2(new_n686), .A3(new_n783), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT62), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n632), .A2(new_n686), .A3(KEYINPUT62), .A4(new_n783), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n903), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(new_n622), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n345), .A2(new_n909), .A3(new_n688), .A4(new_n780), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n401), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n901), .B(new_n902), .C1(new_n911), .C2(new_n890), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n906), .A2(new_n907), .ZN(new_n913));
  INV_X1    g727(.A(new_n903), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n913), .A2(new_n910), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n890), .B1(new_n915), .B2(new_n249), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n897), .A2(new_n899), .A3(new_n401), .ZN(new_n917));
  INV_X1    g731(.A(new_n890), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n917), .A2(new_n918), .A3(new_n891), .ZN(new_n919));
  OAI21_X1  g733(.A(KEYINPUT127), .B1(new_n916), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n249), .B1(G227), .B2(G900), .ZN(new_n921));
  AND3_X1   g735(.A1(new_n912), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n921), .B1(new_n912), .B2(new_n920), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n922), .A2(new_n923), .ZN(G72));
  NAND2_X1  g738(.A1(G472), .A2(G902), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT63), .Z(new_n926));
  OAI21_X1  g740(.A(new_n926), .B1(new_n915), .B2(new_n883), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n614), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n926), .B1(new_n900), .B2(new_n883), .ZN(new_n929));
  INV_X1    g743(.A(new_n274), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n928), .A2(new_n855), .A3(new_n931), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n798), .A2(new_n801), .ZN(new_n933));
  INV_X1    g747(.A(new_n926), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n930), .A2(new_n614), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n932), .B1(new_n933), .B2(new_n935), .ZN(G57));
endmodule


