//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 1 0 0 0 0 0 0 0 1 0 1 1 0 1 0 0 0 0 0 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 1 1 1 1 0 1 0 1 0 0 1 1 1 1 0 0 0 1 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n598, new_n599, new_n600, new_n601,
    new_n603, new_n604, new_n605, new_n606, new_n608, new_n609, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n656, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n762, new_n763, new_n764, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n833, new_n834, new_n836, new_n837, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n855, new_n856,
    new_n857, new_n858, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n887, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  OAI21_X1  g001(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT64), .ZN(new_n204));
  NAND2_X1  g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205));
  OR2_X1    g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206));
  OAI211_X1 g005(.A(new_n204), .B(new_n205), .C1(KEYINPUT26), .C2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT65), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n207), .A2(KEYINPUT65), .A3(new_n208), .ZN(new_n212));
  XNOR2_X1  g011(.A(KEYINPUT27), .B(G183gat), .ZN(new_n213));
  INV_X1    g012(.A(G190gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  XOR2_X1   g014(.A(new_n215), .B(KEYINPUT28), .Z(new_n216));
  NAND3_X1  g015(.A1(new_n211), .A2(new_n212), .A3(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(G127gat), .B(G134gat), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n218), .B(KEYINPUT68), .ZN(new_n219));
  XOR2_X1   g018(.A(KEYINPUT67), .B(G120gat), .Z(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G113gat), .ZN(new_n221));
  INV_X1    g020(.A(G113gat), .ZN(new_n222));
  INV_X1    g021(.A(G120gat), .ZN(new_n223));
  AOI21_X1  g022(.A(KEYINPUT1), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n219), .A2(new_n221), .A3(new_n224), .ZN(new_n225));
  XOR2_X1   g024(.A(KEYINPUT66), .B(G127gat), .Z(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(G134gat), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n224), .B1(new_n222), .B2(new_n223), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n227), .B(new_n228), .C1(G127gat), .C2(G134gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n225), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n206), .B(KEYINPUT23), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n208), .A2(KEYINPUT24), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n233), .B1(G169gat), .B2(G176gat), .ZN(new_n234));
  OR2_X1    g033(.A1(G183gat), .A2(G190gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n235), .A2(KEYINPUT24), .A3(new_n208), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n232), .A2(new_n234), .A3(new_n236), .ZN(new_n237));
  XOR2_X1   g036(.A(new_n237), .B(KEYINPUT25), .Z(new_n238));
  NAND3_X1  g037(.A1(new_n217), .A2(new_n231), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT69), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n217), .A2(KEYINPUT69), .A3(new_n238), .A4(new_n231), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n217), .A2(new_n238), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(new_n230), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n241), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(G227gat), .A2(G233gat), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  OR3_X1    g046(.A1(new_n245), .A2(KEYINPUT34), .A3(new_n247), .ZN(new_n248));
  OAI21_X1  g047(.A(KEYINPUT34), .B1(new_n245), .B2(new_n247), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT33), .B1(new_n245), .B2(new_n247), .ZN(new_n251));
  XNOR2_X1  g050(.A(G71gat), .B(G99gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n252), .B(KEYINPUT70), .ZN(new_n253));
  INV_X1    g052(.A(G15gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n255), .B(G43gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n251), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n250), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n245), .A2(new_n247), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT32), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n248), .B(new_n249), .C1(new_n251), .C2(new_n256), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n258), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n261), .B1(new_n258), .B2(new_n262), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n202), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n265), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n267), .A2(KEYINPUT36), .A3(new_n263), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  AND2_X1   g068(.A1(G226gat), .A2(G233gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n243), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(KEYINPUT29), .B1(new_n217), .B2(new_n238), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n271), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(G197gat), .B(G204gat), .ZN(new_n274));
  INV_X1    g073(.A(G211gat), .ZN(new_n275));
  INV_X1    g074(.A(G218gat), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n274), .B1(KEYINPUT22), .B2(new_n277), .ZN(new_n278));
  XOR2_X1   g077(.A(G211gat), .B(G218gat), .Z(new_n279));
  XNOR2_X1  g078(.A(new_n278), .B(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n280), .B(KEYINPUT71), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n273), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n281), .ZN(new_n283));
  OAI211_X1 g082(.A(new_n271), .B(new_n283), .C1(new_n270), .C2(new_n272), .ZN(new_n284));
  XNOR2_X1  g083(.A(G8gat), .B(G36gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(G64gat), .B(G92gat), .ZN(new_n286));
  XOR2_X1   g085(.A(new_n285), .B(new_n286), .Z(new_n287));
  AND3_X1   g086(.A1(new_n282), .A2(new_n284), .A3(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT72), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT30), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n282), .A2(new_n284), .ZN(new_n292));
  INV_X1    g091(.A(new_n287), .ZN(new_n293));
  OAI21_X1  g092(.A(KEYINPUT72), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n290), .A2(new_n291), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n287), .B1(new_n282), .B2(new_n284), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n296), .B1(new_n288), .B2(KEYINPUT30), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(G155gat), .ZN(new_n299));
  INV_X1    g098(.A(G162gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(G155gat), .A2(G162gat), .ZN(new_n302));
  AND2_X1   g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  XOR2_X1   g102(.A(KEYINPUT73), .B(KEYINPUT2), .Z(new_n304));
  XNOR2_X1  g103(.A(G141gat), .B(G148gat), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n303), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT74), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n306), .B(new_n307), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n302), .B1(new_n301), .B2(KEYINPUT2), .ZN(new_n309));
  INV_X1    g108(.A(G141gat), .ZN(new_n310));
  OAI21_X1  g109(.A(KEYINPUT75), .B1(new_n310), .B2(G148gat), .ZN(new_n311));
  INV_X1    g110(.A(G148gat), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n311), .B1(G141gat), .B2(new_n312), .ZN(new_n313));
  NOR3_X1   g112(.A1(new_n310), .A2(KEYINPUT75), .A3(G148gat), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n309), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  AND2_X1   g114(.A1(new_n308), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(new_n231), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(KEYINPUT4), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT4), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n316), .A2(new_n319), .A3(new_n231), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n308), .A2(new_n315), .ZN(new_n322));
  OR2_X1    g121(.A1(new_n322), .A2(KEYINPUT3), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(KEYINPUT3), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n323), .A2(new_n324), .A3(new_n230), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT39), .ZN(new_n327));
  NAND2_X1  g126(.A1(G225gat), .A2(G233gat), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n326), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  XOR2_X1   g129(.A(G1gat), .B(G29gat), .Z(new_n331));
  XNOR2_X1  g130(.A(G57gat), .B(G85gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n331), .B(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n334));
  XOR2_X1   g133(.A(new_n333), .B(new_n334), .Z(new_n335));
  NAND2_X1  g134(.A1(new_n330), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n231), .B(new_n322), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(new_n328), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(KEYINPUT39), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n339), .B1(new_n329), .B2(new_n326), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT40), .ZN(new_n341));
  OR3_X1    g140(.A1(new_n336), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n341), .B1(new_n336), .B2(new_n340), .ZN(new_n343));
  INV_X1    g142(.A(new_n335), .ZN(new_n344));
  OAI21_X1  g143(.A(KEYINPUT5), .B1(new_n337), .B2(new_n328), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT77), .ZN(new_n346));
  OR2_X1    g145(.A1(new_n320), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n318), .A2(KEYINPUT76), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n320), .A2(new_n346), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT76), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n317), .A2(new_n350), .A3(KEYINPUT4), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n347), .A2(new_n348), .A3(new_n349), .A4(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n325), .A2(new_n328), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n345), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n321), .ZN(new_n356));
  NOR3_X1   g155(.A1(new_n356), .A2(new_n353), .A3(KEYINPUT5), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n344), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  AND2_X1   g157(.A1(new_n343), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n298), .A2(new_n342), .A3(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT29), .ZN(new_n361));
  AOI21_X1  g160(.A(KEYINPUT3), .B1(new_n280), .B2(new_n361), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n316), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n323), .A2(new_n361), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n363), .B1(new_n364), .B2(new_n281), .ZN(new_n365));
  XNOR2_X1  g164(.A(G78gat), .B(G106gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n365), .B(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(G228gat), .A2(G233gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n368), .B(G22gat), .ZN(new_n369));
  XOR2_X1   g168(.A(KEYINPUT31), .B(G50gat), .Z(new_n370));
  XNOR2_X1  g169(.A(new_n369), .B(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n367), .B(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n287), .B1(new_n292), .B2(KEYINPUT37), .ZN(new_n374));
  XOR2_X1   g173(.A(KEYINPUT81), .B(KEYINPUT38), .Z(new_n375));
  INV_X1    g174(.A(KEYINPUT37), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n282), .A2(new_n376), .A3(new_n284), .ZN(new_n377));
  AND3_X1   g176(.A1(new_n374), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n375), .B1(new_n374), .B2(new_n377), .ZN(new_n379));
  OAI211_X1 g178(.A(new_n294), .B(new_n290), .C1(new_n378), .C2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT80), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT6), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n381), .B1(new_n358), .B2(new_n382), .ZN(new_n383));
  OR3_X1    g182(.A1(new_n356), .A2(new_n353), .A3(KEYINPUT5), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n348), .A2(new_n351), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n320), .B(KEYINPUT77), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n353), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n335), .B(new_n384), .C1(new_n387), .C2(new_n345), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n388), .A2(new_n358), .A3(new_n382), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n384), .B1(new_n387), .B2(new_n345), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n390), .A2(KEYINPUT80), .A3(KEYINPUT6), .A4(new_n344), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n383), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n360), .B(new_n373), .C1(new_n380), .C2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n389), .A2(KEYINPUT79), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT79), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n388), .A2(new_n358), .A3(new_n395), .A4(new_n382), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  AND2_X1   g196(.A1(new_n383), .A2(new_n391), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n298), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n269), .B(new_n393), .C1(new_n399), .C2(new_n373), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n397), .A2(new_n398), .ZN(new_n402));
  NOR3_X1   g201(.A1(new_n264), .A2(new_n265), .A3(new_n372), .ZN(new_n403));
  INV_X1    g202(.A(new_n298), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT35), .ZN(new_n406));
  AND3_X1   g205(.A1(new_n392), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  AOI22_X1  g206(.A1(new_n405), .A2(KEYINPUT35), .B1(new_n403), .B2(new_n407), .ZN(new_n408));
  OR2_X1    g207(.A1(new_n401), .A2(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(G113gat), .B(G141gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n410), .B(G197gat), .ZN(new_n411));
  XOR2_X1   g210(.A(KEYINPUT11), .B(G169gat), .Z(new_n412));
  XNOR2_X1  g211(.A(new_n411), .B(new_n412), .ZN(new_n413));
  XOR2_X1   g212(.A(new_n413), .B(KEYINPUT12), .Z(new_n414));
  XNOR2_X1  g213(.A(KEYINPUT83), .B(G36gat), .ZN(new_n415));
  INV_X1    g214(.A(G29gat), .ZN(new_n416));
  OAI21_X1  g215(.A(KEYINPUT84), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT84), .ZN(new_n418));
  INV_X1    g217(.A(G36gat), .ZN(new_n419));
  AND2_X1   g218(.A1(new_n419), .A2(KEYINPUT83), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n419), .A2(KEYINPUT83), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n418), .B(G29gat), .C1(new_n420), .C2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT14), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n423), .B(KEYINPUT82), .C1(G29gat), .C2(G36gat), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT82), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n425), .A2(new_n416), .A3(new_n419), .ZN(new_n426));
  OAI21_X1  g225(.A(KEYINPUT82), .B1(G29gat), .B2(G36gat), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n426), .A2(KEYINPUT14), .A3(new_n427), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n417), .A2(new_n422), .A3(new_n424), .A4(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(G43gat), .B(G50gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n430), .B(KEYINPUT15), .ZN(new_n431));
  OR2_X1    g230(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  AND2_X1   g231(.A1(new_n430), .A2(KEYINPUT15), .ZN(new_n433));
  AND3_X1   g232(.A1(new_n429), .A2(KEYINPUT85), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(KEYINPUT85), .B1(new_n429), .B2(new_n433), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n432), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT86), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT86), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n438), .B(new_n432), .C1(new_n434), .C2(new_n435), .ZN(new_n439));
  XNOR2_X1  g238(.A(KEYINPUT87), .B(KEYINPUT17), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n437), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(KEYINPUT88), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT88), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n437), .A2(new_n443), .A3(new_n439), .A4(new_n440), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(G8gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(G15gat), .B(G22gat), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT89), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n447), .B(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(G1gat), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT16), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n446), .B1(new_n452), .B2(KEYINPUT90), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n452), .B1(G1gat), .B2(new_n449), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OAI221_X1 g254(.A(new_n452), .B1(KEYINPUT90), .B2(new_n446), .C1(G1gat), .C2(new_n449), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n436), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n457), .B1(new_n458), .B2(KEYINPUT17), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n445), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT91), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n455), .A2(KEYINPUT91), .A3(new_n456), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n462), .A2(new_n437), .A3(new_n439), .A4(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(G229gat), .A2(G233gat), .ZN(new_n465));
  AND2_X1   g264(.A1(new_n465), .A2(KEYINPUT18), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n460), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  XOR2_X1   g266(.A(new_n465), .B(KEYINPUT13), .Z(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n462), .A2(new_n463), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n437), .A2(new_n439), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n469), .B1(new_n472), .B2(new_n464), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n467), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n464), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n478), .B1(new_n445), .B2(new_n459), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n477), .B1(new_n479), .B2(new_n465), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n414), .B1(new_n475), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT93), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n460), .A2(new_n465), .A3(new_n464), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(new_n476), .ZN(new_n484));
  INV_X1    g283(.A(new_n414), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n473), .B1(new_n479), .B2(new_n466), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n481), .A2(new_n482), .A3(new_n487), .ZN(new_n488));
  OAI211_X1 g287(.A(KEYINPUT93), .B(new_n414), .C1(new_n475), .C2(new_n480), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT94), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n488), .A2(new_n489), .A3(KEYINPUT94), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AND2_X1   g293(.A1(new_n409), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n496), .B(KEYINPUT95), .ZN(new_n497));
  XOR2_X1   g296(.A(G57gat), .B(G64gat), .Z(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  XOR2_X1   g298(.A(G71gat), .B(G78gat), .Z(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n500), .ZN(new_n502));
  INV_X1    g301(.A(G57gat), .ZN(new_n503));
  INV_X1    g302(.A(G64gat), .ZN(new_n504));
  OR3_X1    g303(.A1(new_n503), .A2(new_n504), .A3(KEYINPUT96), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n504), .B1(new_n503), .B2(KEYINPUT96), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n497), .A2(new_n502), .A3(new_n505), .A4(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n501), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT97), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT97), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n501), .A2(new_n510), .A3(new_n507), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n512), .A2(KEYINPUT21), .ZN(new_n513));
  NAND2_X1  g312(.A1(G231gat), .A2(G233gat), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n513), .B(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n515), .B(G127gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n512), .A2(KEYINPUT21), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n470), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n516), .B(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n520), .B(G155gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(G183gat), .B(G211gat), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n521), .B(new_n522), .ZN(new_n523));
  OR2_X1    g322(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n519), .A2(new_n523), .ZN(new_n525));
  AND2_X1   g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(G232gat), .A2(G233gat), .ZN(new_n528));
  XOR2_X1   g327(.A(new_n528), .B(KEYINPUT98), .Z(new_n529));
  INV_X1    g328(.A(KEYINPUT41), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(G134gat), .B(G162gat), .ZN(new_n532));
  XOR2_X1   g331(.A(new_n531), .B(new_n532), .Z(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  XOR2_X1   g333(.A(KEYINPUT100), .B(G85gat), .Z(new_n535));
  INV_X1    g334(.A(G92gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(G99gat), .A2(G106gat), .ZN(new_n537));
  AOI22_X1  g336(.A1(new_n535), .A2(new_n536), .B1(KEYINPUT8), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT99), .ZN(new_n539));
  INV_X1    g338(.A(G85gat), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n539), .B1(new_n540), .B2(new_n536), .ZN(new_n541));
  NAND3_X1  g340(.A1(KEYINPUT99), .A2(G85gat), .A3(G92gat), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n541), .A2(KEYINPUT7), .A3(new_n542), .ZN(new_n543));
  OR2_X1    g342(.A1(new_n541), .A2(KEYINPUT7), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n538), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(G99gat), .B(G106gat), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT101), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n538), .A2(new_n546), .A3(new_n543), .A4(new_n544), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n545), .A2(KEYINPUT101), .A3(new_n547), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n553), .B1(new_n458), .B2(KEYINPUT17), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n445), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n553), .ZN(new_n556));
  OAI22_X1  g355(.A1(new_n471), .A2(new_n556), .B1(new_n530), .B2(new_n529), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(G190gat), .B(G218gat), .ZN(new_n560));
  XOR2_X1   g359(.A(new_n560), .B(KEYINPUT102), .Z(new_n561));
  NAND2_X1  g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n559), .A2(new_n561), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n534), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n564), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n566), .A2(new_n533), .A3(new_n562), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n527), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(G230gat), .A2(G233gat), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT10), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n548), .A2(new_n501), .A3(new_n507), .A4(new_n550), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n572), .B(new_n573), .C1(new_n553), .C2(new_n512), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n553), .A2(new_n512), .A3(KEYINPUT10), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n571), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n573), .B1(new_n553), .B2(new_n512), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n576), .B1(new_n571), .B2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT104), .ZN(new_n579));
  XOR2_X1   g378(.A(G120gat), .B(G148gat), .Z(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(KEYINPUT103), .ZN(new_n581));
  XNOR2_X1  g380(.A(G176gat), .B(G204gat), .ZN(new_n582));
  XOR2_X1   g381(.A(new_n581), .B(new_n582), .Z(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n578), .A2(new_n579), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n577), .A2(new_n571), .ZN(new_n586));
  AND2_X1   g385(.A1(new_n574), .A2(new_n575), .ZN(new_n587));
  OAI211_X1 g386(.A(new_n586), .B(new_n584), .C1(new_n587), .C2(new_n571), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(KEYINPUT104), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  OR2_X1    g389(.A1(new_n578), .A2(new_n584), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n569), .A2(new_n592), .ZN(new_n593));
  AND2_X1   g392(.A1(new_n495), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n402), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g396(.A(KEYINPUT16), .B(G8gat), .Z(new_n598));
  AND3_X1   g397(.A1(new_n594), .A2(new_n298), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n446), .B1(new_n594), .B2(new_n298), .ZN(new_n600));
  OAI21_X1  g399(.A(KEYINPUT42), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n601), .B1(KEYINPUT42), .B2(new_n599), .ZN(G1325gat));
  NOR2_X1   g401(.A1(new_n264), .A2(new_n265), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n594), .A2(new_n254), .A3(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n269), .ZN(new_n605));
  AND2_X1   g404(.A1(new_n594), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n604), .B1(new_n606), .B2(new_n254), .ZN(G1326gat));
  NAND2_X1  g406(.A1(new_n594), .A2(new_n372), .ZN(new_n608));
  XNOR2_X1  g407(.A(KEYINPUT43), .B(G22gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(G1327gat));
  INV_X1    g409(.A(new_n592), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n526), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n612), .A2(new_n568), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n495), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n614), .A2(new_n416), .A3(new_n595), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT45), .ZN(new_n616));
  INV_X1    g415(.A(new_n568), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n617), .B1(new_n401), .B2(new_n408), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT44), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI211_X1 g419(.A(KEYINPUT44), .B(new_n617), .C1(new_n401), .C2(new_n408), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NOR3_X1   g421(.A1(new_n622), .A2(new_n490), .A3(new_n612), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g423(.A(G29gat), .B1(new_n624), .B2(new_n402), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n616), .A2(new_n625), .ZN(G1328gat));
  NAND3_X1  g425(.A1(new_n614), .A2(new_n298), .A3(new_n415), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n627), .B(KEYINPUT46), .Z(new_n628));
  NOR2_X1   g427(.A1(new_n624), .A2(new_n404), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n628), .B1(new_n415), .B2(new_n629), .ZN(G1329gat));
  OAI21_X1  g429(.A(G43gat), .B1(new_n624), .B2(new_n269), .ZN(new_n631));
  INV_X1    g430(.A(new_n603), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n632), .A2(G43gat), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n495), .A2(new_n613), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT105), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT47), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(G1330gat));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n372), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n373), .A2(G50gat), .ZN(new_n640));
  AOI22_X1  g439(.A1(new_n639), .A2(G50gat), .B1(new_n614), .B2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g441(.A(new_n490), .ZN(new_n643));
  NOR3_X1   g442(.A1(new_n569), .A2(new_n643), .A3(new_n611), .ZN(new_n644));
  AND2_X1   g443(.A1(new_n409), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(new_n595), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(G57gat), .ZN(G1332gat));
  INV_X1    g446(.A(KEYINPUT49), .ZN(new_n648));
  OAI211_X1 g447(.A(new_n645), .B(new_n298), .C1(new_n648), .C2(new_n504), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n504), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(G1333gat));
  NAND2_X1  g450(.A1(new_n645), .A2(new_n605), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n632), .A2(G71gat), .ZN(new_n653));
  AOI22_X1  g452(.A1(new_n652), .A2(G71gat), .B1(new_n645), .B2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g454(.A1(new_n645), .A2(new_n372), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g456(.A1(new_n526), .A2(new_n490), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT106), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n526), .A2(KEYINPUT106), .A3(new_n490), .ZN(new_n661));
  AND2_X1   g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n662), .A2(new_n611), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n620), .A2(new_n621), .A3(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT107), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n620), .A2(new_n663), .A3(KEYINPUT107), .A4(new_n621), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n666), .A2(new_n595), .A3(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT108), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n535), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n670), .B1(new_n669), .B2(new_n668), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT51), .ZN(new_n672));
  OR3_X1    g471(.A1(new_n618), .A2(new_n672), .A3(new_n662), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n672), .B1(new_n618), .B2(new_n662), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n611), .B1(new_n675), .B2(KEYINPUT109), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n676), .B1(KEYINPUT109), .B2(new_n675), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n595), .A2(new_n535), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n671), .B1(new_n677), .B2(new_n678), .ZN(G1336gat));
  AOI21_X1  g478(.A(new_n611), .B1(new_n673), .B2(new_n674), .ZN(new_n680));
  AND3_X1   g479(.A1(new_n680), .A2(new_n536), .A3(new_n298), .ZN(new_n681));
  INV_X1    g480(.A(new_n664), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n536), .B1(new_n682), .B2(new_n298), .ZN(new_n683));
  OR3_X1    g482(.A1(new_n681), .A2(KEYINPUT52), .A3(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n666), .A2(new_n298), .A3(new_n667), .ZN(new_n685));
  AND3_X1   g484(.A1(new_n685), .A2(KEYINPUT110), .A3(G92gat), .ZN(new_n686));
  AOI21_X1  g485(.A(KEYINPUT110), .B1(new_n685), .B2(G92gat), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n686), .A2(new_n687), .A3(new_n681), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT52), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n684), .B1(new_n688), .B2(new_n689), .ZN(G1337gat));
  NAND3_X1  g489(.A1(new_n666), .A2(new_n605), .A3(new_n667), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(G99gat), .ZN(new_n692));
  OR2_X1    g491(.A1(new_n632), .A2(G99gat), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n692), .B1(new_n677), .B2(new_n693), .ZN(G1338gat));
  NOR2_X1   g493(.A1(new_n373), .A2(G106gat), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n695), .ZN(new_n696));
  OR2_X1    g495(.A1(new_n696), .A2(KEYINPUT112), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(KEYINPUT112), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n372), .ZN(new_n699));
  AOI21_X1  g498(.A(KEYINPUT53), .B1(new_n699), .B2(G106gat), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n697), .A2(new_n698), .A3(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n666), .A2(new_n372), .A3(new_n667), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(G106gat), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(new_n696), .ZN(new_n704));
  AOI21_X1  g503(.A(KEYINPUT111), .B1(new_n704), .B2(KEYINPUT53), .ZN(new_n705));
  AOI22_X1  g504(.A1(new_n702), .A2(G106gat), .B1(new_n680), .B2(new_n695), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT111), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT53), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n706), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n701), .B1(new_n705), .B2(new_n709), .ZN(G1339gat));
  INV_X1    g509(.A(KEYINPUT113), .ZN(new_n711));
  AOI211_X1 g510(.A(KEYINPUT54), .B(new_n571), .C1(new_n574), .C2(new_n575), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n711), .B1(new_n712), .B2(new_n584), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT54), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n576), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n715), .A2(KEYINPUT113), .A3(new_n583), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT55), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n576), .A2(new_n714), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n587), .A2(new_n571), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n718), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n717), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n590), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n719), .A2(new_n720), .ZN(new_n724));
  AOI21_X1  g523(.A(KEYINPUT55), .B1(new_n717), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(KEYINPUT114), .B1(new_n723), .B2(new_n725), .ZN(new_n726));
  AOI22_X1  g525(.A1(new_n717), .A2(new_n721), .B1(new_n585), .B2(new_n589), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT114), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n717), .A2(new_n724), .ZN(new_n729));
  OAI211_X1 g528(.A(new_n727), .B(new_n728), .C1(new_n729), .C2(KEYINPUT55), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n726), .A2(new_n730), .A3(new_n488), .A4(new_n489), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n472), .A2(new_n464), .A3(new_n469), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n732), .B1(new_n479), .B2(new_n465), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n413), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n487), .A2(new_n592), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n731), .A2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT116), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n731), .A2(KEYINPUT116), .A3(new_n735), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n738), .A2(new_n568), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n487), .A2(new_n734), .ZN(new_n741));
  XOR2_X1   g540(.A(new_n741), .B(KEYINPUT115), .Z(new_n742));
  AND2_X1   g541(.A1(new_n726), .A2(new_n730), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n742), .A2(new_n617), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n740), .A2(new_n744), .ZN(new_n745));
  AOI22_X1  g544(.A1(new_n745), .A2(new_n526), .B1(new_n490), .B2(new_n593), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n746), .A2(new_n372), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n595), .A2(new_n404), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n748), .A2(new_n632), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(new_n494), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n750), .A2(new_n222), .A3(new_n751), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n746), .A2(new_n402), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n403), .A2(new_n404), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n643), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n752), .B1(new_n222), .B2(new_n757), .ZN(G1340gat));
  OAI21_X1  g557(.A(G120gat), .B1(new_n750), .B2(new_n611), .ZN(new_n759));
  OR2_X1    g558(.A1(new_n611), .A2(new_n220), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n759), .B1(new_n755), .B2(new_n760), .ZN(G1341gat));
  AOI21_X1  g560(.A(new_n226), .B1(new_n756), .B2(new_n527), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n747), .A2(new_n226), .A3(new_n527), .A4(new_n749), .ZN(new_n763));
  AND2_X1   g562(.A1(new_n763), .A2(KEYINPUT117), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n763), .A2(KEYINPUT117), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n762), .A2(new_n764), .A3(new_n765), .ZN(G1342gat));
  OR3_X1    g565(.A1(new_n755), .A2(G134gat), .A3(new_n568), .ZN(new_n767));
  OR2_X1    g566(.A1(new_n767), .A2(KEYINPUT56), .ZN(new_n768));
  OAI21_X1  g567(.A(G134gat), .B1(new_n750), .B2(new_n568), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n767), .A2(KEYINPUT56), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n768), .A2(new_n769), .A3(new_n770), .ZN(G1343gat));
  AND3_X1   g570(.A1(new_n731), .A2(KEYINPUT116), .A3(new_n735), .ZN(new_n772));
  AOI21_X1  g571(.A(KEYINPUT116), .B1(new_n731), .B2(new_n735), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n772), .A2(new_n773), .A3(new_n617), .ZN(new_n774));
  INV_X1    g573(.A(new_n744), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n526), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n593), .A2(new_n490), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n373), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  OAI21_X1  g577(.A(KEYINPUT118), .B1(new_n778), .B2(KEYINPUT57), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n723), .A2(new_n725), .ZN(new_n780));
  AND3_X1   g579(.A1(new_n488), .A2(KEYINPUT94), .A3(new_n489), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT94), .B1(new_n488), .B2(new_n489), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n780), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n735), .B(KEYINPUT119), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n617), .B1(new_n783), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n526), .B1(new_n786), .B2(new_n775), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT120), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OAI211_X1 g588(.A(KEYINPUT120), .B(new_n526), .C1(new_n786), .C2(new_n775), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n789), .A2(new_n777), .A3(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT57), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n373), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT118), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n795), .B(new_n792), .C1(new_n746), .C2(new_n373), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n779), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n748), .A2(new_n605), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n797), .A2(new_n494), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(G141gat), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n753), .A2(new_n269), .A3(new_n372), .A4(new_n404), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n751), .A2(G141gat), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT58), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n800), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n797), .A2(new_n643), .A3(new_n798), .ZN(new_n806));
  AOI22_X1  g605(.A1(new_n806), .A2(G141gat), .B1(new_n802), .B2(new_n803), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT58), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n805), .B1(new_n807), .B2(new_n808), .ZN(G1344gat));
  NAND3_X1  g608(.A1(new_n802), .A2(new_n312), .A3(new_n592), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT59), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(G148gat), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n797), .A2(new_n798), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n812), .B1(new_n813), .B2(new_n592), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT122), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n617), .A2(KEYINPUT121), .A3(new_n780), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n780), .A2(new_n567), .A3(new_n565), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT121), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  AND3_X1   g618(.A1(new_n742), .A2(new_n816), .A3(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n815), .B1(new_n786), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n742), .A2(new_n816), .A3(new_n819), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n784), .B1(new_n494), .B2(new_n780), .ZN(new_n823));
  OAI211_X1 g622(.A(KEYINPUT122), .B(new_n822), .C1(new_n823), .C2(new_n617), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n821), .A2(new_n824), .A3(new_n526), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n593), .A2(new_n751), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n373), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n372), .A2(KEYINPUT57), .ZN(new_n828));
  OAI22_X1  g627(.A1(new_n827), .A2(KEYINPUT57), .B1(new_n746), .B2(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n829), .A2(new_n592), .A3(new_n798), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n811), .B1(new_n830), .B2(G148gat), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n810), .B1(new_n814), .B2(new_n831), .ZN(G1345gat));
  NAND3_X1  g631(.A1(new_n802), .A2(new_n299), .A3(new_n527), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n813), .A2(new_n527), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n833), .B1(new_n834), .B2(new_n299), .ZN(G1346gat));
  NAND3_X1  g634(.A1(new_n802), .A2(new_n300), .A3(new_n617), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n813), .A2(new_n617), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n836), .B1(new_n837), .B2(new_n300), .ZN(G1347gat));
  NOR2_X1   g637(.A1(new_n746), .A2(new_n595), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n403), .A2(new_n298), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT123), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n839), .A2(KEYINPUT123), .A3(new_n840), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n490), .A2(G169gat), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT124), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n846), .B(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n595), .A2(new_n404), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n850), .A2(new_n632), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n747), .A2(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(G169gat), .B1(new_n852), .B2(new_n751), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n848), .A2(new_n853), .ZN(G1348gat));
  AND2_X1   g653(.A1(new_n843), .A2(new_n844), .ZN(new_n855));
  INV_X1    g654(.A(G176gat), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n855), .A2(new_n856), .A3(new_n592), .ZN(new_n857));
  OAI21_X1  g656(.A(G176gat), .B1(new_n852), .B2(new_n611), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(G1349gat));
  OAI21_X1  g658(.A(G183gat), .B1(new_n852), .B2(new_n526), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n527), .A2(new_n213), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n860), .B1(new_n841), .B2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT60), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n863), .A2(KEYINPUT125), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n862), .B(new_n864), .ZN(G1350gat));
  NAND3_X1  g664(.A1(new_n855), .A2(new_n214), .A3(new_n617), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n214), .B1(KEYINPUT126), .B2(KEYINPUT61), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(new_n852), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n868), .B1(new_n869), .B2(new_n617), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT126), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT61), .ZN(new_n872));
  AND3_X1   g671(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n866), .B1(new_n873), .B2(new_n874), .ZN(G1351gat));
  NOR3_X1   g674(.A1(new_n605), .A2(new_n373), .A3(new_n404), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n839), .A2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(G197gat), .B1(new_n878), .B2(new_n643), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n850), .A2(new_n605), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n829), .A2(new_n880), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n494), .A2(G197gat), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n879), .B1(new_n881), .B2(new_n882), .ZN(G1352gat));
  NAND2_X1  g682(.A1(new_n881), .A2(new_n592), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(G204gat), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n877), .A2(G204gat), .A3(new_n611), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n886), .B(KEYINPUT62), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n885), .A2(new_n887), .ZN(G1353gat));
  NAND3_X1  g687(.A1(new_n878), .A2(new_n275), .A3(new_n527), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n829), .A2(new_n527), .A3(new_n880), .ZN(new_n890));
  AND3_X1   g689(.A1(new_n890), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n891));
  AOI21_X1  g690(.A(KEYINPUT63), .B1(new_n890), .B2(G211gat), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n889), .B1(new_n891), .B2(new_n892), .ZN(G1354gat));
  NAND2_X1  g692(.A1(new_n825), .A2(new_n826), .ZN(new_n894));
  AOI21_X1  g693(.A(KEYINPUT57), .B1(new_n894), .B2(new_n372), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n746), .A2(new_n792), .A3(new_n373), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n617), .B(new_n880), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(G218gat), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n878), .A2(new_n276), .A3(new_n617), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(KEYINPUT127), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT127), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n898), .A2(new_n902), .A3(new_n899), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n901), .A2(new_n903), .ZN(G1355gat));
endmodule


