//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 1 1 0 1 0 0 0 0 0 0 1 1 0 0 1 0 1 1 0 1 1 0 1 0 0 1 0 0 1 0 1 0 0 1 0 1 0 1 0 0 1 0 0 0 1 1 1 1 1 0 1 0 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:24 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT0), .Z(new_n212));
  AOI22_X1  g0012(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n213));
  INV_X1    g0013(.A(G68), .ZN(new_n214));
  INV_X1    g0014(.A(G238), .ZN(new_n215));
  INV_X1    g0015(.A(G264), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n203), .C2(new_n216), .ZN(new_n217));
  AOI21_X1  g0017(.A(new_n217), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G50), .ZN(new_n219));
  INV_X1    g0019(.A(G226), .ZN(new_n220));
  INV_X1    g0020(.A(G77), .ZN(new_n221));
  INV_X1    g0021(.A(G244), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G58), .ZN(new_n224));
  INV_X1    g0024(.A(G232), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n209), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT1), .ZN(new_n228));
  NAND3_X1  g0028(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(KEYINPUT64), .B1(G1), .B2(G13), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n232), .A2(new_n207), .ZN(new_n233));
  NOR2_X1   g0033(.A1(G58), .A2(G68), .ZN(new_n234));
  OR2_X1    g0034(.A1(new_n234), .A2(KEYINPUT65), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n234), .A2(KEYINPUT65), .ZN(new_n236));
  NAND3_X1  g0036(.A1(new_n235), .A2(G50), .A3(new_n236), .ZN(new_n237));
  INV_X1    g0037(.A(new_n237), .ZN(new_n238));
  AOI211_X1 g0038(.A(new_n212), .B(new_n228), .C1(new_n233), .C2(new_n238), .ZN(G361));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G226), .B(G232), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G250), .B(G257), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G264), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(G270), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G358));
  XNOR2_X1  g0048(.A(G87), .B(G97), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(G107), .ZN(new_n250));
  INV_X1    g0050(.A(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(G68), .B(G77), .Z(new_n253));
  XOR2_X1   g0053(.A(G50), .B(G58), .Z(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n252), .B(new_n256), .ZN(G351));
  OR2_X1    g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G1698), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G222), .ZN(new_n262));
  INV_X1    g0062(.A(G223), .ZN(new_n263));
  OAI211_X1 g0063(.A(new_n260), .B(new_n262), .C1(new_n263), .C2(new_n261), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G1), .A2(G13), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT64), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI22_X1  g0067(.A1(new_n267), .A2(new_n229), .B1(G33), .B2(G41), .ZN(new_n268));
  OAI211_X1 g0068(.A(new_n264), .B(new_n268), .C1(G77), .C2(new_n260), .ZN(new_n269));
  AND2_X1   g0069(.A1(KEYINPUT67), .A2(G45), .ZN(new_n270));
  NOR2_X1   g0070(.A1(KEYINPUT67), .A2(G45), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OAI211_X1 g0072(.A(new_n206), .B(G274), .C1(new_n272), .C2(G41), .ZN(new_n273));
  INV_X1    g0073(.A(G33), .ZN(new_n274));
  INV_X1    g0074(.A(G41), .ZN(new_n275));
  OAI211_X1 g0075(.A(G1), .B(G13), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  OAI211_X1 g0078(.A(new_n269), .B(new_n273), .C1(new_n220), .C2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G200), .ZN(new_n280));
  INV_X1    g0080(.A(G190), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT9), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n234), .A2(new_n219), .ZN(new_n283));
  NOR2_X1   g0083(.A1(G20), .A2(G33), .ZN(new_n284));
  AOI22_X1  g0084(.A1(new_n283), .A2(G20), .B1(G150), .B2(new_n284), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT8), .B(G58), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n207), .A2(G33), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n267), .A2(new_n229), .A3(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n207), .A2(G1), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n288), .A2(new_n290), .B1(new_n292), .B2(G50), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n291), .A2(G13), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n293), .B1(G50), .B2(new_n294), .ZN(new_n295));
  OAI221_X1 g0095(.A(new_n280), .B1(new_n281), .B2(new_n279), .C1(new_n282), .C2(new_n295), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n295), .A2(new_n282), .ZN(new_n297));
  OR3_X1    g0097(.A1(new_n296), .A2(KEYINPUT10), .A3(new_n297), .ZN(new_n298));
  OAI21_X1  g0098(.A(KEYINPUT10), .B1(new_n296), .B2(new_n297), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT68), .ZN(new_n301));
  XNOR2_X1  g0101(.A(new_n273), .B(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n278), .A2(new_n215), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n225), .A2(G1698), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n304), .B1(G226), .B2(G1698), .ZN(new_n305));
  AND2_X1   g0105(.A1(KEYINPUT3), .A2(G33), .ZN(new_n306));
  NOR2_X1   g0106(.A1(KEYINPUT3), .A2(G33), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  OAI22_X1  g0108(.A1(new_n305), .A2(new_n308), .B1(new_n274), .B2(new_n202), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n303), .B1(new_n268), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n302), .A2(new_n310), .ZN(new_n311));
  XOR2_X1   g0111(.A(new_n311), .B(KEYINPUT13), .Z(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(G190), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n284), .A2(G50), .ZN(new_n314));
  OAI221_X1 g0114(.A(new_n314), .B1(new_n207), .B2(G68), .C1(new_n221), .C2(new_n287), .ZN(new_n315));
  AND2_X1   g0115(.A1(new_n315), .A2(new_n290), .ZN(new_n316));
  OR2_X1    g0116(.A1(new_n316), .A2(KEYINPUT11), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(KEYINPUT11), .ZN(new_n318));
  INV_X1    g0118(.A(new_n294), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(new_n214), .ZN(new_n320));
  XNOR2_X1  g0120(.A(new_n320), .B(KEYINPUT12), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n292), .A2(G68), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n317), .A2(new_n318), .A3(new_n321), .A4(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  XNOR2_X1  g0124(.A(new_n311), .B(KEYINPUT13), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(G200), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n313), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G169), .ZN(new_n329));
  OAI21_X1  g0129(.A(KEYINPUT14), .B1(new_n312), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n312), .A2(G179), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT14), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n325), .A2(new_n332), .A3(G169), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n330), .A2(new_n331), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n328), .B1(new_n323), .B2(new_n334), .ZN(new_n335));
  OR2_X1    g0135(.A1(new_n279), .A2(G179), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n279), .A2(new_n329), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n336), .A2(new_n295), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n261), .A2(G232), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n260), .B(new_n339), .C1(new_n215), .C2(new_n261), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n340), .B(new_n268), .C1(G107), .C2(new_n260), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n341), .B(new_n273), .C1(new_n222), .C2(new_n278), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n329), .ZN(new_n343));
  INV_X1    g0143(.A(new_n286), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n344), .A2(new_n284), .B1(G20), .B2(G77), .ZN(new_n345));
  OR2_X1    g0145(.A1(KEYINPUT15), .A2(G87), .ZN(new_n346));
  NAND2_X1  g0146(.A1(KEYINPUT15), .A2(G87), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n345), .B1(new_n287), .B2(new_n348), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n349), .A2(new_n290), .B1(G77), .B2(new_n292), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n319), .A2(new_n221), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n343), .B(new_n352), .C1(G179), .C2(new_n342), .ZN(new_n353));
  AND4_X1   g0153(.A1(new_n300), .A2(new_n335), .A3(new_n338), .A4(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT16), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n258), .A2(new_n207), .A3(new_n259), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT7), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n258), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n259), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n214), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n224), .A2(new_n214), .ZN(new_n361));
  OAI21_X1  g0161(.A(G20), .B1(new_n361), .B2(new_n234), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n284), .A2(G159), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n355), .B1(new_n360), .B2(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(KEYINPUT7), .B1(new_n308), .B2(new_n207), .ZN(new_n366));
  NOR4_X1   g0166(.A1(new_n306), .A2(new_n307), .A3(new_n357), .A4(G20), .ZN(new_n367));
  OAI21_X1  g0167(.A(G68), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n364), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n368), .A2(KEYINPUT16), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n365), .A2(new_n370), .A3(new_n290), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n344), .B1(new_n290), .B2(new_n291), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n294), .A2(new_n286), .ZN(new_n373));
  AND3_X1   g0173(.A1(new_n372), .A2(KEYINPUT69), .A3(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(KEYINPUT69), .B1(new_n372), .B2(new_n373), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n371), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n276), .A2(G232), .A3(new_n277), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n273), .A2(new_n378), .ZN(new_n379));
  OAI22_X1  g0179(.A1(new_n230), .A2(new_n231), .B1(new_n274), .B2(new_n275), .ZN(new_n380));
  NAND2_X1  g0180(.A1(G33), .A2(G87), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n263), .A2(new_n261), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n220), .A2(G1698), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n382), .B(new_n383), .C1(new_n306), .C2(new_n307), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n380), .B1(new_n381), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(G169), .B1(new_n379), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n384), .A2(new_n381), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n268), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n388), .A2(G179), .A3(new_n378), .A4(new_n273), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n377), .A2(KEYINPUT18), .A3(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(KEYINPUT18), .B1(new_n377), .B2(new_n390), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(G200), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(new_n379), .B2(new_n385), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n388), .A2(new_n281), .A3(new_n378), .A4(new_n273), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n371), .A2(new_n398), .A3(new_n376), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT17), .ZN(new_n400));
  XNOR2_X1  g0200(.A(new_n399), .B(new_n400), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n350), .B(new_n351), .C1(new_n342), .C2(new_n281), .ZN(new_n402));
  AND2_X1   g0202(.A1(new_n342), .A2(G200), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NOR3_X1   g0204(.A1(new_n394), .A2(new_n401), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n354), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n261), .A2(G257), .ZN(new_n408));
  OAI221_X1 g0208(.A(new_n408), .B1(new_n216), .B2(new_n261), .C1(new_n306), .C2(new_n307), .ZN(new_n409));
  INV_X1    g0209(.A(G303), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n308), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n409), .A2(new_n411), .A3(new_n268), .ZN(new_n412));
  INV_X1    g0212(.A(G45), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n413), .A2(G1), .ZN(new_n414));
  AND2_X1   g0214(.A1(KEYINPUT5), .A2(G41), .ZN(new_n415));
  NOR2_X1   g0215(.A1(KEYINPUT5), .A2(G41), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n414), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n417), .A2(G270), .A3(new_n276), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n414), .B(G274), .C1(new_n416), .C2(new_n415), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n412), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n420), .A2(KEYINPUT21), .A3(G169), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n412), .A2(G179), .A3(new_n418), .A4(new_n419), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n290), .B1(new_n206), .B2(G33), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n424), .A2(KEYINPUT74), .A3(G116), .A4(new_n294), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT74), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n206), .A2(G33), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n232), .A2(new_n294), .A3(new_n289), .A4(new_n427), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n426), .B1(new_n428), .B2(new_n251), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n425), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n251), .A2(G20), .ZN(new_n431));
  NAND2_X1  g0231(.A1(G33), .A2(G283), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n432), .B(new_n207), .C1(G33), .C2(new_n202), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n290), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT20), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n290), .A2(KEYINPUT20), .A3(new_n431), .A4(new_n433), .ZN(new_n437));
  AOI22_X1  g0237(.A1(new_n436), .A2(new_n437), .B1(new_n251), .B2(new_n319), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n430), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n423), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n420), .A2(G169), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n441), .B1(new_n438), .B2(new_n430), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n440), .B1(KEYINPUT21), .B2(new_n442), .ZN(new_n443));
  OR2_X1    g0243(.A1(G250), .A2(G1698), .ZN(new_n444));
  OAI221_X1 g0244(.A(new_n444), .B1(G257), .B2(new_n261), .C1(new_n306), .C2(new_n307), .ZN(new_n445));
  NAND2_X1  g0245(.A1(G33), .A2(G294), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n268), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n417), .A2(G264), .A3(new_n276), .ZN(new_n449));
  INV_X1    g0249(.A(G179), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n448), .A2(new_n449), .A3(new_n450), .A4(new_n419), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n380), .B1(new_n445), .B2(new_n446), .ZN(new_n452));
  INV_X1    g0252(.A(new_n449), .ZN(new_n453));
  INV_X1    g0253(.A(new_n419), .ZN(new_n454));
  NOR3_X1   g0254(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n451), .B1(new_n455), .B2(G169), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n207), .B(G87), .C1(new_n306), .C2(new_n307), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(KEYINPUT22), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT22), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n260), .A2(new_n459), .A3(new_n207), .A4(G87), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT24), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT23), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n463), .B1(new_n207), .B2(G107), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n203), .A2(KEYINPUT23), .A3(G20), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n274), .A2(new_n251), .ZN(new_n466));
  AOI22_X1  g0266(.A1(new_n464), .A2(new_n465), .B1(new_n466), .B2(new_n207), .ZN(new_n467));
  AND3_X1   g0267(.A1(new_n461), .A2(new_n462), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n462), .B1(new_n461), .B2(new_n467), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n290), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n428), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT25), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n472), .B1(new_n294), .B2(G107), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n319), .A2(KEYINPUT25), .A3(new_n203), .ZN(new_n474));
  AOI22_X1  g0274(.A1(new_n471), .A2(G107), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n456), .B1(new_n470), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n443), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n206), .A2(G45), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n276), .A2(G250), .A3(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT71), .ZN(new_n480));
  INV_X1    g0280(.A(G274), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n480), .B1(new_n478), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n414), .A2(KEYINPUT71), .A3(G274), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NOR2_X1   g0284(.A1(G238), .A2(G1698), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n485), .B1(new_n258), .B2(new_n259), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n222), .A2(G1698), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n466), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n479), .B(new_n484), .C1(new_n488), .C2(new_n380), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(G200), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n215), .A2(new_n261), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n491), .B(new_n487), .C1(new_n306), .C2(new_n307), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n268), .B1(new_n493), .B2(new_n466), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n494), .A2(G190), .A3(new_n479), .A4(new_n484), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT19), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n496), .B1(new_n287), .B2(new_n202), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n207), .B(G68), .C1(new_n306), .C2(new_n307), .ZN(new_n498));
  INV_X1    g0298(.A(G87), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(KEYINPUT72), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT72), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(G87), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n204), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n504));
  AND2_X1   g0304(.A1(new_n504), .A2(new_n207), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n497), .B(new_n498), .C1(new_n503), .C2(new_n505), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n506), .A2(new_n290), .B1(new_n319), .B2(new_n348), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n471), .A2(G87), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n490), .A2(new_n495), .A3(new_n507), .A4(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n348), .A2(KEYINPUT73), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT73), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n346), .A2(new_n511), .A3(new_n347), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n424), .A2(new_n513), .A3(new_n294), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n506), .A2(new_n290), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n319), .A2(new_n348), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n489), .A2(new_n329), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n494), .A2(new_n450), .A3(new_n479), .A4(new_n484), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  AND2_X1   g0320(.A1(new_n509), .A2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT4), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n522), .A2(G1698), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n523), .B(G244), .C1(new_n307), .C2(new_n306), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n222), .B1(new_n258), .B2(new_n259), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n524), .B(new_n432), .C1(new_n525), .C2(KEYINPUT4), .ZN(new_n526));
  OAI21_X1  g0326(.A(G250), .B1(new_n306), .B2(new_n307), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n261), .B1(new_n527), .B2(KEYINPUT4), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n268), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n417), .A2(G257), .A3(new_n276), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n419), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n529), .A2(G179), .A3(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(G244), .B1(new_n306), .B2(new_n307), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n534), .A2(new_n522), .B1(G33), .B2(G283), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n522), .B1(new_n260), .B2(G250), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n535), .B(new_n524), .C1(new_n261), .C2(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n531), .B1(new_n537), .B2(new_n268), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n533), .B1(new_n538), .B2(new_n329), .ZN(new_n539));
  OAI21_X1  g0339(.A(G107), .B1(new_n366), .B2(new_n367), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT70), .ZN(new_n541));
  NAND2_X1  g0341(.A1(KEYINPUT6), .A2(G97), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n541), .B1(new_n542), .B2(G107), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n203), .A2(KEYINPUT70), .A3(KEYINPUT6), .A4(G97), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(G97), .A2(G107), .ZN(new_n546));
  AOI21_X1  g0346(.A(KEYINPUT6), .B1(new_n204), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g0347(.A(G20), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n284), .A2(G77), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n540), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n290), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n319), .A2(new_n202), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n471), .A2(G97), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n539), .A2(new_n554), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n550), .A2(new_n290), .B1(new_n471), .B2(G97), .ZN(new_n556));
  AND3_X1   g0356(.A1(new_n529), .A2(new_n281), .A3(new_n532), .ZN(new_n557));
  AOI21_X1  g0357(.A(G200), .B1(new_n529), .B2(new_n532), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n556), .B(new_n552), .C1(new_n557), .C2(new_n558), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n448), .A2(new_n449), .A3(new_n281), .A4(new_n419), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n560), .B1(new_n455), .B2(G200), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n561), .A2(new_n470), .A3(new_n475), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n521), .A2(new_n555), .A3(new_n559), .A4(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n439), .B1(G200), .B2(new_n420), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(new_n281), .B2(new_n420), .ZN(new_n566));
  AND4_X1   g0366(.A1(new_n407), .A2(new_n477), .A3(new_n564), .A4(new_n566), .ZN(G372));
  INV_X1    g0367(.A(KEYINPUT77), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n300), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n298), .A2(new_n299), .A3(KEYINPUT77), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n334), .A2(new_n323), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n328), .B1(new_n572), .B2(new_n353), .ZN(new_n573));
  XNOR2_X1  g0373(.A(new_n399), .B(KEYINPUT17), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n571), .B1(new_n575), .B2(new_n394), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n338), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n470), .A2(new_n475), .ZN(new_n579));
  INV_X1    g0379(.A(new_n455), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n329), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n579), .A2(new_n581), .A3(new_n451), .ZN(new_n582));
  OR2_X1    g0382(.A1(new_n442), .A2(KEYINPUT21), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n582), .A2(new_n583), .A3(new_n440), .ZN(new_n584));
  AND2_X1   g0384(.A1(new_n521), .A2(new_n562), .ZN(new_n585));
  AND2_X1   g0385(.A1(new_n555), .A2(new_n559), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n555), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n521), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(KEYINPUT26), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT76), .ZN(new_n591));
  AND3_X1   g0391(.A1(new_n529), .A2(G179), .A3(new_n532), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n329), .B1(new_n529), .B2(new_n532), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n533), .B(KEYINPUT76), .C1(new_n538), .C2(new_n329), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT26), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n596), .A2(new_n597), .A3(new_n521), .A4(new_n554), .ZN(new_n598));
  XOR2_X1   g0398(.A(new_n520), .B(KEYINPUT75), .Z(new_n599));
  NAND4_X1  g0399(.A1(new_n587), .A2(new_n590), .A3(new_n598), .A4(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n578), .B1(new_n406), .B2(new_n601), .ZN(G369));
  INV_X1    g0402(.A(G13), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n603), .A2(G20), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n206), .ZN(new_n605));
  OR2_X1    g0405(.A1(new_n605), .A2(KEYINPUT27), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(KEYINPUT27), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n606), .A2(G213), .A3(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(G343), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n579), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n476), .B1(new_n611), .B2(new_n562), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n582), .A2(new_n610), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT78), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g0416(.A(KEYINPUT78), .B1(new_n612), .B2(new_n613), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n443), .ZN(new_n620));
  INV_X1    g0420(.A(new_n610), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n621), .B1(new_n438), .B2(new_n430), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n622), .B1(new_n620), .B2(new_n566), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(G330), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n619), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n443), .A2(new_n621), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n629), .B1(new_n616), .B2(new_n617), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n630), .A2(new_n613), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n628), .A2(new_n631), .ZN(G399));
  INV_X1    g0432(.A(new_n210), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n633), .A2(G41), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n503), .A2(new_n251), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n635), .A2(G1), .A3(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n638), .B1(new_n237), .B2(new_n635), .ZN(new_n639));
  XNOR2_X1  g0439(.A(new_n639), .B(KEYINPUT28), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n587), .A2(new_n599), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n589), .A2(KEYINPUT26), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n594), .A2(new_n595), .B1(new_n552), .B2(new_n556), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n597), .B1(new_n643), .B2(new_n521), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n610), .B1(new_n641), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(KEYINPUT29), .ZN(new_n647));
  XOR2_X1   g0447(.A(new_n647), .B(KEYINPUT82), .Z(new_n648));
  NAND2_X1  g0448(.A1(new_n600), .A2(new_n621), .ZN(new_n649));
  XNOR2_X1  g0449(.A(new_n649), .B(KEYINPUT79), .ZN(new_n650));
  XOR2_X1   g0450(.A(KEYINPUT80), .B(KEYINPUT29), .Z(new_n651));
  NAND3_X1  g0451(.A1(new_n650), .A2(KEYINPUT81), .A3(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(KEYINPUT81), .B1(new_n650), .B2(new_n651), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n648), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n564), .A2(new_n477), .A3(new_n566), .A4(new_n621), .ZN(new_n656));
  INV_X1    g0456(.A(new_n420), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n592), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT30), .ZN(new_n659));
  OR3_X1    g0459(.A1(new_n489), .A2(new_n452), .A3(new_n453), .ZN(new_n660));
  OR3_X1    g0460(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n659), .B1(new_n658), .B2(new_n660), .ZN(new_n662));
  INV_X1    g0462(.A(new_n538), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n657), .A2(G179), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n663), .A2(new_n664), .A3(new_n580), .A4(new_n489), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n661), .A2(new_n662), .A3(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n666), .A2(KEYINPUT31), .A3(new_n610), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n656), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(KEYINPUT31), .B1(new_n666), .B2(new_n610), .ZN(new_n669));
  OAI21_X1  g0469(.A(G330), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n655), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n640), .B1(new_n672), .B2(G1), .ZN(G364));
  INV_X1    g0473(.A(new_n625), .ZN(new_n674));
  INV_X1    g0474(.A(G330), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n604), .A2(G45), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n635), .A2(G1), .A3(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n676), .A2(new_n626), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g0479(.A(new_n679), .B(KEYINPUT83), .ZN(new_n680));
  NOR2_X1   g0480(.A1(G13), .A2(G33), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(G20), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n678), .B1(new_n674), .B2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n210), .A2(G355), .A3(new_n260), .ZN(new_n685));
  OAI22_X1  g0485(.A1(new_n256), .A2(new_n413), .B1(new_n237), .B2(new_n272), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n633), .A2(new_n260), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  OAI221_X1 g0488(.A(new_n685), .B1(G116), .B2(new_n210), .C1(new_n686), .C2(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n232), .B1(G20), .B2(new_n329), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(new_n683), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n207), .A2(new_n450), .ZN(new_n693));
  XOR2_X1   g0493(.A(new_n693), .B(KEYINPUT84), .Z(new_n694));
  AND3_X1   g0494(.A1(new_n694), .A2(G190), .A3(new_n395), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(G322), .ZN(new_n696));
  NOR2_X1   g0496(.A1(G179), .A2(G200), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT85), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n698), .A2(G190), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(new_n207), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(new_n698), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n207), .A2(G179), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n703), .A2(new_n281), .A3(G200), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  AOI22_X1  g0505(.A1(new_n702), .A2(G329), .B1(G283), .B2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n700), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(G294), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n693), .A2(G200), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(G190), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(G317), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n712), .A2(KEYINPUT33), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n712), .A2(KEYINPUT33), .ZN(new_n714));
  NOR3_X1   g0514(.A1(new_n711), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n709), .A2(new_n281), .ZN(new_n716));
  XOR2_X1   g0516(.A(KEYINPUT87), .B(G326), .Z(new_n717));
  AOI211_X1 g0517(.A(new_n260), .B(new_n715), .C1(new_n716), .C2(new_n717), .ZN(new_n718));
  AND4_X1   g0518(.A1(new_n696), .A2(new_n706), .A3(new_n708), .A4(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n703), .A2(G190), .A3(G200), .ZN(new_n720));
  INV_X1    g0520(.A(G311), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n694), .A2(new_n281), .A3(new_n395), .ZN(new_n722));
  OAI221_X1 g0522(.A(new_n719), .B1(new_n410), .B2(new_n720), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(G159), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n701), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n725), .B(KEYINPUT32), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n707), .A2(G97), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n500), .A2(new_n502), .ZN(new_n728));
  OAI221_X1 g0528(.A(new_n260), .B1(new_n704), .B2(new_n203), .C1(new_n728), .C2(new_n720), .ZN(new_n729));
  XOR2_X1   g0529(.A(new_n729), .B(KEYINPUT86), .Z(new_n730));
  AOI22_X1  g0530(.A1(new_n710), .A2(G68), .B1(new_n716), .B2(G50), .ZN(new_n731));
  INV_X1    g0531(.A(new_n695), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n731), .B1(new_n732), .B2(new_n224), .ZN(new_n733));
  INV_X1    g0533(.A(new_n722), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n733), .B1(G77), .B2(new_n734), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n726), .A2(new_n727), .A3(new_n730), .A4(new_n735), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n723), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n690), .ZN(new_n738));
  OAI211_X1 g0538(.A(new_n684), .B(new_n692), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n680), .A2(new_n739), .ZN(G396));
  NOR2_X1   g0540(.A1(new_n353), .A2(new_n610), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n352), .A2(new_n610), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n742), .B1(new_n402), .B2(new_n403), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n741), .B1(new_n743), .B2(new_n353), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT89), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n600), .A2(new_n746), .A3(new_n621), .A4(new_n744), .ZN(new_n747));
  OAI211_X1 g0547(.A(new_n598), .B(new_n599), .C1(new_n477), .C2(new_n563), .ZN(new_n748));
  INV_X1    g0548(.A(new_n590), .ZN(new_n749));
  OAI211_X1 g0549(.A(new_n621), .B(new_n744), .C1(new_n748), .C2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(KEYINPUT89), .ZN(new_n751));
  AOI22_X1  g0551(.A1(new_n650), .A2(new_n745), .B1(new_n747), .B2(new_n751), .ZN(new_n752));
  XOR2_X1   g0552(.A(new_n752), .B(new_n670), .Z(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(new_n678), .ZN(new_n754));
  INV_X1    g0554(.A(new_n678), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n308), .B1(new_n701), .B2(new_n721), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n705), .A2(G87), .ZN(new_n757));
  INV_X1    g0557(.A(new_n716), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n757), .B1(new_n758), .B2(new_n410), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n759), .B1(new_n707), .B2(G97), .ZN(new_n760));
  INV_X1    g0560(.A(G294), .ZN(new_n761));
  OAI221_X1 g0561(.A(new_n760), .B1(new_n203), .B2(new_n720), .C1(new_n761), .C2(new_n732), .ZN(new_n762));
  AOI211_X1 g0562(.A(new_n756), .B(new_n762), .C1(G116), .C2(new_n734), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n710), .A2(G283), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n260), .B1(new_n700), .B2(new_n224), .ZN(new_n765));
  INV_X1    g0565(.A(G132), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n701), .A2(new_n766), .B1(new_n219), .B2(new_n720), .ZN(new_n767));
  AOI211_X1 g0567(.A(new_n765), .B(new_n767), .C1(G68), .C2(new_n705), .ZN(new_n768));
  AOI22_X1  g0568(.A1(new_n695), .A2(G143), .B1(G150), .B2(new_n710), .ZN(new_n769));
  INV_X1    g0569(.A(G137), .ZN(new_n770));
  OAI221_X1 g0570(.A(new_n769), .B1(new_n770), .B2(new_n758), .C1(new_n724), .C2(new_n722), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(KEYINPUT34), .ZN(new_n772));
  AOI22_X1  g0572(.A1(new_n763), .A2(new_n764), .B1(new_n768), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n738), .A2(new_n682), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n774), .B(KEYINPUT88), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n773), .A2(new_n738), .B1(G77), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n744), .A2(new_n682), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n755), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n754), .A2(new_n778), .ZN(new_n779));
  AND2_X1   g0579(.A1(new_n779), .A2(KEYINPUT90), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n779), .A2(KEYINPUT90), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(G384));
  NOR2_X1   g0583(.A1(new_n572), .A2(new_n610), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(KEYINPUT39), .ZN(new_n786));
  INV_X1    g0586(.A(KEYINPUT37), .ZN(new_n787));
  AND3_X1   g0587(.A1(new_n371), .A2(new_n398), .A3(new_n376), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n372), .A2(new_n373), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n371), .A2(new_n789), .B1(new_n386), .B2(new_n389), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n608), .B1(new_n371), .B2(new_n789), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n787), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  XNOR2_X1  g0594(.A(new_n608), .B(KEYINPUT92), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n377), .B1(new_n390), .B2(new_n795), .ZN(new_n796));
  AND3_X1   g0596(.A1(new_n796), .A2(new_n787), .A3(new_n399), .ZN(new_n797));
  OAI21_X1  g0597(.A(KEYINPUT93), .B1(new_n794), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n792), .B1(new_n394), .B2(new_n401), .ZN(new_n799));
  INV_X1    g0599(.A(KEYINPUT93), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n796), .A2(new_n787), .A3(new_n399), .ZN(new_n801));
  NOR3_X1   g0601(.A1(new_n788), .A2(new_n790), .A3(new_n792), .ZN(new_n802));
  OAI211_X1 g0602(.A(new_n800), .B(new_n801), .C1(new_n802), .C2(new_n787), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n798), .A2(new_n799), .A3(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(KEYINPUT38), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n798), .A2(KEYINPUT38), .A3(new_n799), .A4(new_n803), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n786), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n377), .A2(new_n795), .ZN(new_n809));
  INV_X1    g0609(.A(new_n393), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(new_n391), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n809), .B1(new_n811), .B2(new_n574), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n787), .B1(new_n796), .B2(new_n399), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n797), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n805), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n807), .A2(new_n786), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(KEYINPUT94), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n808), .A2(new_n817), .ZN(new_n818));
  AOI211_X1 g0618(.A(KEYINPUT94), .B(new_n786), .C1(new_n806), .C2(new_n807), .ZN(new_n819));
  OAI21_X1  g0619(.A(KEYINPUT95), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT94), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n808), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT95), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n822), .B(new_n823), .C1(new_n808), .C2(new_n817), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n785), .B1(new_n820), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n323), .A2(new_n610), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n572), .A2(new_n327), .A3(new_n826), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n334), .A2(new_n323), .A3(new_n610), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n806), .A2(new_n807), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT91), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n751), .A2(new_n747), .ZN(new_n832));
  INV_X1    g0632(.A(new_n741), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n831), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  AOI211_X1 g0634(.A(KEYINPUT91), .B(new_n741), .C1(new_n751), .C2(new_n747), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n829), .B(new_n830), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n811), .A2(new_n795), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n825), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n840), .B(KEYINPUT96), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n647), .B(KEYINPUT82), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n650), .A2(new_n651), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT81), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n842), .B1(new_n845), .B2(new_n652), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(new_n407), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(new_n578), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n841), .B(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n745), .B1(new_n827), .B2(new_n828), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n666), .A2(KEYINPUT97), .A3(new_n610), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT31), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(KEYINPUT97), .B1(new_n666), .B2(new_n610), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n667), .B(new_n656), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n850), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT40), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n857), .A2(new_n858), .A3(new_n830), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n807), .A2(new_n815), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(KEYINPUT40), .B1(new_n856), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n863), .A2(new_n855), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(G330), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n855), .A2(G330), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n406), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n864), .A2(new_n407), .B1(new_n865), .B2(new_n868), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n849), .B(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n870), .B1(new_n206), .B2(new_n604), .ZN(new_n871));
  OR2_X1    g0671(.A1(new_n545), .A2(new_n547), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n251), .B1(new_n872), .B2(KEYINPUT35), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n873), .B(new_n233), .C1(KEYINPUT35), .C2(new_n872), .ZN(new_n874));
  XNOR2_X1  g0674(.A(new_n874), .B(KEYINPUT36), .ZN(new_n875));
  NOR3_X1   g0675(.A1(new_n237), .A2(new_n221), .A3(new_n361), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n214), .A2(G50), .ZN(new_n877));
  OAI211_X1 g0677(.A(G1), .B(new_n603), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n871), .A2(new_n875), .A3(new_n878), .ZN(G367));
  INV_X1    g0679(.A(new_n630), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n554), .A2(new_n610), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n586), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n643), .A2(new_n610), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT98), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n882), .A2(KEYINPUT98), .A3(new_n883), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n880), .A2(new_n889), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n890), .A2(KEYINPUT42), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n890), .A2(KEYINPUT42), .ZN(new_n892));
  OR2_X1    g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n507), .A2(new_n508), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n610), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n521), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n896), .B1(new_n599), .B2(new_n895), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n897), .A2(KEYINPUT43), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n555), .B1(new_n889), .B2(new_n582), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n621), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n893), .A2(KEYINPUT99), .A3(new_n898), .A4(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT99), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n900), .B1(new_n891), .B2(new_n892), .ZN(new_n903));
  INV_X1    g0703(.A(new_n898), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n902), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n897), .A2(KEYINPUT43), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n903), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n901), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT100), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n627), .A2(new_n888), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n910), .A2(new_n909), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n627), .A2(KEYINPUT100), .A3(new_n888), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n914), .B1(new_n908), .B2(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n912), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n634), .B(KEYINPUT41), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT44), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT101), .ZN(new_n921));
  OR2_X1    g0721(.A1(new_n630), .A2(new_n613), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n921), .B1(new_n922), .B2(new_n889), .ZN(new_n923));
  NOR3_X1   g0723(.A1(new_n631), .A2(KEYINPUT101), .A3(new_n888), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n920), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT45), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n922), .B2(new_n889), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n631), .A2(KEYINPUT45), .A3(new_n888), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n922), .A2(new_n921), .A3(new_n889), .ZN(new_n930));
  OAI21_X1  g0730(.A(KEYINPUT101), .B1(new_n631), .B2(new_n888), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n930), .A2(KEYINPUT44), .A3(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n925), .A2(new_n929), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n627), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT102), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT103), .B1(new_n619), .B2(new_n629), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n880), .A2(new_n626), .ZN(new_n938));
  XOR2_X1   g0738(.A(new_n937), .B(new_n938), .Z(new_n939));
  AND3_X1   g0739(.A1(new_n655), .A2(new_n670), .A3(new_n939), .ZN(new_n940));
  NAND4_X1  g0740(.A1(new_n925), .A2(new_n628), .A3(new_n929), .A4(new_n932), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n933), .A2(KEYINPUT102), .A3(new_n627), .ZN(new_n942));
  NAND4_X1  g0742(.A1(new_n936), .A2(new_n940), .A3(new_n941), .A4(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n919), .B1(new_n943), .B2(new_n672), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n677), .A2(G1), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n917), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  AND2_X1   g0746(.A1(new_n247), .A2(new_n687), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n691), .B1(new_n210), .B2(new_n348), .ZN(new_n948));
  INV_X1    g0748(.A(G283), .ZN(new_n949));
  OAI221_X1 g0749(.A(new_n308), .B1(new_n722), .B2(new_n949), .C1(new_n203), .C2(new_n700), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n720), .A2(new_n251), .ZN(new_n951));
  OAI22_X1  g0751(.A1(new_n758), .A2(new_n721), .B1(KEYINPUT46), .B2(new_n951), .ZN(new_n952));
  OAI22_X1  g0752(.A1(new_n711), .A2(new_n761), .B1(new_n202), .B2(new_n704), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n951), .A2(KEYINPUT46), .ZN(new_n954));
  NOR4_X1   g0754(.A1(new_n950), .A2(new_n952), .A3(new_n953), .A4(new_n954), .ZN(new_n955));
  OAI221_X1 g0755(.A(new_n955), .B1(new_n410), .B2(new_n732), .C1(new_n712), .C2(new_n701), .ZN(new_n956));
  INV_X1    g0756(.A(new_n720), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n734), .A2(G50), .B1(G58), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n707), .A2(G68), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n260), .B1(new_n704), .B2(new_n221), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n958), .B(new_n959), .C1(KEYINPUT104), .C2(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n961), .B1(G150), .B2(new_n695), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n716), .A2(G143), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n960), .A2(KEYINPUT104), .B1(new_n710), .B2(G159), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n701), .A2(new_n770), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n956), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n967), .B(KEYINPUT47), .Z(new_n968));
  OAI221_X1 g0768(.A(new_n755), .B1(new_n947), .B2(new_n948), .C1(new_n968), .C2(new_n738), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT105), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n969), .A2(new_n970), .ZN(new_n972));
  INV_X1    g0772(.A(new_n683), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n971), .B(new_n972), .C1(new_n973), .C2(new_n897), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n974), .B(KEYINPUT106), .Z(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n946), .A2(new_n976), .ZN(G387));
  INV_X1    g0777(.A(KEYINPUT107), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n940), .B2(new_n635), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n655), .A2(new_n670), .A3(new_n939), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n980), .A2(KEYINPUT107), .A3(new_n634), .ZN(new_n981));
  OAI211_X1 g0781(.A(new_n979), .B(new_n981), .C1(new_n672), .C2(new_n939), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n707), .A2(new_n513), .ZN(new_n983));
  INV_X1    g0783(.A(G150), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n983), .B1(new_n701), .B2(new_n984), .C1(new_n219), .C2(new_n732), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(G159), .B2(new_n716), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n734), .A2(G68), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n711), .A2(new_n286), .B1(new_n202), .B2(new_n704), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n988), .B1(G77), .B2(new_n957), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n986), .A2(new_n260), .A3(new_n987), .A4(new_n989), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n695), .A2(G317), .B1(G311), .B2(new_n710), .ZN(new_n991));
  INV_X1    g0791(.A(G322), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n991), .B1(new_n410), .B2(new_n722), .C1(new_n992), .C2(new_n758), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT48), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n994), .B1(new_n949), .B2(new_n700), .C1(new_n761), .C2(new_n720), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT49), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n702), .A2(new_n717), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n705), .A2(G116), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n997), .A2(new_n308), .A3(new_n998), .A4(new_n999), .ZN(new_n1000));
  AND2_X1   g0800(.A1(new_n995), .A2(new_n996), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n990), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n286), .A2(G50), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT50), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n636), .B1(G68), .B2(G77), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1004), .A2(new_n1005), .A3(new_n413), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n688), .B1(new_n244), .B2(new_n272), .ZN(new_n1007));
  NOR3_X1   g0807(.A1(new_n637), .A2(new_n633), .A3(new_n308), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1006), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(G107), .B2(new_n210), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n1002), .A2(new_n690), .B1(new_n691), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n755), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(new_n619), .B2(new_n683), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(new_n945), .B2(new_n939), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n982), .A2(new_n1014), .ZN(G393));
  INV_X1    g0815(.A(KEYINPUT108), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n934), .A2(new_n1016), .A3(new_n941), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n933), .A2(KEYINPUT108), .A3(new_n627), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT109), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1017), .A2(KEYINPUT109), .A3(new_n1018), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1021), .A2(new_n945), .A3(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n308), .B1(new_n720), .B2(new_n949), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n695), .A2(G311), .B1(G317), .B2(new_n716), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT52), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n1024), .B(new_n1026), .C1(G107), .C2(new_n705), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n734), .A2(G294), .B1(G303), .B2(new_n710), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n251), .B2(new_n700), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT111), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1027), .B(new_n1030), .C1(new_n992), .C2(new_n701), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT112), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n695), .A2(G159), .B1(G150), .B2(new_n716), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(KEYINPUT110), .B(KEYINPUT51), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1033), .B(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n757), .B1(new_n722), .B2(new_n286), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n700), .A2(new_n221), .B1(new_n214), .B2(new_n720), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n1036), .B(new_n1037), .C1(G50), .C2(new_n710), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n308), .B1(new_n702), .B2(G143), .ZN(new_n1039));
  AND3_X1   g0839(.A1(new_n1035), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n690), .B1(new_n1032), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n889), .A2(new_n683), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n691), .B1(new_n202), .B2(new_n210), .C1(new_n252), .C2(new_n688), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1041), .A2(new_n755), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1017), .A2(new_n980), .A3(new_n1018), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n943), .A2(new_n1045), .A3(new_n634), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1023), .A2(new_n1044), .A3(new_n1046), .ZN(G390));
  NAND2_X1  g0847(.A1(new_n743), .A2(new_n353), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n646), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n833), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT113), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1049), .A2(KEYINPUT113), .A3(new_n833), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1052), .A2(new_n829), .A3(new_n1053), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n861), .A2(new_n784), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n832), .A2(new_n833), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(KEYINPUT91), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n832), .A2(new_n831), .A3(new_n833), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n784), .B1(new_n1060), .B2(new_n829), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n820), .A2(new_n824), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1056), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT114), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n850), .A2(G330), .A3(new_n855), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1065), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1063), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n829), .A2(new_n744), .ZN(new_n1068));
  OR3_X1    g0868(.A1(new_n1068), .A2(KEYINPUT115), .A3(new_n670), .ZN(new_n1069));
  OAI21_X1  g0869(.A(KEYINPUT115), .B1(new_n1068), .B2(new_n670), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1071), .B(new_n1056), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(KEYINPUT114), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n829), .B1(new_n834), .B2(new_n835), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n785), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1075), .A2(new_n820), .A3(new_n824), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1065), .B1(new_n1076), .B2(new_n1056), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1067), .B1(new_n1073), .B2(new_n1077), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n577), .B(new_n867), .C1(new_n846), .C2(new_n407), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n829), .ZN(new_n1080));
  AND2_X1   g0880(.A1(new_n866), .A2(KEYINPUT117), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n744), .B1(new_n866), .B2(KEYINPUT117), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1080), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1071), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT116), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n670), .A2(new_n745), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1065), .B1(new_n1087), .B2(new_n829), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1060), .A2(new_n1086), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1086), .B1(new_n1060), .B2(new_n1088), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1085), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  AND2_X1   g0892(.A1(new_n1079), .A2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(KEYINPUT118), .B1(new_n1078), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1078), .A2(new_n1093), .ZN(new_n1095));
  AND2_X1   g0895(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1096));
  AND2_X1   g0896(.A1(new_n820), .A2(new_n824), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1096), .B1(new_n1097), .B2(new_n1075), .ZN(new_n1098));
  OAI211_X1 g0898(.A(KEYINPUT114), .B(new_n1072), .C1(new_n1098), .C2(new_n1065), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT118), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1079), .A2(new_n1092), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .A4(new_n1067), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1094), .A2(new_n634), .A3(new_n1095), .A4(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n702), .A2(G125), .ZN(new_n1104));
  XOR2_X1   g0904(.A(KEYINPUT54), .B(G143), .Z(new_n1105));
  AOI22_X1  g0905(.A1(new_n734), .A2(new_n1105), .B1(G128), .B2(new_n716), .ZN(new_n1106));
  AND2_X1   g0906(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  OAI221_X1 g0907(.A(new_n1107), .B1(new_n766), .B2(new_n732), .C1(new_n724), .C2(new_n700), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n704), .A2(new_n219), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n957), .A2(G150), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT53), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n260), .B1(new_n711), .B2(new_n770), .ZN(new_n1112));
  NOR4_X1   g0912(.A1(new_n1108), .A2(new_n1109), .A3(new_n1111), .A4(new_n1112), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n722), .A2(new_n202), .B1(new_n203), .B2(new_n711), .ZN(new_n1114));
  OR2_X1    g0914(.A1(new_n1114), .A2(KEYINPUT119), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n260), .B1(new_n1114), .B2(KEYINPUT119), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n707), .A2(G77), .B1(G283), .B2(new_n716), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n957), .A2(G87), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n695), .A2(G116), .B1(G68), .B2(new_n705), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1117), .A2(new_n1118), .A3(new_n1119), .A4(new_n1120), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n1116), .B(new_n1121), .C1(G294), .C2(new_n702), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n690), .B1(new_n1113), .B2(new_n1122), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n755), .B(new_n1123), .C1(new_n1062), .C2(new_n682), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n775), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1124), .B1(new_n286), .B2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1126), .B1(new_n1078), .B2(new_n945), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1103), .A2(new_n1127), .ZN(G378));
  INV_X1    g0928(.A(KEYINPUT57), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT121), .ZN(new_n1130));
  OR2_X1    g0930(.A1(new_n808), .A2(new_n817), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n823), .B1(new_n1131), .B2(new_n822), .ZN(new_n1132));
  NOR3_X1   g0932(.A1(new_n818), .A2(KEYINPUT95), .A3(new_n819), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n784), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  AND2_X1   g0934(.A1(new_n836), .A2(new_n838), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1134), .A2(new_n1135), .A3(new_n865), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n675), .B1(new_n859), .B2(new_n862), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1137), .B1(new_n825), .B2(new_n839), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT120), .ZN(new_n1139));
  AND3_X1   g0939(.A1(new_n571), .A2(new_n1139), .A3(new_n338), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1139), .B1(new_n571), .B2(new_n338), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n608), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n295), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  OR3_X1    g0944(.A1(new_n1140), .A2(new_n1141), .A3(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1144), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1147), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  AND3_X1   g0950(.A1(new_n1136), .A2(new_n1138), .A3(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1150), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1130), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1150), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1136), .A2(new_n1138), .A3(new_n1150), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1156), .A2(KEYINPUT121), .A3(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1153), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1079), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(new_n1078), .B2(new_n1093), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1129), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1156), .A2(KEYINPUT57), .A3(new_n1157), .ZN(new_n1163));
  OAI21_X1  g0963(.A(KEYINPUT122), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1164));
  NOR3_X1   g0964(.A1(new_n1151), .A2(new_n1152), .A3(new_n1129), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT122), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1101), .B1(new_n1099), .B2(new_n1067), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1165), .B(new_n1166), .C1(new_n1160), .C2(new_n1167), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1162), .A2(new_n634), .A3(new_n1164), .A4(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1153), .A2(new_n1158), .A3(new_n945), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1155), .A2(new_n681), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n260), .A2(G41), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n710), .A2(G97), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n695), .A2(G107), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n959), .A2(new_n1172), .A3(new_n1173), .A4(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(G77), .B2(new_n957), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n716), .A2(G116), .B1(new_n705), .B2(G58), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1176), .B(new_n1177), .C1(new_n949), .C2(new_n701), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(new_n513), .B2(new_n734), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1179), .B(KEYINPUT58), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n219), .B1(new_n306), .B2(G41), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n707), .A2(G150), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n695), .A2(G128), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n716), .A2(G125), .B1(new_n957), .B2(new_n1105), .ZN(new_n1184));
  AND3_X1   g0984(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n1185), .B1(new_n766), .B2(new_n711), .C1(new_n770), .C2(new_n722), .ZN(new_n1186));
  OR2_X1    g0986(.A1(new_n1186), .A2(KEYINPUT59), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n705), .A2(G159), .ZN(new_n1188));
  AOI21_X1  g0988(.A(G41), .B1(new_n702), .B2(G124), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1187), .A2(new_n274), .A3(new_n1188), .A4(new_n1189), .ZN(new_n1190));
  AND2_X1   g0990(.A1(new_n1186), .A2(KEYINPUT59), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1181), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n690), .B1(new_n1180), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1125), .A2(new_n219), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n1171), .A2(new_n755), .A3(new_n1193), .A4(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1170), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1169), .A2(new_n1197), .ZN(G375));
  NOR2_X1   g0998(.A1(new_n1079), .A2(new_n1092), .ZN(new_n1199));
  NOR3_X1   g0999(.A1(new_n1093), .A2(new_n1199), .A3(new_n919), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n1200), .B(KEYINPUT123), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n702), .A2(G303), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n260), .B1(new_n695), .B2(G283), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n734), .A2(G107), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1202), .A2(new_n983), .A3(new_n1203), .A4(new_n1204), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n711), .A2(new_n251), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n758), .A2(new_n761), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n704), .A2(new_n221), .B1(new_n720), .B2(new_n202), .ZN(new_n1208));
  NOR4_X1   g1008(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .A4(new_n1208), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n695), .A2(G137), .B1(new_n710), .B2(new_n1105), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1210), .B1(new_n219), .B2(new_n700), .C1(new_n224), .C2(new_n704), .ZN(new_n1211));
  AND2_X1   g1011(.A1(new_n702), .A2(G128), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n720), .A2(new_n724), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n260), .B1(new_n766), .B2(new_n758), .C1(new_n722), .C2(new_n984), .ZN(new_n1214));
  NOR4_X1   g1014(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .A4(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n690), .B1(new_n1209), .B2(new_n1215), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n755), .B(new_n1216), .C1(new_n829), .C2(new_n682), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(new_n214), .B2(new_n1125), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n1092), .B2(new_n945), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1201), .A2(new_n1219), .ZN(G381));
  AND2_X1   g1020(.A1(new_n1164), .A2(new_n1168), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1153), .B(new_n1158), .C1(new_n1167), .C2(new_n1160), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n635), .B1(new_n1222), .B2(new_n1129), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1196), .B1(new_n1221), .B2(new_n1223), .ZN(new_n1224));
  AND2_X1   g1024(.A1(new_n1103), .A2(new_n1127), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  AND2_X1   g1026(.A1(new_n1046), .A2(new_n1044), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n946), .A2(new_n1227), .A3(new_n976), .A4(new_n1023), .ZN(new_n1228));
  INV_X1    g1028(.A(G396), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n982), .A2(new_n1229), .A3(new_n1014), .ZN(new_n1230));
  NOR3_X1   g1030(.A1(new_n1226), .A2(new_n1228), .A3(new_n1230), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1231), .A2(new_n782), .A3(new_n1219), .A4(new_n1201), .ZN(G407));
  OAI211_X1 g1032(.A(G407), .B(G213), .C1(G343), .C2(new_n1226), .ZN(G409));
  INV_X1    g1033(.A(G213), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1234), .A2(G343), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  OR3_X1    g1036(.A1(new_n1159), .A2(new_n919), .A3(new_n1161), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1156), .A2(new_n945), .A3(new_n1157), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1225), .A2(new_n1237), .A3(new_n1195), .A4(new_n1238), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1236), .B(new_n1239), .C1(new_n1224), .C2(new_n1225), .ZN(new_n1240));
  OAI21_X1  g1040(.A(KEYINPUT60), .B1(new_n1093), .B2(new_n1199), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT60), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1242), .B1(new_n1079), .B2(new_n1092), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1241), .A2(new_n634), .A3(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1244), .A2(new_n782), .A3(new_n1219), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n782), .B1(new_n1244), .B2(new_n1219), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(KEYINPUT62), .B1(new_n1240), .B2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1235), .A2(G2897), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1247), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1251), .B1(new_n1252), .B2(new_n1245), .ZN(new_n1253));
  NOR3_X1   g1053(.A1(new_n1246), .A2(new_n1247), .A3(new_n1250), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(KEYINPUT61), .B1(new_n1240), .B2(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1235), .B1(G375), .B2(G378), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT62), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1248), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1257), .A2(new_n1258), .A3(new_n1259), .A4(new_n1239), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1249), .A2(new_n1256), .A3(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n908), .A2(new_n915), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n913), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n911), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n942), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n941), .A2(new_n655), .A3(new_n670), .A4(new_n939), .ZN(new_n1266));
  AOI21_X1  g1066(.A(KEYINPUT102), .B1(new_n933), .B2(new_n627), .ZN(new_n1267));
  NOR3_X1   g1067(.A1(new_n1265), .A2(new_n1266), .A3(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n918), .B1(new_n1268), .B2(new_n671), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n945), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1264), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  OAI21_X1  g1071(.A(G390), .B1(new_n1271), .B2(new_n975), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n1228), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(G393), .A2(G396), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n1230), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1273), .A2(KEYINPUT126), .A3(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT126), .ZN(new_n1278));
  AND3_X1   g1078(.A1(new_n982), .A2(new_n1229), .A3(new_n1014), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1229), .B1(new_n982), .B2(new_n1014), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1278), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1274), .A2(KEYINPUT126), .A3(new_n1230), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1281), .A2(new_n1272), .A3(new_n1282), .A4(new_n1228), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1277), .A2(KEYINPUT127), .A3(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(KEYINPUT127), .B1(new_n1277), .B2(new_n1283), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1261), .A2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1277), .A2(new_n1283), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1225), .B1(new_n1169), .B2(new_n1197), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n1195), .B(new_n1238), .C1(new_n1222), .C2(new_n919), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1291), .A2(G378), .ZN(new_n1292));
  NOR4_X1   g1092(.A1(new_n1290), .A2(new_n1292), .A3(new_n1248), .A4(new_n1235), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1289), .B1(new_n1293), .B2(KEYINPUT63), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(G375), .A2(G378), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1295), .A2(new_n1236), .A3(new_n1259), .A4(new_n1239), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT63), .ZN(new_n1297));
  AOI21_X1  g1097(.A(KEYINPUT61), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT124), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1240), .A2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT125), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1301), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1250), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1252), .A2(new_n1251), .A3(new_n1245), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1303), .A2(new_n1304), .A3(KEYINPUT125), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1302), .A2(new_n1305), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1295), .A2(KEYINPUT124), .A3(new_n1236), .A4(new_n1239), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1300), .A2(new_n1306), .A3(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1294), .A2(new_n1298), .A3(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1288), .A2(new_n1309), .ZN(G405));
  OAI21_X1  g1110(.A(new_n1248), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1311));
  AND2_X1   g1111(.A1(new_n1295), .A2(new_n1226), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT127), .ZN(new_n1313));
  AOI211_X1 g1113(.A(new_n1278), .B(new_n1275), .C1(new_n1272), .C2(new_n1228), .ZN(new_n1314));
  AND4_X1   g1114(.A1(new_n1228), .A2(new_n1281), .A3(new_n1272), .A4(new_n1282), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1313), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1316), .A2(new_n1284), .A3(new_n1259), .ZN(new_n1317));
  AND3_X1   g1117(.A1(new_n1311), .A2(new_n1312), .A3(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1312), .B1(new_n1311), .B2(new_n1317), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1318), .A2(new_n1319), .ZN(G402));
endmodule


