

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U551 ( .A(n816), .B(n971), .ZN(n771) );
  NOR2_X2 U552 ( .A1(n560), .A2(n559), .ZN(G160) );
  NOR2_X2 U553 ( .A1(n545), .A2(n544), .ZN(n556) );
  AND2_X1 U554 ( .A1(n703), .A2(n702), .ZN(n516) );
  XNOR2_X1 U555 ( .A(n630), .B(KEYINPUT27), .ZN(n631) );
  XNOR2_X1 U556 ( .A(n632), .B(n631), .ZN(n634) );
  INV_X1 U557 ( .A(n689), .ZN(n666) );
  INV_X1 U558 ( .A(KEYINPUT29), .ZN(n681) );
  XNOR2_X1 U559 ( .A(n682), .B(n681), .ZN(n685) );
  NAND2_X1 U560 ( .A1(n619), .A2(n618), .ZN(n689) );
  XNOR2_X1 U561 ( .A(G305), .B(n771), .ZN(n774) );
  NOR2_X1 U562 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U563 ( .A(G303), .B(G290), .ZN(n779) );
  XNOR2_X1 U564 ( .A(n780), .B(n779), .ZN(n813) );
  NOR2_X1 U565 ( .A1(G651), .A2(G543), .ZN(n761) );
  NOR2_X1 U566 ( .A1(G651), .A2(n581), .ZN(n765) );
  NAND2_X1 U567 ( .A1(G88), .A2(n761), .ZN(n518) );
  XOR2_X1 U568 ( .A(G543), .B(KEYINPUT0), .Z(n581) );
  INV_X1 U569 ( .A(G651), .ZN(n519) );
  NOR2_X1 U570 ( .A1(n581), .A2(n519), .ZN(n762) );
  NAND2_X1 U571 ( .A1(G75), .A2(n762), .ZN(n517) );
  NAND2_X1 U572 ( .A1(n518), .A2(n517), .ZN(n525) );
  NAND2_X1 U573 ( .A1(G50), .A2(n765), .ZN(n523) );
  NOR2_X1 U574 ( .A1(G543), .A2(n519), .ZN(n520) );
  XOR2_X1 U575 ( .A(KEYINPUT66), .B(n520), .Z(n521) );
  XNOR2_X2 U576 ( .A(KEYINPUT1), .B(n521), .ZN(n759) );
  NAND2_X1 U577 ( .A1(G62), .A2(n759), .ZN(n522) );
  NAND2_X1 U578 ( .A1(n523), .A2(n522), .ZN(n524) );
  NOR2_X1 U579 ( .A1(n525), .A2(n524), .ZN(G166) );
  INV_X1 U580 ( .A(G166), .ZN(G303) );
  NAND2_X1 U581 ( .A1(G47), .A2(n765), .ZN(n527) );
  NAND2_X1 U582 ( .A1(G60), .A2(n759), .ZN(n526) );
  NAND2_X1 U583 ( .A1(n527), .A2(n526), .ZN(n531) );
  NAND2_X1 U584 ( .A1(G85), .A2(n761), .ZN(n529) );
  NAND2_X1 U585 ( .A1(G72), .A2(n762), .ZN(n528) );
  NAND2_X1 U586 ( .A1(n529), .A2(n528), .ZN(n530) );
  OR2_X1 U587 ( .A1(n531), .A2(n530), .ZN(G290) );
  NAND2_X1 U588 ( .A1(G73), .A2(n762), .ZN(n532) );
  XOR2_X1 U589 ( .A(KEYINPUT2), .B(n532), .Z(n535) );
  NAND2_X1 U590 ( .A1(G61), .A2(n759), .ZN(n533) );
  XOR2_X1 U591 ( .A(KEYINPUT80), .B(n533), .Z(n534) );
  NOR2_X1 U592 ( .A1(n535), .A2(n534), .ZN(n537) );
  NAND2_X1 U593 ( .A1(n761), .A2(G86), .ZN(n536) );
  NAND2_X1 U594 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U595 ( .A(n538), .B(KEYINPUT81), .ZN(n540) );
  NAND2_X1 U596 ( .A1(G48), .A2(n765), .ZN(n539) );
  NAND2_X1 U597 ( .A1(n540), .A2(n539), .ZN(G305) );
  XNOR2_X1 U598 ( .A(KEYINPUT64), .B(G2104), .ZN(n545) );
  INV_X1 U599 ( .A(G2105), .ZN(n544) );
  AND2_X2 U600 ( .A1(n545), .A2(n544), .ZN(n870) );
  NAND2_X1 U601 ( .A1(n870), .A2(G102), .ZN(n543) );
  NOR2_X1 U602 ( .A1(G2104), .A2(G2105), .ZN(n541) );
  XOR2_X2 U603 ( .A(KEYINPUT17), .B(n541), .Z(n869) );
  NAND2_X1 U604 ( .A1(n869), .A2(G138), .ZN(n542) );
  NAND2_X1 U605 ( .A1(n543), .A2(n542), .ZN(n550) );
  AND2_X1 U606 ( .A1(G2104), .A2(G2105), .ZN(n873) );
  NAND2_X1 U607 ( .A1(G114), .A2(n873), .ZN(n547) );
  NAND2_X1 U608 ( .A1(G126), .A2(n556), .ZN(n546) );
  NAND2_X1 U609 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U610 ( .A(KEYINPUT85), .B(n548), .Z(n549) );
  NOR2_X1 U611 ( .A1(n550), .A2(n549), .ZN(G164) );
  INV_X1 U612 ( .A(KEYINPUT23), .ZN(n552) );
  NAND2_X1 U613 ( .A1(G101), .A2(n870), .ZN(n551) );
  XNOR2_X1 U614 ( .A(n552), .B(n551), .ZN(n555) );
  NAND2_X1 U615 ( .A1(G113), .A2(n873), .ZN(n553) );
  XOR2_X1 U616 ( .A(KEYINPUT65), .B(n553), .Z(n554) );
  NAND2_X1 U617 ( .A1(n555), .A2(n554), .ZN(n560) );
  NAND2_X1 U618 ( .A1(G125), .A2(n556), .ZN(n558) );
  NAND2_X1 U619 ( .A1(G137), .A2(n869), .ZN(n557) );
  NAND2_X1 U620 ( .A1(n558), .A2(n557), .ZN(n559) );
  NAND2_X1 U621 ( .A1(G89), .A2(n761), .ZN(n561) );
  XOR2_X1 U622 ( .A(KEYINPUT75), .B(n561), .Z(n562) );
  XNOR2_X1 U623 ( .A(n562), .B(KEYINPUT4), .ZN(n564) );
  NAND2_X1 U624 ( .A1(G76), .A2(n762), .ZN(n563) );
  NAND2_X1 U625 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U626 ( .A(n565), .B(KEYINPUT5), .ZN(n570) );
  NAND2_X1 U627 ( .A1(G51), .A2(n765), .ZN(n567) );
  NAND2_X1 U628 ( .A1(G63), .A2(n759), .ZN(n566) );
  NAND2_X1 U629 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U630 ( .A(KEYINPUT6), .B(n568), .Z(n569) );
  NAND2_X1 U631 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U632 ( .A(n571), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U633 ( .A1(G64), .A2(n759), .ZN(n572) );
  XOR2_X1 U634 ( .A(KEYINPUT67), .B(n572), .Z(n574) );
  NAND2_X1 U635 ( .A1(n765), .A2(G52), .ZN(n573) );
  NAND2_X1 U636 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U637 ( .A(KEYINPUT68), .B(n575), .ZN(n580) );
  NAND2_X1 U638 ( .A1(G90), .A2(n761), .ZN(n577) );
  NAND2_X1 U639 ( .A1(G77), .A2(n762), .ZN(n576) );
  NAND2_X1 U640 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U641 ( .A(KEYINPUT9), .B(n578), .Z(n579) );
  NOR2_X1 U642 ( .A1(n580), .A2(n579), .ZN(G171) );
  INV_X1 U643 ( .A(G171), .ZN(G301) );
  XOR2_X1 U644 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U645 ( .A1(G87), .A2(n581), .ZN(n583) );
  NAND2_X1 U646 ( .A1(G74), .A2(G651), .ZN(n582) );
  NAND2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U648 ( .A1(n759), .A2(n584), .ZN(n586) );
  NAND2_X1 U649 ( .A1(n765), .A2(G49), .ZN(n585) );
  NAND2_X1 U650 ( .A1(n586), .A2(n585), .ZN(G288) );
  NAND2_X1 U651 ( .A1(G107), .A2(n873), .ZN(n588) );
  NAND2_X1 U652 ( .A1(G131), .A2(n869), .ZN(n587) );
  NAND2_X1 U653 ( .A1(n588), .A2(n587), .ZN(n592) );
  NAND2_X1 U654 ( .A1(G119), .A2(n556), .ZN(n590) );
  NAND2_X1 U655 ( .A1(G95), .A2(n870), .ZN(n589) );
  NAND2_X1 U656 ( .A1(n590), .A2(n589), .ZN(n591) );
  OR2_X1 U657 ( .A1(n592), .A2(n591), .ZN(n886) );
  NAND2_X1 U658 ( .A1(G1991), .A2(n886), .ZN(n602) );
  NAND2_X1 U659 ( .A1(G105), .A2(n870), .ZN(n593) );
  XNOR2_X1 U660 ( .A(n593), .B(KEYINPUT38), .ZN(n600) );
  NAND2_X1 U661 ( .A1(G129), .A2(n556), .ZN(n595) );
  NAND2_X1 U662 ( .A1(G141), .A2(n869), .ZN(n594) );
  NAND2_X1 U663 ( .A1(n595), .A2(n594), .ZN(n598) );
  NAND2_X1 U664 ( .A1(G117), .A2(n873), .ZN(n596) );
  XNOR2_X1 U665 ( .A(KEYINPUT89), .B(n596), .ZN(n597) );
  NOR2_X1 U666 ( .A1(n598), .A2(n597), .ZN(n599) );
  NAND2_X1 U667 ( .A1(n600), .A2(n599), .ZN(n865) );
  NAND2_X1 U668 ( .A1(G1996), .A2(n865), .ZN(n601) );
  NAND2_X1 U669 ( .A1(n602), .A2(n601), .ZN(n929) );
  NOR2_X1 U670 ( .A1(G164), .A2(G1384), .ZN(n619) );
  NAND2_X1 U671 ( .A1(G160), .A2(G40), .ZN(n617) );
  NOR2_X1 U672 ( .A1(n619), .A2(n617), .ZN(n744) );
  NAND2_X1 U673 ( .A1(n929), .A2(n744), .ZN(n603) );
  XOR2_X1 U674 ( .A(KEYINPUT90), .B(n603), .Z(n737) );
  INV_X1 U675 ( .A(n737), .ZN(n616) );
  XNOR2_X1 U676 ( .A(G2067), .B(KEYINPUT37), .ZN(n742) );
  NAND2_X1 U677 ( .A1(G140), .A2(n869), .ZN(n605) );
  NAND2_X1 U678 ( .A1(G104), .A2(n870), .ZN(n604) );
  NAND2_X1 U679 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U680 ( .A(KEYINPUT34), .B(n606), .ZN(n614) );
  NAND2_X1 U681 ( .A1(n873), .A2(G116), .ZN(n607) );
  XNOR2_X1 U682 ( .A(KEYINPUT87), .B(n607), .ZN(n610) );
  NAND2_X1 U683 ( .A1(n556), .A2(G128), .ZN(n608) );
  XOR2_X1 U684 ( .A(n608), .B(KEYINPUT86), .Z(n609) );
  NOR2_X1 U685 ( .A1(n610), .A2(n609), .ZN(n611) );
  XOR2_X1 U686 ( .A(KEYINPUT35), .B(n611), .Z(n612) );
  XOR2_X1 U687 ( .A(KEYINPUT88), .B(n612), .Z(n613) );
  NOR2_X1 U688 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U689 ( .A(KEYINPUT36), .B(n615), .ZN(n887) );
  NOR2_X1 U690 ( .A1(n742), .A2(n887), .ZN(n932) );
  NAND2_X1 U691 ( .A1(n744), .A2(n932), .ZN(n740) );
  NAND2_X1 U692 ( .A1(n616), .A2(n740), .ZN(n730) );
  INV_X1 U693 ( .A(n617), .ZN(n618) );
  NAND2_X1 U694 ( .A1(G8), .A2(n689), .ZN(n725) );
  NOR2_X1 U695 ( .A1(G1966), .A2(n725), .ZN(n697) );
  NOR2_X1 U696 ( .A1(n689), .A2(G2084), .ZN(n620) );
  XNOR2_X1 U697 ( .A(n620), .B(KEYINPUT91), .ZN(n699) );
  NAND2_X1 U698 ( .A1(G8), .A2(n699), .ZN(n621) );
  NOR2_X1 U699 ( .A1(n697), .A2(n621), .ZN(n622) );
  XNOR2_X1 U700 ( .A(n622), .B(KEYINPUT30), .ZN(n624) );
  INV_X1 U701 ( .A(G168), .ZN(n623) );
  NAND2_X1 U702 ( .A1(n624), .A2(n623), .ZN(n628) );
  XOR2_X1 U703 ( .A(G2078), .B(KEYINPUT25), .Z(n945) );
  NOR2_X1 U704 ( .A1(n945), .A2(n689), .ZN(n626) );
  NOR2_X1 U705 ( .A1(n666), .A2(G1961), .ZN(n625) );
  NOR2_X1 U706 ( .A1(n626), .A2(n625), .ZN(n683) );
  NAND2_X1 U707 ( .A1(n683), .A2(G301), .ZN(n627) );
  NAND2_X1 U708 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U709 ( .A(n629), .B(KEYINPUT31), .ZN(n687) );
  NAND2_X1 U710 ( .A1(G2072), .A2(n666), .ZN(n632) );
  INV_X1 U711 ( .A(KEYINPUT93), .ZN(n630) );
  INV_X1 U712 ( .A(G1956), .ZN(n996) );
  NOR2_X1 U713 ( .A1(n666), .A2(n996), .ZN(n633) );
  NOR2_X1 U714 ( .A1(n634), .A2(n633), .ZN(n676) );
  NAND2_X1 U715 ( .A1(G53), .A2(n765), .ZN(n636) );
  NAND2_X1 U716 ( .A1(G65), .A2(n759), .ZN(n635) );
  NAND2_X1 U717 ( .A1(n636), .A2(n635), .ZN(n640) );
  NAND2_X1 U718 ( .A1(G91), .A2(n761), .ZN(n638) );
  NAND2_X1 U719 ( .A1(G78), .A2(n762), .ZN(n637) );
  NAND2_X1 U720 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U721 ( .A1(n640), .A2(n639), .ZN(n971) );
  NAND2_X1 U722 ( .A1(n676), .A2(n971), .ZN(n675) );
  NAND2_X1 U723 ( .A1(n762), .A2(G79), .ZN(n647) );
  NAND2_X1 U724 ( .A1(G54), .A2(n765), .ZN(n642) );
  NAND2_X1 U725 ( .A1(G66), .A2(n759), .ZN(n641) );
  NAND2_X1 U726 ( .A1(n642), .A2(n641), .ZN(n645) );
  NAND2_X1 U727 ( .A1(G92), .A2(n761), .ZN(n643) );
  XNOR2_X1 U728 ( .A(KEYINPUT73), .B(n643), .ZN(n644) );
  NOR2_X1 U729 ( .A1(n645), .A2(n644), .ZN(n646) );
  NAND2_X1 U730 ( .A1(n647), .A2(n646), .ZN(n648) );
  XOR2_X1 U731 ( .A(KEYINPUT15), .B(n648), .Z(n976) );
  NAND2_X1 U732 ( .A1(G43), .A2(n765), .ZN(n658) );
  NAND2_X1 U733 ( .A1(G56), .A2(n759), .ZN(n649) );
  XNOR2_X1 U734 ( .A(n649), .B(KEYINPUT14), .ZN(n655) );
  NAND2_X1 U735 ( .A1(n761), .A2(G81), .ZN(n650) );
  XNOR2_X1 U736 ( .A(n650), .B(KEYINPUT12), .ZN(n652) );
  NAND2_X1 U737 ( .A1(G68), .A2(n762), .ZN(n651) );
  NAND2_X1 U738 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U739 ( .A(KEYINPUT13), .B(n653), .ZN(n654) );
  NAND2_X1 U740 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U741 ( .A(n656), .B(KEYINPUT71), .ZN(n657) );
  NAND2_X1 U742 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U743 ( .A(n659), .B(KEYINPUT72), .ZN(n981) );
  XOR2_X1 U744 ( .A(KEYINPUT26), .B(KEYINPUT96), .Z(n661) );
  XOR2_X1 U745 ( .A(G1996), .B(KEYINPUT95), .Z(n943) );
  NAND2_X1 U746 ( .A1(n943), .A2(n666), .ZN(n660) );
  XNOR2_X1 U747 ( .A(n661), .B(n660), .ZN(n662) );
  NOR2_X1 U748 ( .A1(n981), .A2(n662), .ZN(n664) );
  NAND2_X1 U749 ( .A1(G1341), .A2(n689), .ZN(n663) );
  NAND2_X1 U750 ( .A1(n664), .A2(n663), .ZN(n671) );
  OR2_X1 U751 ( .A1(n976), .A2(n671), .ZN(n670) );
  AND2_X1 U752 ( .A1(n689), .A2(G1348), .ZN(n665) );
  XNOR2_X1 U753 ( .A(n665), .B(KEYINPUT97), .ZN(n668) );
  NAND2_X1 U754 ( .A1(n666), .A2(G2067), .ZN(n667) );
  NAND2_X1 U755 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U756 ( .A1(n670), .A2(n669), .ZN(n673) );
  NAND2_X1 U757 ( .A1(n976), .A2(n671), .ZN(n672) );
  NAND2_X1 U758 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U759 ( .A1(n675), .A2(n674), .ZN(n680) );
  NOR2_X1 U760 ( .A1(n676), .A2(n971), .ZN(n678) );
  XOR2_X1 U761 ( .A(KEYINPUT28), .B(KEYINPUT94), .Z(n677) );
  XNOR2_X1 U762 ( .A(n678), .B(n677), .ZN(n679) );
  NAND2_X1 U763 ( .A1(n680), .A2(n679), .ZN(n682) );
  OR2_X1 U764 ( .A1(G301), .A2(n683), .ZN(n684) );
  NAND2_X1 U765 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U766 ( .A1(n687), .A2(n686), .ZN(n698) );
  NAND2_X1 U767 ( .A1(n698), .A2(G286), .ZN(n694) );
  NOR2_X1 U768 ( .A1(G1971), .A2(n725), .ZN(n688) );
  XNOR2_X1 U769 ( .A(KEYINPUT99), .B(n688), .ZN(n692) );
  NOR2_X1 U770 ( .A1(G2090), .A2(n689), .ZN(n690) );
  NOR2_X1 U771 ( .A1(G166), .A2(n690), .ZN(n691) );
  NAND2_X1 U772 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U773 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U774 ( .A1(n695), .A2(G8), .ZN(n696) );
  XNOR2_X1 U775 ( .A(n696), .B(KEYINPUT32), .ZN(n706) );
  INV_X1 U776 ( .A(n697), .ZN(n704) );
  XNOR2_X1 U777 ( .A(n698), .B(KEYINPUT98), .ZN(n703) );
  INV_X1 U778 ( .A(n699), .ZN(n700) );
  NAND2_X1 U779 ( .A1(n700), .A2(G8), .ZN(n701) );
  XNOR2_X1 U780 ( .A(n701), .B(KEYINPUT92), .ZN(n702) );
  NAND2_X1 U781 ( .A1(n704), .A2(n516), .ZN(n705) );
  NAND2_X1 U782 ( .A1(n706), .A2(n705), .ZN(n719) );
  NOR2_X1 U783 ( .A1(G1976), .A2(G288), .ZN(n712) );
  NOR2_X1 U784 ( .A1(G1971), .A2(G303), .ZN(n707) );
  NOR2_X1 U785 ( .A1(n712), .A2(n707), .ZN(n972) );
  NAND2_X1 U786 ( .A1(n719), .A2(n972), .ZN(n710) );
  INV_X1 U787 ( .A(n725), .ZN(n708) );
  NAND2_X1 U788 ( .A1(G1976), .A2(G288), .ZN(n970) );
  AND2_X1 U789 ( .A1(n708), .A2(n970), .ZN(n709) );
  AND2_X1 U790 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U791 ( .A1(n711), .A2(KEYINPUT33), .ZN(n715) );
  NAND2_X1 U792 ( .A1(n712), .A2(KEYINPUT33), .ZN(n713) );
  NOR2_X1 U793 ( .A1(n713), .A2(n725), .ZN(n714) );
  NOR2_X1 U794 ( .A1(n715), .A2(n714), .ZN(n716) );
  XOR2_X1 U795 ( .A(G1981), .B(G305), .Z(n966) );
  NAND2_X1 U796 ( .A1(n716), .A2(n966), .ZN(n722) );
  NOR2_X1 U797 ( .A1(G2090), .A2(G303), .ZN(n717) );
  NAND2_X1 U798 ( .A1(G8), .A2(n717), .ZN(n718) );
  NAND2_X1 U799 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U800 ( .A1(n720), .A2(n725), .ZN(n721) );
  NAND2_X1 U801 ( .A1(n722), .A2(n721), .ZN(n727) );
  NOR2_X1 U802 ( .A1(G1981), .A2(G305), .ZN(n723) );
  XOR2_X1 U803 ( .A(n723), .B(KEYINPUT24), .Z(n724) );
  NOR2_X1 U804 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U805 ( .A(n728), .B(KEYINPUT100), .ZN(n729) );
  NOR2_X1 U806 ( .A1(n730), .A2(n729), .ZN(n732) );
  XNOR2_X1 U807 ( .A(G1986), .B(G290), .ZN(n978) );
  NAND2_X1 U808 ( .A1(n978), .A2(n744), .ZN(n731) );
  NAND2_X1 U809 ( .A1(n732), .A2(n731), .ZN(n747) );
  NOR2_X1 U810 ( .A1(G1996), .A2(n865), .ZN(n921) );
  NOR2_X1 U811 ( .A1(G1991), .A2(n886), .ZN(n733) );
  XOR2_X1 U812 ( .A(KEYINPUT101), .B(n733), .Z(n927) );
  NOR2_X1 U813 ( .A1(G1986), .A2(G290), .ZN(n734) );
  NOR2_X1 U814 ( .A1(n927), .A2(n734), .ZN(n735) );
  XNOR2_X1 U815 ( .A(n735), .B(KEYINPUT102), .ZN(n736) );
  NOR2_X1 U816 ( .A1(n737), .A2(n736), .ZN(n738) );
  NOR2_X1 U817 ( .A1(n921), .A2(n738), .ZN(n739) );
  XNOR2_X1 U818 ( .A(KEYINPUT39), .B(n739), .ZN(n741) );
  NAND2_X1 U819 ( .A1(n741), .A2(n740), .ZN(n743) );
  NAND2_X1 U820 ( .A1(n742), .A2(n887), .ZN(n918) );
  NAND2_X1 U821 ( .A1(n743), .A2(n918), .ZN(n745) );
  NAND2_X1 U822 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U823 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U824 ( .A(n748), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U825 ( .A(G2435), .B(G2454), .Z(n750) );
  XNOR2_X1 U826 ( .A(KEYINPUT103), .B(G2438), .ZN(n749) );
  XNOR2_X1 U827 ( .A(n750), .B(n749), .ZN(n757) );
  XOR2_X1 U828 ( .A(G2446), .B(G2430), .Z(n752) );
  XNOR2_X1 U829 ( .A(G2451), .B(G2443), .ZN(n751) );
  XNOR2_X1 U830 ( .A(n752), .B(n751), .ZN(n753) );
  XOR2_X1 U831 ( .A(n753), .B(G2427), .Z(n755) );
  XNOR2_X1 U832 ( .A(G1341), .B(G1348), .ZN(n754) );
  XNOR2_X1 U833 ( .A(n755), .B(n754), .ZN(n756) );
  XNOR2_X1 U834 ( .A(n757), .B(n756), .ZN(n758) );
  AND2_X1 U835 ( .A1(n758), .A2(G14), .ZN(G401) );
  AND2_X1 U836 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U837 ( .A(G108), .ZN(G238) );
  INV_X1 U838 ( .A(G132), .ZN(G219) );
  INV_X1 U839 ( .A(G82), .ZN(G220) );
  NAND2_X1 U840 ( .A1(n759), .A2(G67), .ZN(n760) );
  XNOR2_X1 U841 ( .A(n760), .B(KEYINPUT78), .ZN(n770) );
  NAND2_X1 U842 ( .A1(G93), .A2(n761), .ZN(n764) );
  NAND2_X1 U843 ( .A1(G80), .A2(n762), .ZN(n763) );
  NAND2_X1 U844 ( .A1(n764), .A2(n763), .ZN(n768) );
  NAND2_X1 U845 ( .A1(G55), .A2(n765), .ZN(n766) );
  XNOR2_X1 U846 ( .A(KEYINPUT79), .B(n766), .ZN(n767) );
  NOR2_X1 U847 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U848 ( .A1(n770), .A2(n769), .ZN(n816) );
  INV_X1 U849 ( .A(n774), .ZN(n773) );
  INV_X1 U850 ( .A(KEYINPUT82), .ZN(n772) );
  NAND2_X1 U851 ( .A1(n773), .A2(n772), .ZN(n776) );
  NAND2_X1 U852 ( .A1(KEYINPUT82), .A2(n774), .ZN(n775) );
  NAND2_X1 U853 ( .A1(n776), .A2(n775), .ZN(n778) );
  XNOR2_X1 U854 ( .A(G288), .B(KEYINPUT19), .ZN(n777) );
  XNOR2_X1 U855 ( .A(n778), .B(n777), .ZN(n780) );
  XOR2_X1 U856 ( .A(n813), .B(G286), .Z(n783) );
  INV_X1 U857 ( .A(n976), .ZN(n809) );
  XNOR2_X1 U858 ( .A(G171), .B(n809), .ZN(n781) );
  XNOR2_X1 U859 ( .A(n781), .B(n981), .ZN(n782) );
  XNOR2_X1 U860 ( .A(n783), .B(n782), .ZN(n784) );
  NOR2_X1 U861 ( .A1(G37), .A2(n784), .ZN(G397) );
  XOR2_X1 U862 ( .A(KEYINPUT69), .B(KEYINPUT10), .Z(n786) );
  NAND2_X1 U863 ( .A1(G7), .A2(G661), .ZN(n785) );
  XNOR2_X1 U864 ( .A(n786), .B(n785), .ZN(G223) );
  XOR2_X1 U865 ( .A(G223), .B(KEYINPUT70), .Z(n835) );
  NAND2_X1 U866 ( .A1(n835), .A2(G567), .ZN(n787) );
  XOR2_X1 U867 ( .A(KEYINPUT11), .B(n787), .Z(G234) );
  INV_X1 U868 ( .A(G860), .ZN(n794) );
  OR2_X1 U869 ( .A1(n794), .A2(n981), .ZN(G153) );
  NOR2_X1 U870 ( .A1(G868), .A2(n976), .ZN(n789) );
  INV_X1 U871 ( .A(G868), .ZN(n817) );
  NOR2_X1 U872 ( .A1(n817), .A2(G301), .ZN(n788) );
  NOR2_X1 U873 ( .A1(n789), .A2(n788), .ZN(n790) );
  XNOR2_X1 U874 ( .A(KEYINPUT74), .B(n790), .ZN(G284) );
  INV_X1 U875 ( .A(n971), .ZN(G299) );
  XNOR2_X1 U876 ( .A(KEYINPUT76), .B(n817), .ZN(n791) );
  NOR2_X1 U877 ( .A1(G286), .A2(n791), .ZN(n793) );
  NOR2_X1 U878 ( .A1(G868), .A2(G299), .ZN(n792) );
  NOR2_X1 U879 ( .A1(n793), .A2(n792), .ZN(G297) );
  NAND2_X1 U880 ( .A1(n794), .A2(G559), .ZN(n795) );
  NAND2_X1 U881 ( .A1(n795), .A2(n809), .ZN(n796) );
  XNOR2_X1 U882 ( .A(n796), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U883 ( .A1(n981), .A2(G868), .ZN(n799) );
  NAND2_X1 U884 ( .A1(G868), .A2(n809), .ZN(n797) );
  NOR2_X1 U885 ( .A1(G559), .A2(n797), .ZN(n798) );
  NOR2_X1 U886 ( .A1(n799), .A2(n798), .ZN(G282) );
  NAND2_X1 U887 ( .A1(G111), .A2(n873), .ZN(n801) );
  NAND2_X1 U888 ( .A1(G135), .A2(n869), .ZN(n800) );
  NAND2_X1 U889 ( .A1(n801), .A2(n800), .ZN(n804) );
  NAND2_X1 U890 ( .A1(n556), .A2(G123), .ZN(n802) );
  XOR2_X1 U891 ( .A(KEYINPUT18), .B(n802), .Z(n803) );
  NOR2_X1 U892 ( .A1(n804), .A2(n803), .ZN(n806) );
  NAND2_X1 U893 ( .A1(n870), .A2(G99), .ZN(n805) );
  NAND2_X1 U894 ( .A1(n806), .A2(n805), .ZN(n867) );
  INV_X1 U895 ( .A(n867), .ZN(n926) );
  XNOR2_X1 U896 ( .A(n926), .B(G2096), .ZN(n808) );
  INV_X1 U897 ( .A(G2100), .ZN(n807) );
  NAND2_X1 U898 ( .A1(n808), .A2(n807), .ZN(G156) );
  NAND2_X1 U899 ( .A1(G559), .A2(n809), .ZN(n810) );
  XNOR2_X1 U900 ( .A(n810), .B(n981), .ZN(n814) );
  NOR2_X1 U901 ( .A1(G860), .A2(n814), .ZN(n811) );
  XNOR2_X1 U902 ( .A(n811), .B(KEYINPUT77), .ZN(n812) );
  XNOR2_X1 U903 ( .A(n816), .B(n812), .ZN(G145) );
  XNOR2_X1 U904 ( .A(n814), .B(n813), .ZN(n815) );
  NAND2_X1 U905 ( .A1(n815), .A2(G868), .ZN(n819) );
  NAND2_X1 U906 ( .A1(n817), .A2(n816), .ZN(n818) );
  NAND2_X1 U907 ( .A1(n819), .A2(n818), .ZN(G295) );
  NAND2_X1 U908 ( .A1(G2084), .A2(G2078), .ZN(n820) );
  XOR2_X1 U909 ( .A(KEYINPUT20), .B(n820), .Z(n821) );
  NAND2_X1 U910 ( .A1(G2090), .A2(n821), .ZN(n823) );
  XOR2_X1 U911 ( .A(KEYINPUT83), .B(KEYINPUT21), .Z(n822) );
  XNOR2_X1 U912 ( .A(n823), .B(n822), .ZN(n824) );
  NAND2_X1 U913 ( .A1(G2072), .A2(n824), .ZN(G158) );
  XNOR2_X1 U914 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U915 ( .A1(G220), .A2(G219), .ZN(n825) );
  XOR2_X1 U916 ( .A(KEYINPUT22), .B(n825), .Z(n826) );
  NOR2_X1 U917 ( .A1(G218), .A2(n826), .ZN(n827) );
  NAND2_X1 U918 ( .A1(G96), .A2(n827), .ZN(n841) );
  AND2_X1 U919 ( .A1(G2106), .A2(n841), .ZN(n832) );
  NAND2_X1 U920 ( .A1(G120), .A2(G69), .ZN(n828) );
  NOR2_X1 U921 ( .A1(G238), .A2(n828), .ZN(n829) );
  NAND2_X1 U922 ( .A1(G57), .A2(n829), .ZN(n840) );
  NAND2_X1 U923 ( .A1(G567), .A2(n840), .ZN(n830) );
  XOR2_X1 U924 ( .A(KEYINPUT84), .B(n830), .Z(n831) );
  NOR2_X1 U925 ( .A1(n832), .A2(n831), .ZN(G319) );
  INV_X1 U926 ( .A(G319), .ZN(n834) );
  NAND2_X1 U927 ( .A1(G661), .A2(G483), .ZN(n833) );
  NOR2_X1 U928 ( .A1(n834), .A2(n833), .ZN(n839) );
  NAND2_X1 U929 ( .A1(n839), .A2(G36), .ZN(G176) );
  NAND2_X1 U930 ( .A1(n835), .A2(G2106), .ZN(n836) );
  XNOR2_X1 U931 ( .A(n836), .B(KEYINPUT104), .ZN(G217) );
  AND2_X1 U932 ( .A1(G15), .A2(G2), .ZN(n837) );
  NAND2_X1 U933 ( .A1(G661), .A2(n837), .ZN(G259) );
  NAND2_X1 U934 ( .A1(G3), .A2(G1), .ZN(n838) );
  NAND2_X1 U935 ( .A1(n839), .A2(n838), .ZN(G188) );
  XNOR2_X1 U936 ( .A(G120), .B(KEYINPUT105), .ZN(G236) );
  XOR2_X1 U937 ( .A(G69), .B(KEYINPUT106), .Z(G235) );
  INV_X1 U939 ( .A(G96), .ZN(G221) );
  NOR2_X1 U940 ( .A1(n841), .A2(n840), .ZN(G325) );
  INV_X1 U941 ( .A(G325), .ZN(G261) );
  NAND2_X1 U942 ( .A1(G136), .A2(n869), .ZN(n842) );
  XNOR2_X1 U943 ( .A(n842), .B(KEYINPUT108), .ZN(n846) );
  XOR2_X1 U944 ( .A(KEYINPUT107), .B(KEYINPUT44), .Z(n844) );
  NAND2_X1 U945 ( .A1(G124), .A2(n556), .ZN(n843) );
  XNOR2_X1 U946 ( .A(n844), .B(n843), .ZN(n845) );
  NAND2_X1 U947 ( .A1(n846), .A2(n845), .ZN(n851) );
  NAND2_X1 U948 ( .A1(G112), .A2(n873), .ZN(n848) );
  NAND2_X1 U949 ( .A1(G100), .A2(n870), .ZN(n847) );
  NAND2_X1 U950 ( .A1(n848), .A2(n847), .ZN(n849) );
  XOR2_X1 U951 ( .A(KEYINPUT109), .B(n849), .Z(n850) );
  NOR2_X1 U952 ( .A1(n851), .A2(n850), .ZN(G162) );
  XOR2_X1 U953 ( .A(KEYINPUT48), .B(KEYINPUT113), .Z(n853) );
  XNOR2_X1 U954 ( .A(KEYINPUT114), .B(KEYINPUT115), .ZN(n852) );
  XNOR2_X1 U955 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U956 ( .A(n854), .B(KEYINPUT46), .Z(n856) );
  XNOR2_X1 U957 ( .A(G162), .B(KEYINPUT112), .ZN(n855) );
  XNOR2_X1 U958 ( .A(n856), .B(n855), .ZN(n884) );
  NAND2_X1 U959 ( .A1(G118), .A2(n873), .ZN(n858) );
  NAND2_X1 U960 ( .A1(G130), .A2(n556), .ZN(n857) );
  NAND2_X1 U961 ( .A1(n858), .A2(n857), .ZN(n864) );
  NAND2_X1 U962 ( .A1(G142), .A2(n869), .ZN(n860) );
  NAND2_X1 U963 ( .A1(G106), .A2(n870), .ZN(n859) );
  NAND2_X1 U964 ( .A1(n860), .A2(n859), .ZN(n861) );
  XOR2_X1 U965 ( .A(KEYINPUT45), .B(n861), .Z(n862) );
  XNOR2_X1 U966 ( .A(KEYINPUT110), .B(n862), .ZN(n863) );
  NOR2_X1 U967 ( .A1(n864), .A2(n863), .ZN(n866) );
  XNOR2_X1 U968 ( .A(n866), .B(n865), .ZN(n868) );
  XNOR2_X1 U969 ( .A(n868), .B(n867), .ZN(n880) );
  NAND2_X1 U970 ( .A1(G139), .A2(n869), .ZN(n872) );
  NAND2_X1 U971 ( .A1(G103), .A2(n870), .ZN(n871) );
  NAND2_X1 U972 ( .A1(n872), .A2(n871), .ZN(n879) );
  NAND2_X1 U973 ( .A1(n873), .A2(G115), .ZN(n874) );
  XOR2_X1 U974 ( .A(KEYINPUT111), .B(n874), .Z(n876) );
  NAND2_X1 U975 ( .A1(n556), .A2(G127), .ZN(n875) );
  NAND2_X1 U976 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U977 ( .A(KEYINPUT47), .B(n877), .Z(n878) );
  NOR2_X1 U978 ( .A1(n879), .A2(n878), .ZN(n914) );
  XOR2_X1 U979 ( .A(n880), .B(n914), .Z(n882) );
  XNOR2_X1 U980 ( .A(G164), .B(G160), .ZN(n881) );
  XNOR2_X1 U981 ( .A(n882), .B(n881), .ZN(n883) );
  XOR2_X1 U982 ( .A(n884), .B(n883), .Z(n885) );
  XNOR2_X1 U983 ( .A(n886), .B(n885), .ZN(n888) );
  XOR2_X1 U984 ( .A(n888), .B(n887), .Z(n889) );
  NOR2_X1 U985 ( .A1(G37), .A2(n889), .ZN(G395) );
  XOR2_X1 U986 ( .A(G2100), .B(G2096), .Z(n891) );
  XNOR2_X1 U987 ( .A(KEYINPUT42), .B(G2678), .ZN(n890) );
  XNOR2_X1 U988 ( .A(n891), .B(n890), .ZN(n895) );
  XOR2_X1 U989 ( .A(KEYINPUT43), .B(G2090), .Z(n893) );
  XNOR2_X1 U990 ( .A(G2067), .B(G2072), .ZN(n892) );
  XNOR2_X1 U991 ( .A(n893), .B(n892), .ZN(n894) );
  XOR2_X1 U992 ( .A(n895), .B(n894), .Z(n897) );
  XNOR2_X1 U993 ( .A(G2084), .B(G2078), .ZN(n896) );
  XNOR2_X1 U994 ( .A(n897), .B(n896), .ZN(G227) );
  XOR2_X1 U995 ( .A(G1976), .B(G1981), .Z(n899) );
  XNOR2_X1 U996 ( .A(G1966), .B(G1971), .ZN(n898) );
  XNOR2_X1 U997 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U998 ( .A(n900), .B(G2474), .Z(n902) );
  XNOR2_X1 U999 ( .A(G1996), .B(G1991), .ZN(n901) );
  XNOR2_X1 U1000 ( .A(n902), .B(n901), .ZN(n906) );
  XOR2_X1 U1001 ( .A(KEYINPUT41), .B(G1956), .Z(n904) );
  XNOR2_X1 U1002 ( .A(G1986), .B(G1961), .ZN(n903) );
  XNOR2_X1 U1003 ( .A(n904), .B(n903), .ZN(n905) );
  XNOR2_X1 U1004 ( .A(n906), .B(n905), .ZN(G229) );
  NOR2_X1 U1005 ( .A1(G395), .A2(G397), .ZN(n907) );
  XOR2_X1 U1006 ( .A(KEYINPUT116), .B(n907), .Z(n908) );
  NOR2_X1 U1007 ( .A1(G401), .A2(n908), .ZN(n909) );
  NAND2_X1 U1008 ( .A1(G319), .A2(n909), .ZN(n912) );
  NOR2_X1 U1009 ( .A1(G227), .A2(G229), .ZN(n910) );
  XNOR2_X1 U1010 ( .A(KEYINPUT49), .B(n910), .ZN(n911) );
  NOR2_X1 U1011 ( .A1(n912), .A2(n911), .ZN(n913) );
  XNOR2_X1 U1012 ( .A(n913), .B(KEYINPUT117), .ZN(G225) );
  INV_X1 U1013 ( .A(G225), .ZN(G308) );
  INV_X1 U1014 ( .A(G57), .ZN(G237) );
  XOR2_X1 U1015 ( .A(G2072), .B(n914), .Z(n916) );
  XOR2_X1 U1016 ( .A(G164), .B(G2078), .Z(n915) );
  NOR2_X1 U1017 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1018 ( .A(n917), .B(KEYINPUT50), .ZN(n919) );
  NAND2_X1 U1019 ( .A1(n919), .A2(n918), .ZN(n925) );
  XOR2_X1 U1020 ( .A(G2090), .B(G162), .Z(n920) );
  NOR2_X1 U1021 ( .A1(n921), .A2(n920), .ZN(n922) );
  XOR2_X1 U1022 ( .A(KEYINPUT51), .B(n922), .Z(n923) );
  XOR2_X1 U1023 ( .A(KEYINPUT118), .B(n923), .Z(n924) );
  NOR2_X1 U1024 ( .A1(n925), .A2(n924), .ZN(n935) );
  NOR2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(n931) );
  XOR2_X1 U1026 ( .A(G160), .B(G2084), .Z(n928) );
  NOR2_X1 U1027 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n933) );
  NOR2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1031 ( .A(KEYINPUT52), .B(n936), .ZN(n937) );
  XNOR2_X1 U1032 ( .A(KEYINPUT119), .B(n937), .ZN(n938) );
  INV_X1 U1033 ( .A(KEYINPUT55), .ZN(n962) );
  NAND2_X1 U1034 ( .A1(n938), .A2(n962), .ZN(n939) );
  NAND2_X1 U1035 ( .A1(n939), .A2(G29), .ZN(n1022) );
  XNOR2_X1 U1036 ( .A(G2090), .B(G35), .ZN(n957) );
  XOR2_X1 U1037 ( .A(G1991), .B(G25), .Z(n940) );
  XNOR2_X1 U1038 ( .A(KEYINPUT120), .B(n940), .ZN(n941) );
  NAND2_X1 U1039 ( .A1(n941), .A2(G28), .ZN(n942) );
  XNOR2_X1 U1040 ( .A(n942), .B(KEYINPUT121), .ZN(n952) );
  XNOR2_X1 U1041 ( .A(G2067), .B(G26), .ZN(n950) );
  XNOR2_X1 U1042 ( .A(n943), .B(KEYINPUT122), .ZN(n944) );
  XNOR2_X1 U1043 ( .A(n944), .B(G32), .ZN(n947) );
  XNOR2_X1 U1044 ( .A(G27), .B(n945), .ZN(n946) );
  NOR2_X1 U1045 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1046 ( .A(n948), .B(KEYINPUT123), .ZN(n949) );
  NOR2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n954) );
  XNOR2_X1 U1049 ( .A(G33), .B(G2072), .ZN(n953) );
  NOR2_X1 U1050 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1051 ( .A(KEYINPUT53), .B(n955), .ZN(n956) );
  NOR2_X1 U1052 ( .A1(n957), .A2(n956), .ZN(n960) );
  XOR2_X1 U1053 ( .A(G2084), .B(G34), .Z(n958) );
  XNOR2_X1 U1054 ( .A(KEYINPUT54), .B(n958), .ZN(n959) );
  NAND2_X1 U1055 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1056 ( .A(n962), .B(n961), .ZN(n964) );
  INV_X1 U1057 ( .A(G29), .ZN(n963) );
  NAND2_X1 U1058 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1059 ( .A1(G11), .A2(n965), .ZN(n1020) );
  XNOR2_X1 U1060 ( .A(G16), .B(KEYINPUT56), .ZN(n989) );
  XNOR2_X1 U1061 ( .A(G1966), .B(G168), .ZN(n967) );
  NAND2_X1 U1062 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1063 ( .A(n968), .B(KEYINPUT57), .ZN(n987) );
  NAND2_X1 U1064 ( .A1(G1971), .A2(G303), .ZN(n969) );
  NAND2_X1 U1065 ( .A1(n970), .A2(n969), .ZN(n975) );
  XNOR2_X1 U1066 ( .A(n971), .B(G1956), .ZN(n973) );
  NAND2_X1 U1067 ( .A1(n973), .A2(n972), .ZN(n974) );
  NOR2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n980) );
  XNOR2_X1 U1069 ( .A(G1348), .B(n976), .ZN(n977) );
  NOR2_X1 U1070 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1071 ( .A1(n980), .A2(n979), .ZN(n985) );
  XOR2_X1 U1072 ( .A(n981), .B(G1341), .Z(n983) );
  XNOR2_X1 U1073 ( .A(G171), .B(G1961), .ZN(n982) );
  NAND2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n984) );
  NOR2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1076 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1077 ( .A1(n989), .A2(n988), .ZN(n1018) );
  INV_X1 U1078 ( .A(G16), .ZN(n1016) );
  XOR2_X1 U1079 ( .A(G1986), .B(G24), .Z(n992) );
  XNOR2_X1 U1080 ( .A(G22), .B(KEYINPUT127), .ZN(n990) );
  XNOR2_X1 U1081 ( .A(n990), .B(G1971), .ZN(n991) );
  NAND2_X1 U1082 ( .A1(n992), .A2(n991), .ZN(n994) );
  XNOR2_X1 U1083 ( .A(G23), .B(G1976), .ZN(n993) );
  NOR2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n995) );
  XOR2_X1 U1085 ( .A(KEYINPUT58), .B(n995), .Z(n1013) );
  XOR2_X1 U1086 ( .A(G1961), .B(G5), .Z(n1008) );
  XNOR2_X1 U1087 ( .A(G20), .B(n996), .ZN(n1003) );
  XOR2_X1 U1088 ( .A(KEYINPUT125), .B(G4), .Z(n998) );
  XNOR2_X1 U1089 ( .A(G1348), .B(KEYINPUT59), .ZN(n997) );
  XNOR2_X1 U1090 ( .A(n998), .B(n997), .ZN(n999) );
  XOR2_X1 U1091 ( .A(KEYINPUT124), .B(n999), .Z(n1001) );
  XNOR2_X1 U1092 ( .A(G1981), .B(G6), .ZN(n1000) );
  NOR2_X1 U1093 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1005) );
  XNOR2_X1 U1095 ( .A(G19), .B(G1341), .ZN(n1004) );
  NOR2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1097 ( .A(KEYINPUT60), .B(n1006), .ZN(n1007) );
  NAND2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1010) );
  XNOR2_X1 U1099 ( .A(G21), .B(G1966), .ZN(n1009) );
  NOR2_X1 U1100 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XOR2_X1 U1101 ( .A(KEYINPUT126), .B(n1011), .Z(n1012) );
  NOR2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1103 ( .A(KEYINPUT61), .B(n1014), .ZN(n1015) );
  NAND2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1107 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1108 ( .A(KEYINPUT62), .B(n1023), .Z(G311) );
  INV_X1 U1109 ( .A(G311), .ZN(G150) );
endmodule

