

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778;

  XNOR2_X1 U373 ( .A(n590), .B(n589), .ZN(n594) );
  OR2_X1 U374 ( .A1(n584), .A2(n638), .ZN(n589) );
  XNOR2_X1 U375 ( .A(n652), .B(KEYINPUT6), .ZN(n607) );
  BUF_X1 U376 ( .A(n550), .Z(n652) );
  XNOR2_X1 U377 ( .A(n433), .B(n514), .ZN(n550) );
  OR2_X1 U378 ( .A1(n705), .A2(G902), .ZN(n433) );
  NOR2_X1 U379 ( .A1(n750), .A2(G902), .ZN(n501) );
  BUF_X1 U380 ( .A(G107), .Z(n377) );
  BUF_X1 U381 ( .A(G146), .Z(n425) );
  XNOR2_X1 U382 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n353) );
  AND2_X2 U383 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X2 U384 ( .A(n583), .B(KEYINPUT71), .ZN(n606) );
  XNOR2_X2 U385 ( .A(n572), .B(KEYINPUT45), .ZN(n573) );
  XNOR2_X2 U386 ( .A(n631), .B(KEYINPUT75), .ZN(n685) );
  XNOR2_X2 U387 ( .A(G902), .B(KEYINPUT15), .ZN(n680) );
  AND2_X2 U388 ( .A1(n566), .A2(KEYINPUT34), .ZN(n417) );
  XNOR2_X2 U389 ( .A(n351), .B(KEYINPUT35), .ZN(n704) );
  NAND2_X1 U390 ( .A1(n448), .A2(n447), .ZN(n351) );
  XNOR2_X1 U391 ( .A(n354), .B(n353), .ZN(n352) );
  NOR2_X1 U392 ( .A1(G953), .A2(G237), .ZN(n520) );
  XNOR2_X1 U393 ( .A(n352), .B(n454), .ZN(n356) );
  XNOR2_X1 U394 ( .A(n557), .B(KEYINPUT32), .ZN(n701) );
  BUF_X1 U395 ( .A(G143), .Z(n429) );
  XNOR2_X2 U396 ( .A(n548), .B(n547), .ZN(n556) );
  XNOR2_X2 U397 ( .A(G104), .B(G107), .ZN(n368) );
  NOR2_X1 U398 ( .A1(n777), .A2(n778), .ZN(n428) );
  NOR2_X1 U399 ( .A1(n560), .A2(n607), .ZN(n362) );
  XNOR2_X1 U400 ( .A(n550), .B(n549), .ZN(n584) );
  NOR2_X1 U401 ( .A1(n612), .A2(n388), .ZN(n614) );
  INV_X1 U402 ( .A(n600), .ZN(n635) );
  INV_X1 U403 ( .A(G469), .ZN(n359) );
  INV_X2 U404 ( .A(G146), .ZN(n446) );
  INV_X1 U405 ( .A(KEYINPUT3), .ZN(n373) );
  AND2_X1 U406 ( .A1(n406), .A2(n407), .ZN(n405) );
  AND2_X1 U407 ( .A1(n404), .A2(n402), .ZN(n401) );
  XNOR2_X1 U408 ( .A(n596), .B(n595), .ZN(n620) );
  AND2_X1 U409 ( .A1(n594), .A2(n397), .ZN(n596) );
  XNOR2_X1 U410 ( .A(KEYINPUT107), .B(n610), .ZN(n621) );
  NOR2_X1 U411 ( .A1(n435), .A2(n605), .ZN(n725) );
  XNOR2_X1 U412 ( .A(n362), .B(KEYINPUT33), .ZN(n668) );
  NOR2_X1 U413 ( .A1(n568), .A2(n543), .ZN(n464) );
  XNOR2_X1 U414 ( .A(n380), .B(n381), .ZN(n746) );
  XNOR2_X1 U415 ( .A(n485), .B(n425), .ZN(n372) );
  XNOR2_X1 U416 ( .A(n369), .B(n368), .ZN(n383) );
  XOR2_X2 U417 ( .A(KEYINPUT11), .B(KEYINPUT98), .Z(n518) );
  INV_X2 U418 ( .A(G146), .ZN(n355) );
  INV_X1 U419 ( .A(KEYINPUT46), .ZN(n427) );
  INV_X1 U420 ( .A(G953), .ZN(n490) );
  NAND2_X1 U421 ( .A1(n367), .A2(n366), .ZN(n365) );
  XNOR2_X2 U422 ( .A(n355), .B(G125), .ZN(n354) );
  XNOR2_X2 U423 ( .A(n486), .B(n356), .ZN(n364) );
  XNOR2_X2 U424 ( .A(n535), .B(KEYINPUT4), .ZN(n486) );
  XNOR2_X2 U425 ( .A(n357), .B(n467), .ZN(n535) );
  XNOR2_X2 U426 ( .A(G143), .B(KEYINPUT65), .ZN(n357) );
  NAND2_X1 U427 ( .A1(n358), .A2(n680), .ZN(n363) );
  XNOR2_X1 U428 ( .A(n358), .B(n695), .ZN(n696) );
  XNOR2_X2 U429 ( .A(n364), .B(n760), .ZN(n358) );
  XNOR2_X2 U430 ( .A(n360), .B(n359), .ZN(n586) );
  OR2_X2 U431 ( .A1(n741), .A2(G902), .ZN(n360) );
  XNOR2_X1 U432 ( .A(n361), .B(n487), .ZN(n741) );
  XNOR2_X1 U433 ( .A(n382), .B(n425), .ZN(n361) );
  NAND2_X1 U434 ( .A1(n668), .A2(KEYINPUT34), .ZN(n416) );
  OR2_X2 U435 ( .A1(n646), .A2(n645), .ZN(n560) );
  XNOR2_X2 U436 ( .A(n363), .B(n391), .ZN(n603) );
  XNOR2_X2 U437 ( .A(n365), .B(n466), .ZN(n760) );
  NAND2_X1 U438 ( .A1(n414), .A2(n511), .ZN(n366) );
  NAND2_X1 U439 ( .A1(n384), .A2(n383), .ZN(n367) );
  INV_X1 U440 ( .A(n383), .ZN(n414) );
  XNOR2_X2 U441 ( .A(G101), .B(G110), .ZN(n369) );
  NAND2_X1 U442 ( .A1(n370), .A2(n445), .ZN(n441) );
  OR2_X1 U443 ( .A1(n386), .A2(n444), .ZN(n370) );
  XNOR2_X1 U444 ( .A(n486), .B(n372), .ZN(n456) );
  XNOR2_X2 U445 ( .A(n374), .B(n373), .ZN(n511) );
  XNOR2_X2 U446 ( .A(G119), .B(G113), .ZN(n374) );
  BUF_X1 U447 ( .A(n418), .Z(n375) );
  BUF_X1 U448 ( .A(n414), .Z(n376) );
  XNOR2_X1 U449 ( .A(n446), .B(G125), .ZN(n378) );
  BUF_X1 U450 ( .A(n603), .Z(n379) );
  XNOR2_X1 U451 ( .A(n540), .B(n539), .ZN(n380) );
  AND2_X1 U452 ( .A1(G217), .A2(n541), .ZN(n381) );
  XNOR2_X1 U453 ( .A(n486), .B(n485), .ZN(n382) );
  AND2_X1 U454 ( .A1(n460), .A2(n625), .ZN(n421) );
  INV_X1 U455 ( .A(n511), .ZN(n384) );
  INV_X1 U456 ( .A(n597), .ZN(n385) );
  INV_X1 U457 ( .A(n385), .ZN(n386) );
  BUF_X1 U458 ( .A(n704), .Z(n387) );
  BUF_X1 U459 ( .A(n611), .Z(n388) );
  NOR2_X1 U460 ( .A1(n725), .A2(n403), .ZN(n402) );
  NOR2_X1 U461 ( .A1(KEYINPUT82), .A2(KEYINPUT47), .ZN(n403) );
  NAND2_X1 U462 ( .A1(n405), .A2(n401), .ZN(n438) );
  INV_X1 U463 ( .A(KEYINPUT10), .ZN(n494) );
  XOR2_X1 U464 ( .A(KEYINPUT12), .B(KEYINPUT99), .Z(n522) );
  XNOR2_X1 U465 ( .A(n429), .B(G131), .ZN(n526) );
  XOR2_X1 U466 ( .A(G137), .B(G140), .Z(n495) );
  NAND2_X1 U467 ( .A1(n490), .A2(G224), .ZN(n455) );
  NOR2_X2 U468 ( .A1(n420), .A2(n419), .ZN(n628) );
  XNOR2_X1 U469 ( .A(G119), .B(G128), .ZN(n488) );
  XNOR2_X1 U470 ( .A(KEYINPUT76), .B(KEYINPUT24), .ZN(n462) );
  XNOR2_X1 U471 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U472 ( .A(KEYINPUT93), .B(KEYINPUT25), .ZN(n498) );
  BUF_X1 U473 ( .A(n490), .Z(n769) );
  AND2_X1 U474 ( .A1(n633), .A2(n632), .ZN(n673) );
  INV_X1 U475 ( .A(KEYINPUT74), .ZN(n459) );
  XNOR2_X1 U476 ( .A(KEYINPUT101), .B(KEYINPUT100), .ZN(n517) );
  XOR2_X1 U477 ( .A(G116), .B(KEYINPUT95), .Z(n506) );
  INV_X1 U478 ( .A(KEYINPUT5), .ZN(n507) );
  XNOR2_X1 U479 ( .A(G137), .B(G101), .ZN(n508) );
  XOR2_X1 U480 ( .A(G116), .B(G122), .Z(n536) );
  INV_X1 U481 ( .A(G237), .ZN(n468) );
  NAND2_X1 U482 ( .A1(n389), .A2(KEYINPUT79), .ZN(n439) );
  INV_X1 U483 ( .A(G902), .ZN(n530) );
  XNOR2_X1 U484 ( .A(n586), .B(KEYINPUT1), .ZN(n646) );
  XOR2_X1 U485 ( .A(G140), .B(G122), .Z(n527) );
  XNOR2_X1 U486 ( .A(G134), .B(G131), .ZN(n485) );
  XNOR2_X1 U487 ( .A(n455), .B(KEYINPUT77), .ZN(n454) );
  BUF_X1 U488 ( .A(n646), .Z(n430) );
  XNOR2_X1 U489 ( .A(n707), .B(n706), .ZN(n708) );
  XNOR2_X1 U490 ( .A(n489), .B(n462), .ZN(n493) );
  XOR2_X1 U491 ( .A(KEYINPUT59), .B(n687), .Z(n688) );
  XNOR2_X1 U492 ( .A(n690), .B(KEYINPUT89), .ZN(n744) );
  XNOR2_X1 U493 ( .A(n434), .B(n399), .ZN(n777) );
  INV_X1 U494 ( .A(n656), .ZN(n432) );
  NOR2_X1 U495 ( .A1(n673), .A2(n672), .ZN(n674) );
  OR2_X1 U496 ( .A1(n386), .A2(n586), .ZN(n389) );
  XOR2_X1 U497 ( .A(KEYINPUT23), .B(G110), .Z(n390) );
  AND2_X1 U498 ( .A1(n469), .A2(G210), .ZN(n391) );
  XNOR2_X1 U499 ( .A(n604), .B(KEYINPUT78), .ZN(n392) );
  NOR2_X1 U500 ( .A1(n413), .A2(KEYINPUT2), .ZN(n393) );
  AND2_X1 U501 ( .A1(n635), .A2(n408), .ZN(n394) );
  AND2_X1 U502 ( .A1(n607), .A2(n559), .ZN(n395) );
  AND2_X1 U503 ( .A1(n464), .A2(n545), .ZN(n396) );
  AND2_X1 U504 ( .A1(n593), .A2(n436), .ZN(n397) );
  AND2_X1 U505 ( .A1(n584), .A2(n430), .ZN(n398) );
  XNOR2_X1 U506 ( .A(KEYINPUT109), .B(KEYINPUT40), .ZN(n399) );
  AND2_X1 U507 ( .A1(KEYINPUT82), .A2(KEYINPUT47), .ZN(n400) );
  NAND2_X1 U508 ( .A1(n721), .A2(n635), .ZN(n409) );
  NAND2_X1 U509 ( .A1(n721), .A2(n394), .ZN(n407) );
  NAND2_X1 U510 ( .A1(n601), .A2(n602), .ZN(n404) );
  NAND2_X1 U511 ( .A1(n409), .A2(n400), .ZN(n406) );
  INV_X1 U512 ( .A(KEYINPUT47), .ZN(n408) );
  BUF_X1 U513 ( .A(n382), .Z(n410) );
  XNOR2_X1 U514 ( .A(n418), .B(KEYINPUT91), .ZN(n566) );
  NOR2_X2 U515 ( .A1(n568), .A2(n567), .ZN(n722) );
  XNOR2_X2 U516 ( .A(G478), .B(n542), .ZN(n567) );
  NOR2_X2 U517 ( .A1(n430), .A2(n615), .ZN(n735) );
  NOR2_X1 U518 ( .A1(n618), .A2(KEYINPUT48), .ZN(n423) );
  XNOR2_X1 U519 ( .A(n428), .B(n427), .ZN(n618) );
  NAND2_X1 U520 ( .A1(n440), .A2(n439), .ZN(n411) );
  NAND2_X1 U521 ( .A1(n440), .A2(n439), .ZN(n721) );
  BUF_X1 U522 ( .A(n431), .Z(n412) );
  NAND2_X1 U523 ( .A1(n679), .A2(n413), .ZN(n426) );
  XNOR2_X1 U524 ( .A(n413), .B(n767), .ZN(n768) );
  XNOR2_X2 U525 ( .A(n628), .B(KEYINPUT86), .ZN(n413) );
  XNOR2_X1 U526 ( .A(n484), .B(n376), .ZN(n487) );
  NOR2_X1 U527 ( .A1(n417), .A2(n415), .ZN(n448) );
  NAND2_X1 U528 ( .A1(n416), .A2(n392), .ZN(n415) );
  XNOR2_X2 U529 ( .A(n451), .B(KEYINPUT0), .ZN(n418) );
  NAND2_X1 U530 ( .A1(n418), .A2(n396), .ZN(n548) );
  NAND2_X1 U531 ( .A1(n432), .A2(n375), .ZN(n562) );
  XNOR2_X1 U532 ( .A(n378), .B(n494), .ZN(n515) );
  AND2_X1 U533 ( .A1(n461), .A2(KEYINPUT48), .ZN(n419) );
  NAND2_X1 U534 ( .A1(n422), .A2(n421), .ZN(n420) );
  NAND2_X1 U535 ( .A1(n424), .A2(n423), .ZN(n422) );
  INV_X1 U536 ( .A(n461), .ZN(n424) );
  NAND2_X1 U537 ( .A1(n552), .A2(n582), .ZN(n431) );
  NAND2_X1 U538 ( .A1(n426), .A2(n682), .ZN(n684) );
  NAND2_X1 U539 ( .A1(n437), .A2(n616), .ZN(n617) );
  XNOR2_X1 U540 ( .A(n617), .B(KEYINPUT70), .ZN(n461) );
  XNOR2_X1 U541 ( .A(n438), .B(n459), .ZN(n437) );
  XNOR2_X1 U542 ( .A(n452), .B(KEYINPUT67), .ZN(n552) );
  NOR2_X2 U543 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U544 ( .A1(n620), .A2(n727), .ZN(n434) );
  NOR2_X2 U545 ( .A1(n677), .A2(n680), .ZN(n678) );
  XNOR2_X2 U546 ( .A(n574), .B(n573), .ZN(n677) );
  NAND2_X1 U547 ( .A1(n431), .A2(n701), .ZN(n558) );
  XNOR2_X1 U548 ( .A(n412), .B(n703), .ZN(G12) );
  NAND2_X1 U549 ( .A1(n594), .A2(n593), .ZN(n435) );
  INV_X1 U550 ( .A(n639), .ZN(n436) );
  XNOR2_X1 U551 ( .A(n410), .B(n766), .ZN(n771) );
  NAND2_X1 U552 ( .A1(n442), .A2(n441), .ZN(n440) );
  NAND2_X1 U553 ( .A1(n443), .A2(n599), .ZN(n442) );
  INV_X1 U554 ( .A(n445), .ZN(n443) );
  XNOR2_X2 U555 ( .A(n585), .B(KEYINPUT28), .ZN(n445) );
  NAND2_X1 U556 ( .A1(n445), .A2(n587), .ZN(n598) );
  NAND2_X1 U557 ( .A1(n587), .A2(n599), .ZN(n444) );
  NAND2_X1 U558 ( .A1(n450), .A2(n449), .ZN(n447) );
  INV_X1 U559 ( .A(n668), .ZN(n449) );
  NOR2_X1 U560 ( .A1(n566), .A2(KEYINPUT34), .ZN(n450) );
  NOR2_X2 U561 ( .A1(n584), .A2(n606), .ZN(n585) );
  NOR2_X2 U562 ( .A1(n597), .A2(n481), .ZN(n451) );
  XNOR2_X2 U563 ( .A(n611), .B(n474), .ZN(n597) );
  XNOR2_X2 U564 ( .A(n453), .B(n473), .ZN(n611) );
  AND2_X1 U565 ( .A1(n556), .A2(n430), .ZN(n551) );
  NAND2_X1 U566 ( .A1(n556), .A2(n398), .ZN(n452) );
  NAND2_X1 U567 ( .A1(n603), .A2(n472), .ZN(n453) );
  NAND2_X1 U568 ( .A1(n551), .A2(n395), .ZN(n713) );
  XNOR2_X1 U569 ( .A(n456), .B(n513), .ZN(n705) );
  NAND2_X1 U570 ( .A1(n457), .A2(n571), .ZN(n574) );
  XNOR2_X1 U571 ( .A(n458), .B(KEYINPUT44), .ZN(n457) );
  NOR2_X2 U572 ( .A1(n558), .A2(n704), .ZN(n458) );
  NAND2_X1 U573 ( .A1(n618), .A2(KEYINPUT48), .ZN(n460) );
  BUF_X1 U574 ( .A(n677), .Z(n629) );
  XOR2_X1 U575 ( .A(n524), .B(n523), .Z(n463) );
  XOR2_X1 U576 ( .A(n623), .B(KEYINPUT43), .Z(n465) );
  XNOR2_X1 U577 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U578 ( .A(n510), .B(n509), .ZN(n512) );
  INV_X1 U579 ( .A(n638), .ZN(n472) );
  INV_X1 U580 ( .A(KEYINPUT66), .ZN(n683) );
  BUF_X1 U581 ( .A(n705), .Z(n707) );
  XNOR2_X1 U582 ( .A(n493), .B(n492), .ZN(n496) );
  INV_X1 U583 ( .A(KEYINPUT36), .ZN(n613) );
  INV_X1 U584 ( .A(KEYINPUT79), .ZN(n599) );
  XNOR2_X1 U585 ( .A(n741), .B(n740), .ZN(n742) );
  BUF_X1 U586 ( .A(n411), .Z(n726) );
  XNOR2_X1 U587 ( .A(n743), .B(n742), .ZN(n745) );
  XNOR2_X1 U588 ( .A(n676), .B(n675), .ZN(G75) );
  XNOR2_X1 U589 ( .A(n536), .B(KEYINPUT16), .ZN(n466) );
  INV_X1 U590 ( .A(G128), .ZN(n467) );
  NAND2_X1 U591 ( .A1(n530), .A2(n468), .ZN(n469) );
  NAND2_X1 U592 ( .A1(n469), .A2(G214), .ZN(n471) );
  INV_X1 U593 ( .A(KEYINPUT90), .ZN(n470) );
  XNOR2_X1 U594 ( .A(n471), .B(n470), .ZN(n638) );
  INV_X1 U595 ( .A(KEYINPUT87), .ZN(n473) );
  XNOR2_X1 U596 ( .A(KEYINPUT69), .B(KEYINPUT19), .ZN(n474) );
  NAND2_X1 U597 ( .A1(G234), .A2(G237), .ZN(n475) );
  XNOR2_X1 U598 ( .A(n475), .B(KEYINPUT14), .ZN(n634) );
  INV_X1 U599 ( .A(G952), .ZN(n476) );
  NAND2_X1 U600 ( .A1(n769), .A2(n476), .ZN(n478) );
  OR2_X1 U601 ( .A1(n769), .A2(G902), .ZN(n477) );
  AND2_X1 U602 ( .A1(n478), .A2(n477), .ZN(n479) );
  AND2_X1 U603 ( .A1(n634), .A2(n479), .ZN(n580) );
  NAND2_X1 U604 ( .A1(G953), .A2(G898), .ZN(n480) );
  NAND2_X1 U605 ( .A1(n580), .A2(n480), .ZN(n481) );
  XOR2_X1 U606 ( .A(n495), .B(KEYINPUT92), .Z(n483) );
  NAND2_X1 U607 ( .A1(G227), .A2(n769), .ZN(n482) );
  XNOR2_X1 U608 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U609 ( .A(n390), .B(n488), .ZN(n489) );
  NAND2_X1 U610 ( .A1(G234), .A2(n490), .ZN(n491) );
  XOR2_X1 U611 ( .A(KEYINPUT8), .B(n491), .Z(n541) );
  NAND2_X1 U612 ( .A1(G221), .A2(n541), .ZN(n492) );
  XNOR2_X1 U613 ( .A(n495), .B(n515), .ZN(n766) );
  XNOR2_X1 U614 ( .A(n496), .B(n766), .ZN(n750) );
  NAND2_X1 U615 ( .A1(G234), .A2(n680), .ZN(n497) );
  XNOR2_X1 U616 ( .A(KEYINPUT20), .B(n497), .ZN(n502) );
  NAND2_X1 U617 ( .A1(n502), .A2(G217), .ZN(n499) );
  XNOR2_X2 U618 ( .A(n501), .B(n500), .ZN(n582) );
  NAND2_X1 U619 ( .A1(n502), .A2(G221), .ZN(n503) );
  XNOR2_X1 U620 ( .A(n503), .B(KEYINPUT21), .ZN(n648) );
  XNOR2_X1 U621 ( .A(n648), .B(KEYINPUT94), .ZN(n544) );
  NOR2_X1 U622 ( .A1(n582), .A2(n544), .ZN(n504) );
  INV_X1 U623 ( .A(n504), .ZN(n645) );
  NAND2_X1 U624 ( .A1(n520), .A2(G210), .ZN(n505) );
  XNOR2_X1 U625 ( .A(n506), .B(n505), .ZN(n510) );
  XNOR2_X1 U626 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U627 ( .A(G472), .B(KEYINPUT72), .ZN(n514) );
  XNOR2_X1 U628 ( .A(n515), .B(G104), .ZN(n516) );
  XNOR2_X1 U629 ( .A(n516), .B(KEYINPUT97), .ZN(n525) );
  XNOR2_X1 U630 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U631 ( .A(G113), .B(n519), .ZN(n524) );
  NAND2_X1 U632 ( .A1(G214), .A2(n520), .ZN(n521) );
  XNOR2_X1 U633 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U634 ( .A(n525), .B(n463), .ZN(n529) );
  XOR2_X1 U635 ( .A(n527), .B(n526), .Z(n528) );
  XNOR2_X1 U636 ( .A(n529), .B(n528), .ZN(n687) );
  NAND2_X1 U637 ( .A1(n687), .A2(n530), .ZN(n532) );
  XOR2_X1 U638 ( .A(KEYINPUT13), .B(G475), .Z(n531) );
  XNOR2_X2 U639 ( .A(n532), .B(n531), .ZN(n568) );
  XOR2_X1 U640 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n534) );
  XNOR2_X1 U641 ( .A(G134), .B(KEYINPUT7), .ZN(n533) );
  XNOR2_X1 U642 ( .A(n534), .B(n533), .ZN(n540) );
  XOR2_X1 U643 ( .A(n535), .B(n377), .Z(n538) );
  XOR2_X1 U644 ( .A(KEYINPUT9), .B(n536), .Z(n537) );
  XNOR2_X1 U645 ( .A(n538), .B(n537), .ZN(n539) );
  NOR2_X1 U646 ( .A1(G902), .A2(n746), .ZN(n542) );
  INV_X1 U647 ( .A(n567), .ZN(n543) );
  AND2_X1 U648 ( .A1(n568), .A2(n543), .ZN(n604) );
  INV_X1 U649 ( .A(n544), .ZN(n545) );
  XNOR2_X1 U650 ( .A(KEYINPUT73), .B(KEYINPUT22), .ZN(n546) );
  XNOR2_X1 U651 ( .A(n546), .B(KEYINPUT68), .ZN(n547) );
  INV_X1 U652 ( .A(KEYINPUT106), .ZN(n549) );
  INV_X1 U653 ( .A(KEYINPUT105), .ZN(n553) );
  XNOR2_X1 U654 ( .A(n582), .B(n553), .ZN(n649) );
  INV_X1 U655 ( .A(n649), .ZN(n559) );
  NOR2_X1 U656 ( .A1(n430), .A2(n559), .ZN(n554) );
  AND2_X1 U657 ( .A1(n554), .A2(n607), .ZN(n555) );
  NAND2_X1 U658 ( .A1(n556), .A2(n555), .ZN(n557) );
  INV_X1 U659 ( .A(n652), .ZN(n563) );
  OR2_X1 U660 ( .A1(n560), .A2(n563), .ZN(n656) );
  XOR2_X1 U661 ( .A(KEYINPUT96), .B(KEYINPUT31), .Z(n561) );
  XNOR2_X1 U662 ( .A(n562), .B(n561), .ZN(n733) );
  OR2_X1 U663 ( .A1(n586), .A2(n645), .ZN(n591) );
  INV_X1 U664 ( .A(n591), .ZN(n564) );
  NAND2_X1 U665 ( .A1(n564), .A2(n563), .ZN(n565) );
  OR2_X1 U666 ( .A1(n566), .A2(n565), .ZN(n715) );
  NAND2_X1 U667 ( .A1(n733), .A2(n715), .ZN(n569) );
  XNOR2_X1 U668 ( .A(KEYINPUT104), .B(n722), .ZN(n619) );
  NAND2_X1 U669 ( .A1(n568), .A2(n567), .ZN(n730) );
  INV_X1 U670 ( .A(n730), .ZN(n727) );
  NOR2_X1 U671 ( .A1(n619), .A2(n727), .ZN(n600) );
  NAND2_X1 U672 ( .A1(n569), .A2(n635), .ZN(n570) );
  AND2_X1 U673 ( .A1(n713), .A2(n570), .ZN(n571) );
  INV_X1 U674 ( .A(KEYINPUT64), .ZN(n572) );
  INV_X1 U675 ( .A(KEYINPUT2), .ZN(n575) );
  NAND2_X1 U676 ( .A1(n629), .A2(n575), .ZN(n576) );
  XNOR2_X1 U677 ( .A(n576), .B(KEYINPUT83), .ZN(n626) );
  INV_X1 U678 ( .A(n379), .ZN(n624) );
  INV_X1 U679 ( .A(KEYINPUT38), .ZN(n577) );
  XNOR2_X1 U680 ( .A(n624), .B(n577), .ZN(n639) );
  NOR2_X1 U681 ( .A1(n639), .A2(n638), .ZN(n636) );
  NAND2_X1 U682 ( .A1(n464), .A2(n636), .ZN(n578) );
  XOR2_X1 U683 ( .A(KEYINPUT41), .B(n578), .Z(n667) );
  NAND2_X1 U684 ( .A1(G953), .A2(G900), .ZN(n579) );
  NAND2_X1 U685 ( .A1(n580), .A2(n579), .ZN(n592) );
  NOR2_X1 U686 ( .A1(n648), .A2(n592), .ZN(n581) );
  INV_X1 U687 ( .A(n586), .ZN(n587) );
  NOR2_X1 U688 ( .A1(n667), .A2(n598), .ZN(n588) );
  XNOR2_X1 U689 ( .A(n588), .B(KEYINPUT42), .ZN(n778) );
  XOR2_X1 U690 ( .A(KEYINPUT108), .B(KEYINPUT30), .Z(n590) );
  INV_X1 U691 ( .A(KEYINPUT39), .ZN(n595) );
  INV_X1 U692 ( .A(KEYINPUT82), .ZN(n602) );
  NAND2_X1 U693 ( .A1(n411), .A2(n600), .ZN(n601) );
  NAND2_X1 U694 ( .A1(n604), .A2(n379), .ZN(n605) );
  INV_X1 U695 ( .A(n606), .ZN(n609) );
  NOR2_X1 U696 ( .A1(n730), .A2(n607), .ZN(n608) );
  NAND2_X1 U697 ( .A1(n609), .A2(n608), .ZN(n610) );
  INV_X1 U698 ( .A(n621), .ZN(n612) );
  XNOR2_X1 U699 ( .A(n614), .B(n613), .ZN(n615) );
  INV_X1 U700 ( .A(n735), .ZN(n616) );
  NAND2_X1 U701 ( .A1(n620), .A2(n619), .ZN(n738) );
  NAND2_X1 U702 ( .A1(n430), .A2(n621), .ZN(n622) );
  NOR2_X1 U703 ( .A1(n638), .A2(n622), .ZN(n623) );
  NAND2_X1 U704 ( .A1(n465), .A2(n624), .ZN(n702) );
  AND2_X1 U705 ( .A1(n738), .A2(n702), .ZN(n625) );
  NOR2_X1 U706 ( .A1(n626), .A2(n393), .ZN(n627) );
  XNOR2_X1 U707 ( .A(n627), .B(KEYINPUT80), .ZN(n633) );
  AND2_X1 U708 ( .A1(n628), .A2(KEYINPUT2), .ZN(n630) );
  INV_X1 U709 ( .A(n629), .ZN(n756) );
  NAND2_X1 U710 ( .A1(n630), .A2(n756), .ZN(n631) );
  INV_X1 U711 ( .A(n685), .ZN(n632) );
  NAND2_X1 U712 ( .A1(G952), .A2(n634), .ZN(n666) );
  NAND2_X1 U713 ( .A1(n636), .A2(n635), .ZN(n637) );
  XOR2_X1 U714 ( .A(KEYINPUT119), .B(n637), .Z(n643) );
  NAND2_X1 U715 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U716 ( .A(KEYINPUT118), .B(n640), .ZN(n641) );
  NAND2_X1 U717 ( .A1(n641), .A2(n464), .ZN(n642) );
  NAND2_X1 U718 ( .A1(n643), .A2(n642), .ZN(n644) );
  NAND2_X1 U719 ( .A1(n644), .A2(n449), .ZN(n662) );
  NAND2_X1 U720 ( .A1(n430), .A2(n645), .ZN(n647) );
  XNOR2_X1 U721 ( .A(KEYINPUT50), .B(n647), .ZN(n654) );
  NAND2_X1 U722 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U723 ( .A(KEYINPUT49), .B(n650), .ZN(n651) );
  NOR2_X1 U724 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U725 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U726 ( .A(n655), .B(KEYINPUT116), .ZN(n657) );
  NAND2_X1 U727 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U728 ( .A(KEYINPUT51), .B(n658), .ZN(n659) );
  NOR2_X1 U729 ( .A1(n667), .A2(n659), .ZN(n660) );
  XNOR2_X1 U730 ( .A(KEYINPUT117), .B(n660), .ZN(n661) );
  NAND2_X1 U731 ( .A1(n662), .A2(n661), .ZN(n663) );
  XOR2_X1 U732 ( .A(KEYINPUT52), .B(n663), .Z(n664) );
  XNOR2_X1 U733 ( .A(KEYINPUT120), .B(n664), .ZN(n665) );
  NOR2_X1 U734 ( .A1(n666), .A2(n665), .ZN(n670) );
  NOR2_X1 U735 ( .A1(n668), .A2(n667), .ZN(n669) );
  NOR2_X1 U736 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U737 ( .A(n671), .B(KEYINPUT121), .ZN(n672) );
  NAND2_X1 U738 ( .A1(n769), .A2(n674), .ZN(n676) );
  INV_X1 U739 ( .A(KEYINPUT53), .ZN(n675) );
  XNOR2_X1 U740 ( .A(n678), .B(KEYINPUT84), .ZN(n679) );
  XNOR2_X1 U741 ( .A(n680), .B(KEYINPUT85), .ZN(n681) );
  NAND2_X1 U742 ( .A1(n681), .A2(KEYINPUT2), .ZN(n682) );
  XNOR2_X1 U743 ( .A(n684), .B(n683), .ZN(n686) );
  NOR2_X2 U744 ( .A1(n686), .A2(n685), .ZN(n739) );
  NAND2_X1 U745 ( .A1(n739), .A2(G475), .ZN(n689) );
  XNOR2_X1 U746 ( .A(n689), .B(n688), .ZN(n691) );
  NOR2_X1 U747 ( .A1(n769), .A2(G952), .ZN(n690) );
  NAND2_X1 U748 ( .A1(n691), .A2(n744), .ZN(n693) );
  INV_X1 U749 ( .A(KEYINPUT60), .ZN(n692) );
  XNOR2_X1 U750 ( .A(n693), .B(n692), .ZN(G60) );
  NAND2_X1 U751 ( .A1(n739), .A2(G210), .ZN(n697) );
  XNOR2_X1 U752 ( .A(KEYINPUT55), .B(KEYINPUT81), .ZN(n694) );
  XNOR2_X1 U753 ( .A(n694), .B(KEYINPUT54), .ZN(n695) );
  XNOR2_X1 U754 ( .A(n697), .B(n696), .ZN(n698) );
  NAND2_X1 U755 ( .A1(n698), .A2(n744), .ZN(n700) );
  INV_X1 U756 ( .A(KEYINPUT56), .ZN(n699) );
  XNOR2_X1 U757 ( .A(n700), .B(n699), .ZN(G51) );
  XNOR2_X1 U758 ( .A(n701), .B(G119), .ZN(G21) );
  XNOR2_X1 U759 ( .A(n702), .B(G140), .ZN(G42) );
  XOR2_X1 U760 ( .A(G110), .B(KEYINPUT113), .Z(n703) );
  XOR2_X1 U761 ( .A(G122), .B(n387), .Z(G24) );
  NAND2_X1 U762 ( .A1(n739), .A2(G472), .ZN(n709) );
  XOR2_X1 U763 ( .A(KEYINPUT110), .B(KEYINPUT62), .Z(n706) );
  XNOR2_X1 U764 ( .A(n709), .B(n708), .ZN(n710) );
  NAND2_X1 U765 ( .A1(n710), .A2(n744), .ZN(n712) );
  XNOR2_X1 U766 ( .A(KEYINPUT88), .B(KEYINPUT63), .ZN(n711) );
  XNOR2_X1 U767 ( .A(n712), .B(n711), .ZN(G57) );
  XNOR2_X1 U768 ( .A(G101), .B(n713), .ZN(G3) );
  NOR2_X1 U769 ( .A1(n730), .A2(n715), .ZN(n714) );
  XOR2_X1 U770 ( .A(G104), .B(n714), .Z(G6) );
  INV_X1 U771 ( .A(n722), .ZN(n732) );
  NOR2_X1 U772 ( .A1(n732), .A2(n715), .ZN(n720) );
  XOR2_X1 U773 ( .A(KEYINPUT112), .B(KEYINPUT27), .Z(n717) );
  XNOR2_X1 U774 ( .A(n377), .B(KEYINPUT26), .ZN(n716) );
  XNOR2_X1 U775 ( .A(n717), .B(n716), .ZN(n718) );
  XNOR2_X1 U776 ( .A(KEYINPUT111), .B(n718), .ZN(n719) );
  XNOR2_X1 U777 ( .A(n720), .B(n719), .ZN(G9) );
  XOR2_X1 U778 ( .A(G128), .B(KEYINPUT29), .Z(n724) );
  NAND2_X1 U779 ( .A1(n726), .A2(n722), .ZN(n723) );
  XNOR2_X1 U780 ( .A(n724), .B(n723), .ZN(G30) );
  XOR2_X1 U781 ( .A(n429), .B(n725), .Z(G45) );
  XNOR2_X1 U782 ( .A(n425), .B(KEYINPUT114), .ZN(n729) );
  NAND2_X1 U783 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U784 ( .A(n729), .B(n728), .ZN(G48) );
  NOR2_X1 U785 ( .A1(n733), .A2(n730), .ZN(n731) );
  XOR2_X1 U786 ( .A(G113), .B(n731), .Z(G15) );
  NOR2_X1 U787 ( .A1(n733), .A2(n732), .ZN(n734) );
  XOR2_X1 U788 ( .A(G116), .B(n734), .Z(G18) );
  XOR2_X1 U789 ( .A(KEYINPUT37), .B(KEYINPUT115), .Z(n737) );
  XNOR2_X1 U790 ( .A(G125), .B(n735), .ZN(n736) );
  XNOR2_X1 U791 ( .A(n737), .B(n736), .ZN(G27) );
  XNOR2_X1 U792 ( .A(G134), .B(n738), .ZN(G36) );
  BUF_X2 U793 ( .A(n739), .Z(n749) );
  NAND2_X1 U794 ( .A1(n749), .A2(G469), .ZN(n743) );
  XOR2_X1 U795 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n740) );
  INV_X1 U796 ( .A(n744), .ZN(n753) );
  NOR2_X1 U797 ( .A1(n745), .A2(n753), .ZN(G54) );
  NAND2_X1 U798 ( .A1(n749), .A2(G478), .ZN(n747) );
  XNOR2_X1 U799 ( .A(n747), .B(n746), .ZN(n748) );
  NOR2_X1 U800 ( .A1(n753), .A2(n748), .ZN(G63) );
  NAND2_X1 U801 ( .A1(n749), .A2(G217), .ZN(n751) );
  XNOR2_X1 U802 ( .A(n751), .B(n750), .ZN(n752) );
  NOR2_X1 U803 ( .A1(n753), .A2(n752), .ZN(G66) );
  NAND2_X1 U804 ( .A1(G953), .A2(G224), .ZN(n754) );
  XNOR2_X1 U805 ( .A(KEYINPUT61), .B(n754), .ZN(n755) );
  NAND2_X1 U806 ( .A1(n755), .A2(G898), .ZN(n759) );
  NAND2_X1 U807 ( .A1(n756), .A2(n769), .ZN(n757) );
  XNOR2_X1 U808 ( .A(n757), .B(KEYINPUT122), .ZN(n758) );
  NAND2_X1 U809 ( .A1(n759), .A2(n758), .ZN(n765) );
  NOR2_X1 U810 ( .A1(G898), .A2(n769), .ZN(n762) );
  XOR2_X1 U811 ( .A(n760), .B(KEYINPUT124), .Z(n761) );
  NOR2_X1 U812 ( .A1(n762), .A2(n761), .ZN(n763) );
  XOR2_X1 U813 ( .A(KEYINPUT123), .B(n763), .Z(n764) );
  XNOR2_X1 U814 ( .A(n765), .B(n764), .ZN(G69) );
  XNOR2_X1 U815 ( .A(n771), .B(KEYINPUT125), .ZN(n767) );
  NAND2_X1 U816 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U817 ( .A(n770), .B(KEYINPUT126), .ZN(n775) );
  XNOR2_X1 U818 ( .A(G227), .B(n771), .ZN(n772) );
  NAND2_X1 U819 ( .A1(n772), .A2(G900), .ZN(n773) );
  NAND2_X1 U820 ( .A1(n773), .A2(G953), .ZN(n774) );
  NAND2_X1 U821 ( .A1(n775), .A2(n774), .ZN(n776) );
  XOR2_X1 U822 ( .A(KEYINPUT127), .B(n776), .Z(G72) );
  XOR2_X1 U823 ( .A(n777), .B(G131), .Z(G33) );
  XOR2_X1 U824 ( .A(G137), .B(n778), .Z(G39) );
endmodule

