//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 0 0 1 1 1 0 0 1 0 0 1 0 1 1 0 1 1 1 0 1 0 1 0 0 0 1 1 0 0 0 0 0 0 1 1 1 1 0 1 0 1 0 0 0 0 1 1 1 0 0 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:02 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n657, new_n658, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938;
  XNOR2_X1  g000(.A(G116), .B(G119), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XNOR2_X1  g002(.A(KEYINPUT2), .B(G113), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(new_n189), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(new_n187), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT67), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n190), .A2(new_n192), .A3(KEYINPUT67), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  XNOR2_X1  g011(.A(G143), .B(G146), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT1), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n198), .A2(new_n199), .A3(G128), .ZN(new_n200));
  INV_X1    g014(.A(G143), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(KEYINPUT1), .A3(G146), .ZN(new_n202));
  OAI211_X1 g016(.A(new_n200), .B(new_n202), .C1(G128), .C2(new_n198), .ZN(new_n203));
  INV_X1    g017(.A(G134), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G137), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n204), .A2(G137), .ZN(new_n207));
  OAI21_X1  g021(.A(G131), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT11), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n209), .B1(new_n204), .B2(G137), .ZN(new_n210));
  INV_X1    g024(.A(G137), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n211), .A2(KEYINPUT11), .A3(G134), .ZN(new_n212));
  INV_X1    g026(.A(G131), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n210), .A2(new_n212), .A3(new_n213), .A4(new_n205), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT64), .ZN(new_n215));
  AND2_X1   g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n214), .A2(new_n215), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n203), .B(new_n208), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AND2_X1   g032(.A1(new_n197), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n210), .A2(new_n205), .A3(new_n212), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G131), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n221), .B1(new_n216), .B2(new_n217), .ZN(new_n222));
  NAND2_X1  g036(.A1(KEYINPUT0), .A2(G128), .ZN(new_n223));
  OR2_X1    g037(.A1(KEYINPUT0), .A2(G128), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n198), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n198), .A2(new_n223), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n222), .A2(new_n228), .ZN(new_n229));
  AND2_X1   g043(.A1(new_n219), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n230), .A2(KEYINPUT28), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT65), .ZN(new_n232));
  AND2_X1   g046(.A1(new_n220), .A2(G131), .ZN(new_n233));
  AND2_X1   g047(.A1(new_n210), .A2(new_n212), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n234), .A2(KEYINPUT64), .A3(new_n213), .A4(new_n205), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n214), .A2(new_n215), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n233), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n232), .B1(new_n237), .B2(new_n227), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n222), .A2(KEYINPUT65), .A3(new_n228), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n238), .A2(new_n218), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT66), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n241), .B1(new_n237), .B2(new_n227), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n222), .A2(KEYINPUT66), .A3(new_n228), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n240), .A2(new_n193), .B1(new_n244), .B2(new_n219), .ZN(new_n245));
  XOR2_X1   g059(.A(KEYINPUT69), .B(KEYINPUT28), .Z(new_n246));
  OAI21_X1  g060(.A(KEYINPUT70), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n240), .A2(new_n193), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n244), .A2(new_n219), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT70), .ZN(new_n251));
  INV_X1    g065(.A(new_n246), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n250), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n231), .B1(new_n247), .B2(new_n253), .ZN(new_n254));
  NOR2_X1   g068(.A1(G237), .A2(G953), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G210), .ZN(new_n256));
  XOR2_X1   g070(.A(new_n256), .B(G101), .Z(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n258));
  XOR2_X1   g072(.A(new_n257), .B(new_n258), .Z(new_n259));
  OAI21_X1  g073(.A(KEYINPUT71), .B1(new_n254), .B2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n231), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n251), .B1(new_n250), .B2(new_n252), .ZN(new_n262));
  AOI211_X1 g076(.A(KEYINPUT70), .B(new_n246), .C1(new_n248), .C2(new_n249), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n261), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT71), .ZN(new_n265));
  INV_X1    g079(.A(new_n259), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT30), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n238), .A2(new_n239), .A3(new_n268), .A4(new_n218), .ZN(new_n269));
  INV_X1    g083(.A(new_n218), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n270), .B1(new_n242), .B2(new_n243), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n269), .B1(new_n271), .B2(new_n268), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(new_n193), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT68), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT31), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n273), .A2(new_n259), .A3(new_n249), .A4(new_n275), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n274), .A2(KEYINPUT31), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI22_X1  g092(.A1(new_n272), .A2(new_n193), .B1(new_n219), .B2(new_n244), .ZN(new_n279));
  INV_X1    g093(.A(new_n277), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n279), .A2(new_n259), .A3(new_n275), .A4(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n278), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n260), .A2(new_n267), .A3(new_n282), .ZN(new_n283));
  NOR2_X1   g097(.A1(G472), .A2(G902), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(KEYINPUT32), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT32), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n283), .A2(new_n287), .A3(new_n284), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n249), .B1(new_n197), .B2(new_n271), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n231), .B1(new_n289), .B2(KEYINPUT28), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT29), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n266), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(G902), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n291), .B1(new_n264), .B2(new_n266), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n279), .A2(new_n259), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  AOI22_X1  g110(.A1(new_n286), .A2(new_n288), .B1(G472), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(G125), .A2(G140), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  NOR2_X1   g113(.A1(G125), .A2(G140), .ZN(new_n300));
  OAI21_X1  g114(.A(KEYINPUT16), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G125), .ZN(new_n302));
  OR3_X1    g116(.A1(new_n302), .A2(KEYINPUT16), .A3(G140), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n301), .A2(G146), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT73), .ZN(new_n305));
  OR2_X1    g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n301), .A2(new_n303), .ZN(new_n307));
  INV_X1    g121(.A(G146), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n304), .A2(new_n305), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n306), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  XOR2_X1   g125(.A(KEYINPUT24), .B(G110), .Z(new_n312));
  XNOR2_X1  g126(.A(G119), .B(G128), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT23), .ZN(new_n315));
  INV_X1    g129(.A(G119), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n315), .B1(new_n316), .B2(G128), .ZN(new_n317));
  INV_X1    g131(.A(G128), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n318), .A2(KEYINPUT23), .A3(G119), .ZN(new_n319));
  OAI211_X1 g133(.A(new_n317), .B(new_n319), .C1(G119), .C2(new_n318), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G110), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n311), .A2(new_n314), .A3(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n304), .B(KEYINPUT75), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n308), .B1(new_n299), .B2(new_n300), .ZN(new_n324));
  XNOR2_X1  g138(.A(KEYINPUT74), .B(G110), .ZN(new_n325));
  OAI22_X1  g139(.A1(new_n320), .A2(new_n325), .B1(new_n313), .B2(new_n312), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n323), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n322), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT22), .B(G137), .ZN(new_n329));
  INV_X1    g143(.A(G221), .ZN(new_n330));
  INV_X1    g144(.A(G234), .ZN(new_n331));
  NOR3_X1   g145(.A1(new_n330), .A2(new_n331), .A3(G953), .ZN(new_n332));
  XOR2_X1   g146(.A(new_n329), .B(new_n332), .Z(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n328), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n322), .A2(new_n327), .A3(new_n333), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  OR3_X1    g151(.A1(new_n337), .A2(KEYINPUT25), .A3(G902), .ZN(new_n338));
  OAI21_X1  g152(.A(G217), .B1(new_n331), .B2(G902), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n339), .B(KEYINPUT72), .ZN(new_n340));
  OAI21_X1  g154(.A(KEYINPUT25), .B1(new_n337), .B2(G902), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n338), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n337), .ZN(new_n343));
  INV_X1    g157(.A(G902), .ZN(new_n344));
  INV_X1    g158(.A(new_n340), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n347), .B(KEYINPUT76), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n297), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(G104), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n351), .A2(G107), .ZN(new_n352));
  AND2_X1   g166(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n353));
  NOR2_X1   g167(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT78), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n352), .ZN(new_n358));
  INV_X1    g172(.A(G107), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n359), .A2(G104), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n358), .B1(new_n360), .B2(KEYINPUT3), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n352), .B(KEYINPUT78), .C1(new_n354), .C2(new_n353), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n357), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(KEYINPUT79), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT79), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n357), .A2(new_n361), .A3(new_n365), .A4(new_n362), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n364), .A2(G101), .A3(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(KEYINPUT80), .B(G101), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n357), .A2(new_n361), .A3(new_n368), .A4(new_n362), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n367), .A2(KEYINPUT4), .A3(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT4), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n364), .A2(new_n371), .A3(G101), .A4(new_n366), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n370), .A2(new_n228), .A3(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT10), .ZN(new_n374));
  OAI21_X1  g188(.A(G101), .B1(new_n352), .B2(new_n360), .ZN(new_n375));
  AND3_X1   g189(.A1(new_n369), .A2(new_n203), .A3(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT81), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n374), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n369), .A2(new_n203), .A3(new_n375), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n379), .A2(KEYINPUT81), .A3(KEYINPUT10), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  AND3_X1   g195(.A1(new_n373), .A2(new_n237), .A3(new_n381), .ZN(new_n382));
  XNOR2_X1  g196(.A(G110), .B(G140), .ZN(new_n383));
  INV_X1    g197(.A(G227), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n384), .A2(G953), .ZN(new_n385));
  XOR2_X1   g199(.A(new_n383), .B(new_n385), .Z(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(KEYINPUT83), .B1(new_n382), .B2(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n203), .B1(new_n369), .B2(new_n375), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n222), .B1(new_n376), .B2(new_n389), .ZN(new_n390));
  XOR2_X1   g204(.A(new_n390), .B(KEYINPUT12), .Z(new_n391));
  NAND3_X1  g205(.A1(new_n373), .A2(new_n381), .A3(new_n237), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT83), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n392), .A2(new_n393), .A3(new_n386), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n388), .A2(new_n391), .A3(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT84), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n237), .B1(new_n373), .B2(new_n381), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n387), .B1(new_n382), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT85), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OAI211_X1 g215(.A(KEYINPUT85), .B(new_n387), .C1(new_n382), .C2(new_n398), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n388), .A2(KEYINPUT84), .A3(new_n391), .A4(new_n394), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n397), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(G469), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(new_n406), .A3(new_n344), .ZN(new_n407));
  NAND2_X1  g221(.A1(G469), .A2(G902), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n391), .A2(new_n392), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT82), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT82), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n391), .A2(new_n392), .A3(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n410), .A2(new_n387), .A3(new_n412), .ZN(new_n413));
  OR3_X1    g227(.A1(new_n382), .A2(new_n398), .A3(new_n387), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n413), .A2(G469), .A3(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n407), .A2(new_n408), .A3(new_n415), .ZN(new_n416));
  XOR2_X1   g230(.A(KEYINPUT9), .B(G234), .Z(new_n417));
  AOI21_X1  g231(.A(new_n330), .B1(new_n417), .B2(new_n344), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  AND2_X1   g233(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(G214), .B1(G237), .B2(G902), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n370), .A2(new_n193), .A3(new_n372), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT86), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(KEYINPUT87), .B(KEYINPUT5), .ZN(new_n426));
  INV_X1    g240(.A(G116), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n427), .A2(G119), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(G113), .B1(new_n426), .B2(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n430), .B1(new_n187), .B2(new_n426), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n431), .B1(new_n187), .B2(new_n191), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n369), .A2(new_n375), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n370), .A2(KEYINPUT86), .A3(new_n193), .A4(new_n372), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n425), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  XOR2_X1   g251(.A(G110), .B(G122), .Z(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n438), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n425), .A2(new_n440), .A3(new_n435), .A4(new_n436), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n439), .A2(KEYINPUT6), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n203), .A2(new_n302), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n443), .B1(new_n302), .B2(new_n227), .ZN(new_n444));
  XNOR2_X1  g258(.A(KEYINPUT88), .B(G224), .ZN(new_n445));
  INV_X1    g259(.A(G953), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n444), .B(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT6), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n437), .A2(new_n449), .A3(new_n438), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n442), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(KEYINPUT7), .B1(new_n445), .B2(new_n446), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n448), .B(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n432), .A2(new_n433), .ZN(new_n454));
  AND2_X1   g268(.A1(new_n187), .A2(KEYINPUT5), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n192), .B1(new_n430), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n434), .A2(new_n456), .ZN(new_n457));
  XOR2_X1   g271(.A(new_n438), .B(KEYINPUT8), .Z(new_n458));
  NAND3_X1  g272(.A1(new_n454), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n453), .A2(new_n441), .A3(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n451), .A2(new_n344), .A3(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(G210), .B1(G237), .B2(G902), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n451), .A2(new_n344), .A3(new_n462), .A4(new_n460), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n422), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n201), .A2(G128), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n318), .A2(G143), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n204), .ZN(new_n470));
  XNOR2_X1  g284(.A(G116), .B(G122), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n471), .B(new_n359), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT13), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n473), .B1(new_n318), .B2(G143), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(KEYINPUT93), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n201), .A2(KEYINPUT13), .A3(G128), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT93), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n467), .A2(new_n477), .A3(new_n473), .ZN(new_n478));
  AND4_X1   g292(.A1(new_n468), .A2(new_n475), .A3(new_n476), .A4(new_n478), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n470), .B(new_n472), .C1(new_n479), .C2(new_n204), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT94), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n480), .B(new_n481), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n469), .B(new_n204), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n427), .A2(KEYINPUT14), .A3(G122), .ZN(new_n484));
  INV_X1    g298(.A(new_n471), .ZN(new_n485));
  OAI211_X1 g299(.A(G107), .B(new_n484), .C1(new_n485), .C2(KEYINPUT14), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n483), .B(new_n486), .C1(G107), .C2(new_n485), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n482), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n417), .A2(G217), .A3(new_n446), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n489), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n482), .A2(new_n487), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n344), .ZN(new_n494));
  INV_X1    g308(.A(G478), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n495), .A2(KEYINPUT15), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n494), .B(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n311), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT90), .ZN(new_n500));
  INV_X1    g314(.A(G237), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n501), .A2(new_n446), .A3(G214), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n201), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n255), .A2(G143), .A3(G214), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n500), .B1(new_n505), .B2(G131), .ZN(new_n506));
  AOI211_X1 g320(.A(KEYINPUT90), .B(new_n213), .C1(new_n503), .C2(new_n504), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(KEYINPUT17), .ZN(new_n509));
  OAI22_X1  g323(.A1(new_n506), .A2(new_n507), .B1(G131), .B2(new_n505), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n499), .B(new_n509), .C1(KEYINPUT17), .C2(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(G113), .B(G122), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(new_n351), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT89), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT18), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n503), .B(new_n504), .C1(new_n515), .C2(new_n213), .ZN(new_n516));
  INV_X1    g330(.A(new_n300), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n517), .A2(G146), .A3(new_n298), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n324), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  AOI211_X1 g334(.A(new_n515), .B(new_n213), .C1(new_n503), .C2(new_n504), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n514), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n505), .A2(KEYINPUT18), .A3(G131), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n523), .A2(KEYINPUT89), .A3(new_n516), .A4(new_n519), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n511), .A2(new_n513), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n513), .B1(new_n511), .B2(new_n525), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n344), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(G475), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT20), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n517), .A2(new_n298), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n532), .B(KEYINPUT19), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n308), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n510), .A2(new_n323), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n513), .B1(new_n535), .B2(new_n525), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT91), .ZN(new_n537));
  OR2_X1    g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n536), .A2(new_n537), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n538), .A2(new_n526), .A3(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(G475), .ZN(new_n541));
  AND4_X1   g355(.A1(new_n531), .A2(new_n540), .A3(new_n541), .A4(new_n344), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n540), .A2(new_n541), .A3(new_n344), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(KEYINPUT20), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n542), .B1(KEYINPUT92), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT92), .ZN(new_n546));
  NOR3_X1   g360(.A1(new_n543), .A2(new_n546), .A3(KEYINPUT20), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n498), .B(new_n530), .C1(new_n545), .C2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(G952), .ZN(new_n550));
  AOI211_X1 g364(.A(G953), .B(new_n550), .C1(G234), .C2(G237), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  AOI211_X1 g366(.A(new_n344), .B(new_n446), .C1(G234), .C2(G237), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  XOR2_X1   g368(.A(KEYINPUT21), .B(G898), .Z(new_n555));
  OAI21_X1  g369(.A(new_n552), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n556), .B(KEYINPUT95), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n466), .A2(new_n549), .A3(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n350), .A2(new_n420), .A3(new_n560), .ZN(new_n561));
  XOR2_X1   g375(.A(new_n561), .B(new_n368), .Z(G3));
  NAND2_X1  g376(.A1(new_n416), .A2(new_n419), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n283), .A2(new_n344), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(G472), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n285), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT97), .ZN(new_n568));
  OR2_X1    g382(.A1(new_n492), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n492), .A2(new_n568), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n569), .A2(KEYINPUT33), .A3(new_n490), .A4(new_n570), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n495), .A2(G902), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT96), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT33), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n573), .B1(new_n493), .B2(new_n574), .ZN(new_n575));
  AOI211_X1 g389(.A(KEYINPUT96), .B(KEYINPUT33), .C1(new_n490), .C2(new_n492), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n571), .B(new_n572), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n494), .A2(new_n495), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n544), .A2(KEYINPUT92), .ZN(new_n581));
  INV_X1    g395(.A(new_n542), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n547), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n580), .B1(new_n585), .B2(new_n530), .ZN(new_n586));
  AND3_X1   g400(.A1(new_n466), .A2(new_n586), .A3(new_n558), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n567), .A2(new_n348), .A3(new_n587), .ZN(new_n588));
  XOR2_X1   g402(.A(KEYINPUT98), .B(KEYINPUT99), .Z(new_n589));
  XNOR2_X1  g403(.A(KEYINPUT34), .B(G104), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n589), .B(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n588), .B(new_n591), .ZN(G6));
  AOI22_X1  g406(.A1(new_n564), .A2(G472), .B1(new_n284), .B2(new_n283), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n593), .A2(new_n416), .A3(new_n348), .A4(new_n419), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n582), .A2(new_n544), .ZN(new_n595));
  AND3_X1   g409(.A1(new_n595), .A2(new_n497), .A3(new_n530), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n466), .A2(new_n558), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(KEYINPUT100), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT100), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n466), .A2(new_n599), .A3(new_n558), .A4(new_n596), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n594), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(KEYINPUT35), .B(G107), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(G9));
  NOR2_X1   g417(.A1(new_n334), .A2(KEYINPUT36), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n328), .B(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n605), .A2(new_n344), .A3(new_n345), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n342), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n567), .A2(new_n560), .A3(new_n607), .ZN(new_n608));
  XOR2_X1   g422(.A(KEYINPUT37), .B(G110), .Z(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(G12));
  INV_X1    g424(.A(new_n607), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n286), .A2(new_n288), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n296), .A2(G472), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  OR2_X1    g428(.A1(new_n554), .A2(G900), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n552), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n595), .A2(new_n497), .A3(new_n530), .A4(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(KEYINPUT101), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n614), .A2(new_n420), .A3(new_n466), .A4(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(G128), .ZN(G30));
  XNOR2_X1  g434(.A(new_n616), .B(KEYINPUT39), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n420), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT40), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n464), .A2(new_n465), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT38), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n464), .A2(KEYINPUT38), .A3(new_n465), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AOI22_X1  g443(.A1(new_n583), .A2(new_n584), .B1(G475), .B2(new_n529), .ZN(new_n630));
  NOR3_X1   g444(.A1(new_n629), .A2(new_n498), .A3(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n279), .A2(new_n266), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n344), .B1(new_n289), .B2(new_n259), .ZN(new_n633));
  OAI21_X1  g447(.A(G472), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n612), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NOR3_X1   g450(.A1(new_n636), .A2(new_n422), .A3(new_n607), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n624), .A2(new_n631), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(G143), .ZN(G45));
  OAI21_X1  g453(.A(new_n530), .B1(new_n545), .B2(new_n547), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n640), .A2(new_n579), .A3(new_n616), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n614), .A2(new_n420), .A3(new_n466), .A4(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G146), .ZN(G48));
  AND3_X1   g458(.A1(new_n283), .A2(new_n287), .A3(new_n284), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n287), .B1(new_n283), .B2(new_n284), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n613), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT102), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(G469), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n405), .A2(new_n344), .A3(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n649), .B1(new_n405), .B2(new_n344), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n651), .A2(new_n652), .A3(new_n418), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n587), .A2(new_n647), .A3(new_n348), .A4(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT41), .B(G113), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G15));
  NAND3_X1  g470(.A1(new_n653), .A2(new_n647), .A3(new_n348), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n657), .B1(new_n600), .B2(new_n598), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(new_n427), .ZN(G18));
  NAND3_X1  g473(.A1(new_n560), .A2(new_n614), .A3(new_n653), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G119), .ZN(G21));
  INV_X1    g475(.A(new_n284), .ZN(new_n662));
  OR2_X1    g476(.A1(new_n290), .A2(new_n259), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n662), .B1(new_n282), .B2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT103), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n565), .A2(KEYINPUT104), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT104), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n564), .A2(new_n668), .A3(G472), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n666), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  AND4_X1   g484(.A1(new_n497), .A2(new_n625), .A3(new_n640), .A4(new_n421), .ZN(new_n671));
  NOR4_X1   g485(.A1(new_n651), .A2(new_n652), .A3(new_n418), .A4(new_n557), .ZN(new_n672));
  XOR2_X1   g486(.A(new_n347), .B(KEYINPUT105), .Z(new_n673));
  NAND4_X1  g487(.A1(new_n670), .A2(new_n671), .A3(new_n672), .A4(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G122), .ZN(G24));
  INV_X1    g489(.A(new_n652), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n676), .A2(new_n419), .A3(new_n650), .ZN(new_n677));
  INV_X1    g491(.A(new_n466), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n679), .A2(new_n670), .A3(new_n607), .A4(new_n642), .ZN(new_n680));
  XNOR2_X1  g494(.A(KEYINPUT106), .B(G125), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G27));
  XOR2_X1   g496(.A(KEYINPUT107), .B(KEYINPUT42), .Z(new_n683));
  NAND3_X1  g497(.A1(new_n464), .A2(new_n421), .A3(new_n465), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n642), .A2(new_n685), .A3(new_n419), .A4(new_n416), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n647), .A2(new_n348), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n683), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n612), .A2(KEYINPUT108), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT108), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n286), .A2(new_n690), .A3(new_n288), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n689), .A2(new_n613), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n673), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n563), .A2(new_n641), .A3(new_n684), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(KEYINPUT42), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n688), .B1(new_n693), .B2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G131), .ZN(G33));
  NAND4_X1  g511(.A1(new_n350), .A2(new_n420), .A3(new_n618), .A4(new_n685), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G134), .ZN(G36));
  NAND3_X1  g513(.A1(new_n630), .A2(KEYINPUT43), .A3(new_n579), .ZN(new_n700));
  OAI211_X1 g514(.A(new_n579), .B(new_n530), .C1(new_n545), .C2(new_n547), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT43), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(KEYINPUT111), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n593), .A2(new_n611), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT44), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n705), .A2(KEYINPUT44), .A3(new_n706), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g525(.A(KEYINPUT45), .B1(new_n413), .B2(new_n414), .ZN(new_n712));
  OR3_X1    g526(.A1(new_n712), .A2(KEYINPUT109), .A3(new_n406), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n413), .A2(new_n414), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT45), .ZN(new_n715));
  OR3_X1    g529(.A1(new_n714), .A2(KEYINPUT110), .A3(new_n715), .ZN(new_n716));
  OAI21_X1  g530(.A(KEYINPUT110), .B1(new_n714), .B2(new_n715), .ZN(new_n717));
  OAI21_X1  g531(.A(KEYINPUT109), .B1(new_n712), .B2(new_n406), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n713), .A2(new_n716), .A3(new_n717), .A4(new_n718), .ZN(new_n719));
  AND3_X1   g533(.A1(new_n719), .A2(KEYINPUT46), .A3(new_n408), .ZN(new_n720));
  AOI21_X1  g534(.A(KEYINPUT46), .B1(new_n719), .B2(new_n408), .ZN(new_n721));
  INV_X1    g535(.A(new_n407), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n720), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n723), .A2(new_n418), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n684), .B(KEYINPUT112), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n724), .A2(new_n621), .A3(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n711), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(new_n211), .ZN(G39));
  INV_X1    g542(.A(KEYINPUT47), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n729), .B1(new_n723), .B2(new_n418), .ZN(new_n730));
  OR2_X1    g544(.A1(new_n721), .A2(new_n722), .ZN(new_n731));
  OAI211_X1 g545(.A(KEYINPUT47), .B(new_n419), .C1(new_n731), .C2(new_n720), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n647), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n641), .A2(new_n684), .A3(new_n348), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G140), .ZN(G42));
  NAND4_X1  g550(.A1(new_n647), .A2(new_n348), .A3(new_n419), .A4(new_n416), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n640), .A2(new_n580), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n466), .A2(new_n738), .A3(new_n548), .A4(new_n558), .ZN(new_n739));
  OAI22_X1  g553(.A1(new_n737), .A2(new_n559), .B1(new_n594), .B2(new_n739), .ZN(new_n740));
  NOR4_X1   g554(.A1(new_n559), .A2(new_n563), .A3(new_n566), .A4(new_n611), .ZN(new_n741));
  OAI21_X1  g555(.A(KEYINPUT114), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OR2_X1    g556(.A1(new_n594), .A2(new_n739), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT114), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n561), .A2(new_n608), .A3(new_n743), .A4(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n674), .A2(new_n654), .ZN(new_n747));
  NOR4_X1   g561(.A1(new_n559), .A2(new_n297), .A3(new_n677), .A4(new_n611), .ZN(new_n748));
  NOR3_X1   g562(.A1(new_n747), .A2(new_n658), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n664), .B(KEYINPUT103), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n668), .B1(new_n564), .B2(G472), .ZN(new_n752));
  INV_X1    g566(.A(G472), .ZN(new_n753));
  AOI211_X1 g567(.A(KEYINPUT104), .B(new_n753), .C1(new_n283), .C2(new_n344), .ZN(new_n754));
  OAI211_X1 g568(.A(new_n751), .B(new_n607), .C1(new_n752), .C2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n756), .A2(new_n694), .A3(KEYINPUT115), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT115), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n758), .B1(new_n686), .B2(new_n755), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n297), .A2(new_n563), .A3(new_n611), .ZN(new_n761));
  AND3_X1   g575(.A1(new_n685), .A2(new_n530), .A3(new_n595), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n761), .A2(new_n762), .A3(new_n498), .A4(new_n616), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n696), .A2(new_n760), .A3(new_n698), .A4(new_n763), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n750), .A2(new_n764), .ZN(new_n765));
  AND3_X1   g579(.A1(new_n680), .A2(new_n619), .A3(new_n643), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT117), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n607), .B1(new_n552), .B2(new_n615), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n671), .A2(new_n635), .A3(new_n420), .A4(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n766), .A2(new_n767), .A3(KEYINPUT52), .A4(new_n769), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n680), .A2(new_n619), .A3(new_n643), .A4(new_n769), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n761), .B(new_n466), .C1(new_n618), .C2(new_n642), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n774), .A2(KEYINPUT52), .A3(new_n680), .A4(new_n769), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n773), .A2(KEYINPUT117), .A3(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n765), .A2(KEYINPUT53), .A3(new_n770), .A4(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT54), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n598), .A2(new_n600), .ZN(new_n779));
  INV_X1    g593(.A(new_n657), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n781), .A2(new_n654), .A3(new_n660), .A4(new_n674), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n782), .B1(new_n745), .B2(new_n742), .ZN(new_n783));
  AND4_X1   g597(.A1(new_n696), .A2(new_n760), .A3(new_n698), .A4(new_n763), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n773), .A2(new_n775), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n783), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT53), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n777), .A2(new_n778), .A3(new_n788), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n786), .A2(new_n787), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n776), .A2(new_n770), .ZN(new_n791));
  OAI21_X1  g605(.A(KEYINPUT116), .B1(new_n750), .B2(new_n764), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT116), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n783), .A2(new_n784), .A3(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n791), .A2(new_n792), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n790), .B1(new_n795), .B2(new_n787), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n789), .B1(new_n796), .B2(new_n778), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n704), .A2(new_n551), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n799), .A2(new_n673), .A3(new_n670), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n653), .A2(new_n422), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT118), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(new_n629), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT119), .ZN(new_n805));
  OR3_X1    g619(.A1(new_n677), .A2(KEYINPUT118), .A3(new_n421), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n800), .A2(new_n804), .A3(new_n805), .A4(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT120), .ZN(new_n808));
  AOI21_X1  g622(.A(KEYINPUT50), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n636), .A2(new_n551), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n653), .A2(new_n685), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n812), .A2(new_n349), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n811), .A2(new_n630), .A3(new_n580), .A4(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n799), .A2(new_n806), .A3(new_n673), .A4(new_n670), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n815), .A2(new_n803), .ZN(new_n816));
  AOI21_X1  g630(.A(KEYINPUT119), .B1(new_n808), .B2(KEYINPUT50), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n814), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n809), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n651), .A2(new_n652), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(new_n418), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n730), .A2(new_n732), .A3(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n822), .A2(new_n725), .A3(new_n800), .ZN(new_n823));
  OR3_X1    g637(.A1(new_n798), .A2(new_n812), .A3(new_n755), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n819), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT51), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n811), .A2(new_n586), .A3(new_n813), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n819), .A2(new_n823), .A3(KEYINPUT51), .A4(new_n824), .ZN(new_n829));
  AOI211_X1 g643(.A(new_n550), .B(G953), .C1(new_n800), .C2(new_n679), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n693), .A2(new_n812), .A3(new_n798), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT48), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(KEYINPUT121), .ZN(new_n833));
  OR2_X1    g647(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  OR2_X1    g648(.A1(new_n832), .A2(KEYINPUT121), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n831), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n830), .A2(new_n834), .A3(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n827), .A2(new_n828), .A3(new_n829), .A4(new_n837), .ZN(new_n838));
  OAI22_X1  g652(.A1(new_n797), .A2(new_n838), .B1(G952), .B2(G953), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n820), .B(KEYINPUT49), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n840), .A2(new_n419), .A3(new_n421), .A4(new_n673), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n636), .A2(new_n629), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n841), .A2(new_n701), .A3(new_n842), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(KEYINPUT113), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n839), .A2(new_n844), .ZN(G75));
  NAND2_X1  g659(.A1(new_n777), .A2(new_n788), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n846), .A2(G210), .A3(G902), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT56), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n442), .A2(new_n450), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(new_n448), .ZN(new_n850));
  XOR2_X1   g664(.A(new_n850), .B(KEYINPUT55), .Z(new_n851));
  AOI21_X1  g665(.A(new_n851), .B1(KEYINPUT122), .B2(new_n848), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n847), .A2(new_n848), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n852), .B1(new_n847), .B2(new_n848), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n446), .A2(G952), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(G51));
  XOR2_X1   g670(.A(new_n408), .B(KEYINPUT57), .Z(new_n857));
  AND3_X1   g671(.A1(new_n777), .A2(new_n778), .A3(new_n788), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n778), .B1(new_n777), .B2(new_n788), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n857), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(new_n405), .ZN(new_n861));
  INV_X1    g675(.A(new_n846), .ZN(new_n862));
  OR3_X1    g676(.A1(new_n862), .A2(new_n344), .A3(new_n719), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n855), .B1(new_n861), .B2(new_n863), .ZN(G54));
  AOI21_X1  g678(.A(new_n344), .B1(new_n777), .B2(new_n788), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n865), .A2(KEYINPUT58), .A3(G475), .ZN(new_n866));
  INV_X1    g680(.A(new_n540), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n855), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n865), .A2(KEYINPUT58), .A3(G475), .A4(new_n540), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(G60));
  OR2_X1    g685(.A1(new_n575), .A2(new_n576), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n872), .A2(new_n571), .ZN(new_n873));
  NAND2_X1  g687(.A1(G478), .A2(G902), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(KEYINPUT59), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n873), .B1(new_n797), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n873), .A2(new_n875), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n878), .B1(new_n858), .B2(new_n859), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(new_n869), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n876), .A2(new_n880), .ZN(G63));
  NAND2_X1  g695(.A1(G217), .A2(G902), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(KEYINPUT60), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n846), .A2(new_n605), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n883), .B1(new_n777), .B2(new_n788), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n885), .B(new_n869), .C1(new_n343), .C2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT61), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  OR2_X1    g703(.A1(new_n886), .A2(new_n343), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n890), .A2(KEYINPUT61), .A3(new_n869), .A4(new_n885), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n889), .A2(new_n891), .ZN(G66));
  AOI21_X1  g706(.A(new_n446), .B1(new_n555), .B2(new_n445), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n893), .B1(new_n750), .B2(new_n446), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n849), .B1(G898), .B2(new_n446), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n894), .B(new_n895), .Z(G69));
  NAND3_X1  g710(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n272), .B(new_n533), .Z(new_n898));
  INV_X1    g712(.A(KEYINPUT62), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n638), .B(new_n766), .C1(KEYINPUT123), .C2(new_n899), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n899), .A2(KEYINPUT123), .ZN(new_n901));
  OR2_X1    g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n900), .A2(new_n901), .ZN(new_n903));
  AOI22_X1  g717(.A1(new_n902), .A2(new_n903), .B1(new_n733), .B2(new_n734), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n446), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n622), .A2(new_n684), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n906), .A2(new_n350), .A3(new_n548), .A4(new_n738), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT124), .ZN(new_n908));
  OAI21_X1  g722(.A(KEYINPUT125), .B1(new_n727), .B2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT124), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n907), .B(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT125), .ZN(new_n912));
  OAI211_X1 g726(.A(new_n911), .B(new_n912), .C1(new_n711), .C2(new_n726), .ZN(new_n913));
  AND2_X1   g727(.A1(new_n909), .A2(new_n913), .ZN(new_n914));
  OAI211_X1 g728(.A(new_n897), .B(new_n898), .C1(new_n905), .C2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n735), .A2(new_n766), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n696), .A2(new_n698), .ZN(new_n917));
  INV_X1    g731(.A(new_n693), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n724), .A2(new_n918), .A3(new_n621), .A4(new_n671), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n917), .B(new_n919), .C1(new_n711), .C2(new_n726), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n446), .B1(new_n916), .B2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(new_n898), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n384), .A2(G900), .A3(G953), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n915), .A2(new_n924), .ZN(G72));
  AND2_X1   g739(.A1(new_n279), .A2(new_n266), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n916), .A2(new_n920), .A3(new_n750), .ZN(new_n927));
  XOR2_X1   g741(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n928));
  NOR2_X1   g742(.A1(new_n753), .A2(new_n344), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n928), .B(new_n929), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n926), .B1(new_n927), .B2(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n750), .B1(new_n909), .B2(new_n913), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n930), .B1(new_n932), .B2(new_n904), .ZN(new_n933));
  INV_X1    g747(.A(new_n632), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n869), .B(new_n931), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n926), .A2(new_n632), .A3(new_n930), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT127), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n796), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n935), .A2(new_n938), .ZN(G57));
endmodule


