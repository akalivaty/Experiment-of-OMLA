//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 1 0 0 1 1 1 1 0 1 0 1 1 0 0 0 0 0 1 1 1 1 0 1 0 0 1 1 0 1 0 0 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 1 0 0 1 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:33 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n554, new_n556, new_n557, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n626, new_n627, new_n628, new_n631, new_n633,
    new_n634, new_n635, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1180, new_n1181, new_n1182, new_n1183, new_n1185;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT65), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT66), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  AND3_X1   g038(.A1(new_n461), .A2(new_n463), .A3(KEYINPUT67), .ZN(new_n464));
  AOI21_X1  g039(.A(KEYINPUT67), .B1(new_n461), .B2(new_n463), .ZN(new_n465));
  OAI21_X1  g040(.A(G125), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n459), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n461), .A2(new_n463), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G137), .ZN(new_n471));
  NAND2_X1  g046(.A1(G101), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(G2105), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n468), .A2(new_n473), .ZN(G160));
  NOR2_X1   g049(.A1(new_n469), .A2(new_n459), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n469), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  NOR2_X1   g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI21_X1  g054(.A(G2104), .B1(new_n459), .B2(G112), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n476), .B(new_n478), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G162));
  INV_X1    g057(.A(KEYINPUT68), .ZN(new_n483));
  NAND4_X1  g058(.A1(new_n461), .A2(new_n463), .A3(KEYINPUT4), .A4(G138), .ZN(new_n484));
  NAND2_X1  g059(.A1(G102), .A2(G2104), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(new_n459), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n461), .A2(new_n463), .A3(G126), .ZN(new_n488));
  NAND2_X1  g063(.A1(G114), .A2(G2104), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT67), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n462), .A2(G2104), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n461), .A2(new_n463), .A3(KEYINPUT67), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n459), .A2(G138), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g075(.A(KEYINPUT4), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n483), .B1(new_n492), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n500), .B1(new_n464), .B2(new_n465), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT4), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g080(.A(G2105), .B1(new_n484), .B2(new_n485), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n459), .B1(new_n488), .B2(new_n489), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n505), .A2(new_n508), .A3(KEYINPUT68), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n502), .A2(new_n509), .ZN(G164));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  OR2_X1    g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G50), .ZN(new_n515));
  XOR2_X1   g090(.A(new_n515), .B(KEYINPUT69), .Z(new_n516));
  NAND2_X1  g091(.A1(new_n511), .A2(KEYINPUT5), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G543), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n520), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n521));
  INV_X1    g096(.A(G651), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n516), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n512), .A2(new_n513), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n520), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(new_n527));
  XNOR2_X1  g102(.A(KEYINPUT70), .B(G88), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n524), .A2(new_n529), .ZN(G303));
  INV_X1    g105(.A(G303), .ZN(G166));
  NAND2_X1  g106(.A1(new_n525), .A2(G89), .ZN(new_n532));
  INV_X1    g107(.A(G63), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n533), .B2(new_n522), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n534), .A2(new_n520), .B1(G51), .B2(new_n514), .ZN(new_n535));
  XOR2_X1   g110(.A(KEYINPUT71), .B(KEYINPUT7), .Z(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n536), .B(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n535), .A2(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  AOI22_X1  g115(.A1(new_n520), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(new_n522), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n514), .A2(G52), .ZN(new_n543));
  XNOR2_X1  g118(.A(KEYINPUT72), .B(G90), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n526), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n542), .A2(new_n545), .ZN(G171));
  INV_X1    g121(.A(new_n514), .ZN(new_n547));
  XOR2_X1   g122(.A(KEYINPUT73), .B(G43), .Z(new_n548));
  NOR2_X1   g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n520), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n550), .A2(new_n522), .ZN(new_n551));
  AOI211_X1 g126(.A(new_n549), .B(new_n551), .C1(G81), .C2(new_n527), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  AND3_X1   g128(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G36), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n554), .A2(new_n557), .ZN(G188));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT76), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n517), .A2(new_n519), .A3(G65), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(KEYINPUT77), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT77), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n560), .A2(new_n564), .A3(new_n561), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n563), .A2(G651), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(KEYINPUT78), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT78), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n563), .A2(new_n568), .A3(new_n565), .A4(G651), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n527), .A2(G91), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT75), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT74), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT9), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n525), .A2(G53), .A3(G543), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n573), .A2(new_n574), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n575), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n579), .B1(new_n514), .B2(G53), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n572), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n576), .A2(new_n575), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n514), .A2(G53), .B1(new_n573), .B2(new_n574), .ZN(new_n583));
  OAI211_X1 g158(.A(new_n582), .B(KEYINPUT75), .C1(new_n583), .C2(new_n575), .ZN(new_n584));
  AND2_X1   g159(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n570), .A2(new_n571), .A3(new_n585), .ZN(G299));
  INV_X1    g161(.A(G171), .ZN(G301));
  NAND2_X1  g162(.A1(new_n514), .A2(G49), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT79), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n588), .B(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n527), .A2(G87), .ZN(new_n591));
  OAI21_X1  g166(.A(G651), .B1(new_n520), .B2(G74), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(G288));
  AOI22_X1  g168(.A1(new_n520), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n594), .A2(new_n522), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n514), .A2(G48), .ZN(new_n596));
  INV_X1    g171(.A(G86), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n526), .B2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n595), .A2(new_n599), .ZN(G305));
  AOI22_X1  g175(.A1(new_n520), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n601), .A2(new_n522), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n514), .A2(G47), .ZN(new_n603));
  INV_X1    g178(.A(G85), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n526), .B2(new_n604), .ZN(new_n605));
  OR3_X1    g180(.A1(new_n602), .A2(new_n605), .A3(KEYINPUT80), .ZN(new_n606));
  OAI21_X1  g181(.A(KEYINPUT80), .B1(new_n602), .B2(new_n605), .ZN(new_n607));
  AND2_X1   g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(G290));
  NAND2_X1  g184(.A1(G301), .A2(G868), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n527), .A2(G92), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT10), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n514), .A2(G54), .ZN(new_n613));
  XNOR2_X1  g188(.A(KEYINPUT81), .B(G66), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n520), .A2(new_n614), .B1(G79), .B2(G543), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n613), .B1(new_n615), .B2(new_n522), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(KEYINPUT82), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT82), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(new_n612), .B2(new_n616), .ZN(new_n620));
  AND3_X1   g195(.A1(new_n618), .A2(KEYINPUT83), .A3(new_n620), .ZN(new_n621));
  AOI21_X1  g196(.A(KEYINPUT83), .B1(new_n618), .B2(new_n620), .ZN(new_n622));
  NOR2_X1   g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n610), .B1(new_n623), .B2(G868), .ZN(G284));
  OAI21_X1  g199(.A(new_n610), .B1(new_n623), .B2(G868), .ZN(G321));
  NAND2_X1  g200(.A1(G286), .A2(G868), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT84), .Z(new_n627));
  XNOR2_X1  g202(.A(G299), .B(KEYINPUT85), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(new_n628), .B2(G868), .ZN(G297));
  OAI21_X1  g204(.A(new_n627), .B1(new_n628), .B2(G868), .ZN(G280));
  INV_X1    g205(.A(G559), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n623), .B1(new_n631), .B2(G860), .ZN(G148));
  NOR3_X1   g207(.A1(new_n621), .A2(new_n622), .A3(G559), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(G868), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n635), .B1(G868), .B2(new_n552), .ZN(G323));
  XNOR2_X1  g211(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g212(.A1(new_n498), .A2(G2104), .A3(new_n459), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT12), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT13), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2100), .ZN(new_n641));
  INV_X1    g216(.A(new_n477), .ZN(new_n642));
  INV_X1    g217(.A(G135), .ZN(new_n643));
  OR3_X1    g218(.A1(new_n642), .A2(KEYINPUT86), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n475), .A2(G123), .ZN(new_n645));
  OR2_X1    g220(.A1(G99), .A2(G2105), .ZN(new_n646));
  OAI211_X1 g221(.A(new_n646), .B(G2104), .C1(G111), .C2(new_n459), .ZN(new_n647));
  OAI21_X1  g222(.A(KEYINPUT86), .B1(new_n642), .B2(new_n643), .ZN(new_n648));
  NAND4_X1  g223(.A1(new_n644), .A2(new_n645), .A3(new_n647), .A4(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(G2096), .Z(new_n650));
  NAND2_X1  g225(.A1(new_n641), .A2(new_n650), .ZN(G156));
  XNOR2_X1  g226(.A(KEYINPUT15), .B(G2430), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2435), .ZN(new_n653));
  XOR2_X1   g228(.A(G2427), .B(G2438), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n655), .A2(KEYINPUT14), .ZN(new_n656));
  XOR2_X1   g231(.A(G2451), .B(G2454), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT16), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n656), .B(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G1341), .B(G1348), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2443), .B(G2446), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n661), .B(new_n662), .Z(new_n663));
  NAND2_X1  g238(.A1(new_n663), .A2(G14), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(G401));
  XNOR2_X1  g240(.A(G2084), .B(G2090), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT87), .ZN(new_n667));
  XOR2_X1   g242(.A(G2067), .B(G2678), .Z(new_n668));
  NOR2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2072), .B(G2078), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT17), .Z(new_n671));
  AOI21_X1  g246(.A(new_n671), .B1(new_n667), .B2(new_n668), .ZN(new_n672));
  INV_X1    g247(.A(new_n668), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n673), .A2(new_n670), .ZN(new_n674));
  AOI211_X1 g249(.A(new_n669), .B(new_n672), .C1(new_n667), .C2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n669), .A2(new_n670), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT18), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(G2096), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(G2100), .Z(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(G227));
  XOR2_X1   g256(.A(G1956), .B(G2474), .Z(new_n682));
  XOR2_X1   g257(.A(G1961), .B(G1966), .Z(new_n683));
  NOR2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1971), .B(G1976), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT19), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n682), .A2(new_n683), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT20), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n688), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n685), .A2(new_n687), .A3(new_n689), .ZN(new_n693));
  OAI211_X1 g268(.A(new_n692), .B(new_n693), .C1(new_n691), .C2(new_n690), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT21), .B(G1986), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(G1991), .B(G1996), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT22), .B(G1981), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n698), .B(new_n699), .Z(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(G229));
  NAND2_X1  g276(.A1(new_n608), .A2(G16), .ZN(new_n702));
  OR2_X1    g277(.A1(G16), .A2(G24), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(KEYINPUT89), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT89), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n702), .A2(new_n706), .A3(new_n703), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(G1986), .ZN(new_n709));
  INV_X1    g284(.A(G16), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n710), .A2(G22), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(G303), .B2(G16), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(G1971), .ZN(new_n713));
  MUX2_X1   g288(.A(G23), .B(G288), .S(G16), .Z(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT33), .B(G1976), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT90), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n714), .B(new_n716), .ZN(new_n717));
  MUX2_X1   g292(.A(G6), .B(G305), .S(G16), .Z(new_n718));
  XOR2_X1   g293(.A(KEYINPUT32), .B(G1981), .Z(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n713), .A2(new_n717), .A3(new_n720), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n721), .A2(KEYINPUT34), .ZN(new_n722));
  AND3_X1   g297(.A1(new_n721), .A2(KEYINPUT91), .A3(KEYINPUT34), .ZN(new_n723));
  AOI21_X1  g298(.A(KEYINPUT91), .B1(new_n721), .B2(KEYINPUT34), .ZN(new_n724));
  OAI211_X1 g299(.A(new_n709), .B(new_n722), .C1(new_n723), .C2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(G29), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G25), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n475), .A2(G119), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT88), .Z(new_n729));
  NAND2_X1  g304(.A1(new_n477), .A2(G131), .ZN(new_n730));
  NOR2_X1   g305(.A1(G95), .A2(G2105), .ZN(new_n731));
  OAI21_X1  g306(.A(G2104), .B1(new_n459), .B2(G107), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n729), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n727), .B1(new_n734), .B2(new_n726), .ZN(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT35), .B(G1991), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(KEYINPUT36), .B1(new_n725), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n721), .A2(KEYINPUT34), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n721), .A2(KEYINPUT34), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT91), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n721), .A2(KEYINPUT91), .A3(KEYINPUT34), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n739), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT36), .ZN(new_n745));
  INV_X1    g320(.A(new_n737), .ZN(new_n746));
  NAND4_X1  g321(.A1(new_n744), .A2(new_n745), .A3(new_n709), .A4(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n738), .A2(new_n747), .ZN(new_n748));
  AOI22_X1  g323(.A1(G129), .A2(new_n475), .B1(new_n477), .B2(G141), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n459), .A2(G105), .A3(G2104), .ZN(new_n750));
  XOR2_X1   g325(.A(KEYINPUT98), .B(KEYINPUT26), .Z(new_n751));
  NAND3_X1  g326(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  AND3_X1   g328(.A1(new_n749), .A2(new_n750), .A3(new_n753), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT99), .Z(new_n755));
  INV_X1    g330(.A(KEYINPUT100), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n754), .B(KEYINPUT99), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n758), .A2(KEYINPUT100), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n757), .A2(G29), .A3(new_n759), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT27), .B(G1996), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n726), .A2(G32), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n760), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n726), .A2(G35), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G162), .B2(new_n726), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT29), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n763), .B1(G2090), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n761), .B1(new_n760), .B2(new_n762), .ZN(new_n768));
  OR2_X1    g343(.A1(G29), .A2(G33), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n477), .A2(G139), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT25), .Z(new_n772));
  AOI22_X1  g347(.A1(new_n498), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n773));
  OAI211_X1 g348(.A(new_n770), .B(new_n772), .C1(new_n773), .C2(new_n459), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n769), .B1(new_n774), .B2(new_n726), .ZN(new_n775));
  INV_X1    g350(.A(G2072), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT95), .Z(new_n778));
  NOR3_X1   g353(.A1(new_n767), .A2(new_n768), .A3(new_n778), .ZN(new_n779));
  XOR2_X1   g354(.A(KEYINPUT31), .B(G11), .Z(new_n780));
  NAND2_X1  g355(.A1(G168), .A2(G16), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT101), .ZN(new_n782));
  OAI211_X1 g357(.A(new_n781), .B(new_n782), .C1(G16), .C2(G21), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(new_n782), .B2(new_n781), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n780), .B1(new_n784), .B2(G1966), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n784), .A2(G1966), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n786), .A2(KEYINPUT102), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT102), .ZN(new_n788));
  NOR3_X1   g363(.A1(new_n784), .A2(new_n788), .A3(G1966), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n775), .A2(new_n776), .ZN(new_n790));
  NOR3_X1   g365(.A1(new_n787), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n766), .A2(G2090), .ZN(new_n792));
  NOR2_X1   g367(.A1(G5), .A2(G16), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G171), .B2(G16), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G1961), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n649), .A2(new_n726), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT30), .ZN(new_n797));
  AND2_X1   g372(.A1(new_n797), .A2(G28), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n797), .A2(G28), .ZN(new_n799));
  NOR3_X1   g374(.A1(new_n798), .A2(new_n799), .A3(G29), .ZN(new_n800));
  NOR4_X1   g375(.A1(new_n792), .A2(new_n795), .A3(new_n796), .A4(new_n800), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n779), .A2(new_n785), .A3(new_n791), .A4(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(G16), .B1(new_n621), .B2(new_n622), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n710), .A2(G4), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(G1348), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n803), .A2(G1348), .A3(new_n804), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n726), .A2(G26), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n475), .A2(G128), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n811), .A2(KEYINPUT93), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n477), .A2(G140), .ZN(new_n813));
  OR2_X1    g388(.A1(G104), .A2(G2105), .ZN(new_n814));
  OAI211_X1 g389(.A(new_n814), .B(G2104), .C1(G116), .C2(new_n459), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n811), .A2(KEYINPUT93), .ZN(new_n816));
  NAND4_X1  g391(.A1(new_n812), .A2(new_n813), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n810), .B1(new_n818), .B2(new_n726), .ZN(new_n819));
  MUX2_X1   g394(.A(new_n810), .B(new_n819), .S(KEYINPUT28), .Z(new_n820));
  INV_X1    g395(.A(G2067), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n710), .A2(G19), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(new_n552), .B2(new_n710), .ZN(new_n824));
  XOR2_X1   g399(.A(KEYINPUT92), .B(G1341), .Z(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n809), .A2(new_n822), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(KEYINPUT94), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT94), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n809), .A2(new_n829), .A3(new_n822), .A4(new_n826), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n802), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(G27), .ZN(new_n832));
  OAI21_X1  g407(.A(KEYINPUT103), .B1(new_n832), .B2(G29), .ZN(new_n833));
  OR3_X1    g408(.A1(new_n832), .A2(KEYINPUT103), .A3(G29), .ZN(new_n834));
  OAI211_X1 g409(.A(new_n833), .B(new_n834), .C1(G164), .C2(new_n726), .ZN(new_n835));
  INV_X1    g410(.A(G2078), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT24), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n726), .B1(new_n838), .B2(G34), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n839), .A2(KEYINPUT96), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n838), .A2(G34), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n839), .A2(KEYINPUT96), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n843), .A2(KEYINPUT97), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n844), .B1(G160), .B2(G29), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n843), .A2(KEYINPUT97), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(G2084), .ZN(new_n848));
  NAND4_X1  g423(.A1(new_n748), .A2(new_n831), .A3(new_n837), .A4(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n710), .A2(G20), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(KEYINPUT104), .Z(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT23), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n852), .B1(G299), .B2(G16), .ZN(new_n853));
  INV_X1    g428(.A(G1956), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n849), .A2(new_n855), .ZN(G311));
  AND3_X1   g431(.A1(new_n748), .A2(new_n848), .A3(new_n831), .ZN(new_n857));
  INV_X1    g432(.A(new_n855), .ZN(new_n858));
  NAND4_X1  g433(.A1(new_n857), .A2(KEYINPUT105), .A3(new_n858), .A4(new_n837), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT105), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n860), .B1(new_n849), .B2(new_n855), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(new_n861), .ZN(G150));
  NAND2_X1  g437(.A1(new_n514), .A2(G55), .ZN(new_n863));
  INV_X1    g438(.A(G93), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n863), .B1(new_n526), .B2(new_n864), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n865), .B(KEYINPUT108), .Z(new_n866));
  AOI22_X1  g441(.A1(new_n520), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT107), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n868), .A2(new_n522), .ZN(new_n869));
  OAI21_X1  g444(.A(G860), .B1(new_n866), .B2(new_n869), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n870), .B(KEYINPUT37), .Z(new_n871));
  NAND2_X1  g446(.A1(new_n623), .A2(G559), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT109), .ZN(new_n873));
  XOR2_X1   g448(.A(KEYINPUT106), .B(KEYINPUT38), .Z(new_n874));
  XNOR2_X1  g449(.A(new_n873), .B(new_n874), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n866), .A2(new_n869), .ZN(new_n876));
  XOR2_X1   g451(.A(new_n876), .B(new_n552), .Z(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT39), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n875), .B(new_n878), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n871), .B1(new_n879), .B2(G860), .ZN(G145));
  NAND2_X1  g455(.A1(new_n475), .A2(G130), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n477), .A2(G142), .ZN(new_n882));
  NOR2_X1   g457(.A1(G106), .A2(G2105), .ZN(new_n883));
  OAI21_X1  g458(.A(G2104), .B1(new_n459), .B2(G118), .ZN(new_n884));
  OAI211_X1 g459(.A(new_n881), .B(new_n882), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n639), .B(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n734), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n886), .B(new_n887), .ZN(new_n888));
  AND2_X1   g463(.A1(new_n757), .A2(new_n759), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n499), .B1(new_n496), .B2(new_n497), .ZN(new_n890));
  OAI211_X1 g465(.A(new_n487), .B(new_n491), .C1(new_n890), .C2(KEYINPUT4), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n817), .B(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n889), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n757), .A2(new_n759), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(new_n892), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n774), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n755), .A2(new_n892), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(new_n774), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n755), .A2(new_n892), .ZN(new_n900));
  OAI21_X1  g475(.A(KEYINPUT110), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n897), .A2(new_n901), .ZN(new_n902));
  AOI211_X1 g477(.A(KEYINPUT110), .B(new_n774), .C1(new_n894), .C2(new_n896), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n888), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT110), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n897), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n888), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n906), .B(new_n907), .C1(new_n897), .C2(new_n901), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n649), .B(G160), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(G162), .ZN(new_n910));
  AND3_X1   g485(.A1(new_n904), .A2(new_n908), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n910), .B1(new_n904), .B2(new_n908), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(G37), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n915), .B(KEYINPUT40), .ZN(G395));
  OR2_X1    g491(.A1(new_n633), .A2(new_n877), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n633), .A2(new_n877), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(G299), .B(new_n617), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  XOR2_X1   g497(.A(new_n920), .B(KEYINPUT41), .Z(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n924), .A2(new_n917), .A3(new_n918), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n922), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(KEYINPUT42), .ZN(new_n927));
  XOR2_X1   g502(.A(new_n608), .B(G305), .Z(new_n928));
  XNOR2_X1  g503(.A(G303), .B(G288), .ZN(new_n929));
  XOR2_X1   g504(.A(new_n928), .B(new_n929), .Z(new_n930));
  INV_X1    g505(.A(KEYINPUT42), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n922), .A2(new_n931), .A3(new_n925), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n927), .A2(new_n930), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n930), .B1(new_n927), .B2(new_n932), .ZN(new_n934));
  OAI21_X1  g509(.A(G868), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n935), .B1(G868), .B2(new_n876), .ZN(G295));
  OAI21_X1  g511(.A(new_n935), .B1(G868), .B2(new_n876), .ZN(G331));
  XNOR2_X1  g512(.A(G286), .B(G171), .ZN(new_n938));
  OR2_X1    g513(.A1(new_n877), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n877), .A2(new_n938), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(new_n923), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n939), .A2(new_n920), .A3(new_n940), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(KEYINPUT112), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT112), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n942), .A2(new_n943), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n945), .A2(new_n930), .A3(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n914), .B1(new_n944), .B2(new_n930), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT43), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n948), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n944), .A2(new_n930), .ZN(new_n953));
  OAI21_X1  g528(.A(KEYINPUT43), .B1(new_n953), .B2(new_n949), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n952), .A2(KEYINPUT44), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n951), .B1(new_n948), .B2(new_n950), .ZN(new_n956));
  NOR3_X1   g531(.A1(new_n953), .A2(new_n949), .A3(KEYINPUT43), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  XOR2_X1   g533(.A(KEYINPUT111), .B(KEYINPUT44), .Z(new_n959));
  OAI21_X1  g534(.A(new_n955), .B1(new_n958), .B2(new_n959), .ZN(G397));
  INV_X1    g535(.A(G40), .ZN(new_n961));
  NOR3_X1   g536(.A1(new_n468), .A2(new_n961), .A3(new_n473), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT45), .ZN(new_n963));
  INV_X1    g538(.A(G1384), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n964), .B1(new_n492), .B2(new_n501), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n962), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n889), .A2(G1996), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n817), .B(G2067), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n967), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n758), .A2(new_n967), .A3(G1996), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(KEYINPUT113), .ZN(new_n972));
  OR2_X1    g547(.A1(new_n971), .A2(KEYINPUT113), .ZN(new_n973));
  AND3_X1   g548(.A1(new_n970), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n734), .B(new_n736), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n974), .B1(new_n966), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(G1986), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n608), .B(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n976), .B1(new_n978), .B2(new_n967), .ZN(new_n979));
  XNOR2_X1  g554(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n980), .B1(G303), .B2(G8), .ZN(new_n981));
  INV_X1    g556(.A(G8), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n982), .B1(new_n524), .B2(new_n529), .ZN(new_n983));
  NOR2_X1   g558(.A1(KEYINPUT115), .A2(KEYINPUT55), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n981), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT50), .ZN(new_n986));
  AOI211_X1 g561(.A(KEYINPUT114), .B(G1384), .C1(new_n505), .C2(new_n508), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT114), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n988), .B1(new_n891), .B2(new_n964), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n986), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n502), .A2(new_n964), .A3(new_n509), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(KEYINPUT50), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n990), .A2(new_n992), .A3(new_n962), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n993), .A2(G2090), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n891), .A2(KEYINPUT45), .A3(new_n964), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n962), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n996), .B1(new_n963), .B2(new_n991), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n997), .A2(G1971), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n985), .B(G8), .C1(new_n994), .C2(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n962), .B1(new_n987), .B2(new_n989), .ZN(new_n1000));
  INV_X1    g575(.A(G1976), .ZN(new_n1001));
  OR2_X1    g576(.A1(G288), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1000), .A2(G8), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT52), .ZN(new_n1004));
  NAND2_X1  g579(.A1(G305), .A2(G1981), .ZN(new_n1005));
  INV_X1    g580(.A(G1981), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n595), .A2(new_n599), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT49), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1005), .A2(KEYINPUT49), .A3(new_n1007), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1010), .A2(G8), .A3(new_n1000), .A4(new_n1011), .ZN(new_n1012));
  XOR2_X1   g587(.A(KEYINPUT116), .B(G1976), .Z(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT52), .B1(G288), .B2(new_n1013), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1000), .A2(G8), .A3(new_n1002), .A4(new_n1014), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n1004), .A2(new_n1012), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n998), .ZN(new_n1017));
  NOR3_X1   g592(.A1(new_n987), .A2(new_n989), .A3(new_n986), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n502), .A2(new_n986), .A3(new_n964), .A4(new_n509), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(new_n962), .ZN(new_n1020));
  OR3_X1    g595(.A1(new_n1018), .A2(new_n1020), .A3(G2090), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n982), .B1(new_n1017), .B2(new_n1021), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n999), .B(new_n1016), .C1(new_n1022), .C2(new_n985), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n821), .B(new_n962), .C1(new_n987), .C2(new_n989), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1025), .B1(new_n993), .B2(new_n806), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT125), .ZN(new_n1027));
  AND3_X1   g602(.A1(new_n1026), .A2(new_n1027), .A3(KEYINPUT60), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1027), .B1(new_n1026), .B2(KEYINPUT60), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n618), .A2(new_n620), .ZN(new_n1030));
  NOR3_X1   g605(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1026), .A2(KEYINPUT60), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1032), .A2(KEYINPUT125), .A3(new_n1030), .ZN(new_n1033));
  OR2_X1    g608(.A1(new_n1026), .A2(KEYINPUT60), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(KEYINPUT126), .B1(new_n1031), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT122), .ZN(new_n1037));
  INV_X1    g612(.A(new_n473), .ZN(new_n1038));
  AND2_X1   g613(.A1(new_n466), .A2(new_n467), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n1038), .B(G40), .C1(new_n1039), .C2(new_n459), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n965), .A2(KEYINPUT114), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n891), .A2(new_n988), .A3(new_n964), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1040), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g618(.A(KEYINPUT58), .B(G1341), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1037), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n996), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n991), .A2(new_n963), .ZN(new_n1047));
  INV_X1    g622(.A(G1996), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1044), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1000), .A2(KEYINPUT122), .A3(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1045), .A2(new_n1049), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(KEYINPUT123), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT123), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1045), .A2(new_n1054), .A3(new_n1049), .A4(new_n1051), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1053), .A2(new_n552), .A3(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT59), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1053), .A2(KEYINPUT59), .A3(new_n552), .A4(new_n1055), .ZN(new_n1059));
  AND2_X1   g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1041), .A2(KEYINPUT50), .A3(new_n1042), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1061), .A2(new_n962), .A3(new_n1019), .ZN(new_n1062));
  XNOR2_X1  g637(.A(KEYINPUT56), .B(G2072), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n1062), .A2(new_n854), .B1(new_n997), .B2(new_n1063), .ZN(new_n1064));
  AOI22_X1  g639(.A1(new_n567), .A2(new_n569), .B1(G91), .B2(new_n527), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n578), .A2(new_n580), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1066), .A2(KEYINPUT57), .ZN(new_n1067));
  AOI22_X1  g642(.A1(G299), .A2(KEYINPUT57), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1064), .A2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n854), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1046), .A2(new_n1047), .A3(new_n1063), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1068), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT61), .B1(new_n1069), .B2(new_n1074), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1070), .A2(KEYINPUT124), .A3(new_n1068), .A4(new_n1071), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(KEYINPUT61), .ZN(new_n1077));
  OAI21_X1  g652(.A(KEYINPUT121), .B1(new_n1064), .B2(new_n1068), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT121), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1072), .A2(new_n1079), .A3(new_n1073), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1077), .B1(new_n1078), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT124), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1069), .A2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1075), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1032), .A2(KEYINPUT125), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n618), .A2(new_n620), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1026), .A2(new_n1027), .A3(KEYINPUT60), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT126), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1088), .A2(new_n1089), .A3(new_n1034), .A4(new_n1033), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1036), .A2(new_n1060), .A3(new_n1084), .A4(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1026), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(new_n1086), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT120), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1093), .A2(KEYINPUT120), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1069), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1091), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT53), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1100), .B1(new_n1101), .B2(G2078), .ZN(new_n1102));
  INV_X1    g677(.A(G1961), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n993), .A2(new_n1103), .ZN(new_n1104));
  AND2_X1   g679(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1046), .A2(KEYINPUT53), .A3(new_n836), .A4(new_n966), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1105), .A2(KEYINPUT127), .A3(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1102), .A2(new_n1104), .A3(new_n1106), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT127), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(G301), .B1(new_n1107), .B2(new_n1110), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n1102), .A2(new_n1104), .A3(G301), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n962), .B1(new_n991), .B2(new_n963), .ZN(new_n1113));
  NOR3_X1   g688(.A1(new_n987), .A2(new_n989), .A3(KEYINPUT45), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1115), .A2(KEYINPUT53), .A3(new_n836), .ZN(new_n1116));
  AND2_X1   g691(.A1(new_n1112), .A2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(KEYINPUT54), .B1(new_n1111), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1105), .A2(new_n1116), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(G171), .ZN(new_n1120));
  AOI21_X1  g695(.A(KEYINPUT54), .B1(new_n1112), .B2(new_n1106), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(KEYINPUT117), .B1(new_n1115), .B2(G1966), .ZN(new_n1123));
  OR2_X1    g698(.A1(new_n993), .A2(G2084), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT117), .ZN(new_n1125));
  INV_X1    g700(.A(G1966), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1125), .B(new_n1126), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1123), .A2(new_n1124), .A3(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(G8), .B1(new_n1128), .B2(G286), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT51), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1130), .B1(new_n1128), .B2(G286), .ZN(new_n1131));
  OR2_X1    g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1129), .A2(KEYINPUT51), .ZN(new_n1133));
  AOI22_X1  g708(.A1(new_n1118), .A2(new_n1122), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1099), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(KEYINPUT62), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1120), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT62), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1132), .A2(new_n1139), .A3(new_n1133), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1137), .A2(new_n1138), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1023), .B1(new_n1135), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(new_n999), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1012), .A2(new_n1001), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1007), .B1(new_n1144), .B2(G288), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1043), .A2(new_n982), .ZN(new_n1146));
  AOI22_X1  g721(.A1(new_n1143), .A2(new_n1016), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1128), .A2(G8), .A3(G168), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(KEYINPUT118), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT118), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1128), .A2(new_n1150), .A3(G8), .A4(G168), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1023), .ZN(new_n1153));
  AOI21_X1  g728(.A(KEYINPUT119), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT119), .ZN(new_n1155));
  AOI211_X1 g730(.A(new_n1155), .B(new_n1023), .C1(new_n1149), .C2(new_n1151), .ZN(new_n1156));
  NOR3_X1   g731(.A1(new_n1154), .A2(new_n1156), .A3(KEYINPUT63), .ZN(new_n1157));
  INV_X1    g732(.A(new_n994), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n982), .B1(new_n1158), .B2(new_n1017), .ZN(new_n1159));
  OAI211_X1 g734(.A(new_n1152), .B(KEYINPUT63), .C1(new_n985), .C2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n999), .A2(new_n1016), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1147), .B1(new_n1157), .B2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n979), .B1(new_n1142), .B2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n967), .A2(new_n977), .A3(new_n608), .ZN(new_n1165));
  XOR2_X1   g740(.A(new_n1165), .B(KEYINPUT48), .Z(new_n1166));
  NOR2_X1   g741(.A1(new_n976), .A2(new_n1166), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n887), .A2(new_n736), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n974), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n818), .A2(new_n821), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n966), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  OR2_X1    g746(.A1(new_n969), .A2(new_n758), .ZN(new_n1172));
  OAI21_X1  g747(.A(KEYINPUT46), .B1(new_n966), .B2(G1996), .ZN(new_n1173));
  OR3_X1    g748(.A1(new_n966), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1174));
  AOI22_X1  g749(.A1(new_n1172), .A2(new_n967), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  XNOR2_X1  g750(.A(new_n1175), .B(KEYINPUT47), .ZN(new_n1176));
  NOR3_X1   g751(.A1(new_n1167), .A2(new_n1171), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1164), .A2(new_n1177), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g753(.A1(new_n664), .A2(new_n680), .ZN(new_n1180));
  AOI21_X1  g754(.A(new_n1180), .B1(new_n913), .B2(new_n914), .ZN(new_n1181));
  INV_X1    g755(.A(new_n1181), .ZN(new_n1182));
  OAI211_X1 g756(.A(new_n457), .B(new_n700), .C1(new_n956), .C2(new_n957), .ZN(new_n1183));
  NOR2_X1   g757(.A1(new_n1182), .A2(new_n1183), .ZN(G308));
  INV_X1    g758(.A(new_n958), .ZN(new_n1185));
  NAND4_X1  g759(.A1(new_n1185), .A2(new_n457), .A3(new_n700), .A4(new_n1181), .ZN(G225));
endmodule


