//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 1 0 0 1 0 0 1 0 1 0 1 1 0 1 1 1 0 1 0 1 0 0 0 0 0 0 1 1 0 1 1 0 1 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n779, new_n780, new_n781, new_n783, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n852, new_n853, new_n855, new_n856, new_n857,
    new_n858, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965;
  XOR2_X1   g000(.A(G190gat), .B(G218gat), .Z(new_n202));
  INV_X1    g001(.A(KEYINPUT102), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XOR2_X1   g003(.A(KEYINPUT96), .B(KEYINPUT17), .Z(new_n205));
  XOR2_X1   g004(.A(G43gat), .B(G50gat), .Z(new_n206));
  INV_X1    g005(.A(KEYINPUT15), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g007(.A1(G29gat), .A2(G36gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT14), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT14), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n211), .B1(G29gat), .B2(G36gat), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n210), .B1(new_n212), .B2(new_n209), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n208), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT94), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n214), .B(new_n215), .ZN(new_n216));
  AND2_X1   g015(.A1(new_n206), .A2(new_n207), .ZN(new_n217));
  OR3_X1    g016(.A1(new_n217), .A2(new_n208), .A3(new_n213), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n216), .A2(KEYINPUT95), .A3(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(KEYINPUT95), .B1(new_n216), .B2(new_n218), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n205), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n216), .A2(KEYINPUT17), .A3(new_n218), .ZN(new_n223));
  NAND2_X1  g022(.A1(G85gat), .A2(G92gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT7), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n225), .B(KEYINPUT99), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT100), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n227), .B1(new_n224), .B2(KEYINPUT7), .ZN(new_n228));
  OR3_X1    g027(.A1(new_n224), .A2(new_n227), .A3(KEYINPUT7), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n226), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(G99gat), .A2(G106gat), .ZN(new_n231));
  INV_X1    g030(.A(G85gat), .ZN(new_n232));
  INV_X1    g031(.A(G92gat), .ZN(new_n233));
  AOI22_X1  g032(.A1(KEYINPUT8), .A2(new_n231), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n230), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(G99gat), .B(G106gat), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT101), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n230), .A2(new_n236), .A3(new_n234), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n238), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n235), .A2(KEYINPUT101), .A3(new_n237), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n222), .A2(new_n223), .A3(new_n244), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n243), .B1(new_n220), .B2(new_n221), .ZN(new_n246));
  NAND3_X1  g045(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n245), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(G162gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n202), .A2(new_n203), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n248), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n249), .B1(new_n248), .B2(new_n250), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n204), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n253), .ZN(new_n255));
  INV_X1    g054(.A(new_n204), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n255), .A2(new_n256), .A3(new_n251), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n259), .B(G134gat), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n254), .A2(new_n257), .A3(new_n260), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT98), .ZN(new_n265));
  XNOR2_X1  g064(.A(G57gat), .B(G64gat), .ZN(new_n266));
  AND2_X1   g065(.A1(G71gat), .A2(G78gat), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n267), .A2(KEYINPUT9), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n265), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  NOR2_X1   g068(.A1(G71gat), .A2(G78gat), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  XOR2_X1   g070(.A(new_n269), .B(new_n271), .Z(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n273), .A2(KEYINPUT21), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n274), .B(G127gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(G15gat), .B(G22gat), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT16), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n276), .B1(new_n277), .B2(G1gat), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n278), .B1(G1gat), .B2(new_n276), .ZN(new_n279));
  INV_X1    g078(.A(G8gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n282), .B1(KEYINPUT21), .B2(new_n273), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n275), .B(new_n283), .ZN(new_n284));
  XOR2_X1   g083(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n285));
  XNOR2_X1  g084(.A(G155gat), .B(G183gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n284), .B(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(G231gat), .A2(G233gat), .ZN(new_n289));
  INV_X1    g088(.A(G211gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n289), .B(new_n290), .ZN(new_n291));
  XOR2_X1   g090(.A(new_n288), .B(new_n291), .Z(new_n292));
  XNOR2_X1  g091(.A(G120gat), .B(G148gat), .ZN(new_n293));
  INV_X1    g092(.A(G176gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n293), .B(new_n294), .ZN(new_n295));
  XOR2_X1   g094(.A(new_n295), .B(G204gat), .Z(new_n296));
  INV_X1    g095(.A(G230gat), .ZN(new_n297));
  INV_X1    g096(.A(G233gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n273), .A2(new_n238), .A3(new_n240), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT103), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n303), .B1(new_n243), .B2(new_n273), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n241), .A2(new_n272), .A3(KEYINPUT103), .A4(new_n242), .ZN(new_n305));
  AOI211_X1 g104(.A(KEYINPUT10), .B(new_n302), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n243), .A2(KEYINPUT10), .A3(new_n273), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n300), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n304), .A2(new_n305), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(new_n301), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(new_n299), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n309), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT104), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n296), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n296), .ZN(new_n316));
  AOI211_X1 g115(.A(KEYINPUT104), .B(new_n316), .C1(new_n309), .C2(new_n312), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n264), .A2(new_n292), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT97), .ZN(new_n320));
  OR2_X1    g119(.A1(G127gat), .A2(G134gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(G127gat), .A2(G134gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT71), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(G113gat), .ZN(new_n326));
  INV_X1    g125(.A(G120gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT1), .ZN(new_n329));
  NAND2_X1  g128(.A1(G113gat), .A2(G120gat), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n321), .A2(KEYINPUT71), .A3(new_n322), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n325), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  AND2_X1   g132(.A1(G113gat), .A2(G120gat), .ZN(new_n334));
  NOR2_X1   g133(.A1(G113gat), .A2(G120gat), .ZN(new_n335));
  OAI21_X1  g134(.A(KEYINPUT72), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT72), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n328), .A2(new_n337), .A3(new_n330), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n329), .A2(KEYINPUT73), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT73), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT1), .ZN(new_n342));
  AOI22_X1  g141(.A1(new_n340), .A2(new_n342), .B1(new_n321), .B2(new_n322), .ZN(new_n343));
  AND3_X1   g142(.A1(new_n339), .A2(KEYINPUT74), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT74), .B1(new_n339), .B2(new_n343), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n333), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(G155gat), .A2(G162gat), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NOR2_X1   g147(.A1(G155gat), .A2(G162gat), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(G141gat), .B(G148gat), .ZN(new_n351));
  AND2_X1   g150(.A1(new_n347), .A2(KEYINPUT2), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n350), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(G141gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(G148gat), .ZN(new_n355));
  INV_X1    g154(.A(G148gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(G141gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(G155gat), .B(G162gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n347), .A2(KEYINPUT2), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT3), .ZN(new_n362));
  AND3_X1   g161(.A1(new_n353), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n362), .B1(new_n353), .B2(new_n361), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n346), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT4), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT75), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n339), .A2(new_n343), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT74), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n339), .A2(KEYINPUT74), .A3(new_n343), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n368), .B1(new_n373), .B2(new_n333), .ZN(new_n374));
  OAI211_X1 g173(.A(new_n368), .B(new_n333), .C1(new_n344), .C2(new_n345), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n353), .A2(new_n361), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n367), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n378), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n380), .B(new_n333), .C1(new_n344), .C2(new_n345), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT4), .ZN(new_n383));
  AOI21_X1  g182(.A(KEYINPUT85), .B1(new_n379), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n346), .A2(KEYINPUT75), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n378), .B1(new_n385), .B2(new_n375), .ZN(new_n386));
  OAI211_X1 g185(.A(KEYINPUT85), .B(new_n383), .C1(new_n386), .C2(KEYINPUT4), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n366), .B1(new_n384), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(G225gat), .A2(G233gat), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  AND2_X1   g191(.A1(new_n325), .A2(new_n332), .ZN(new_n393));
  AOI22_X1  g192(.A1(new_n371), .A2(new_n372), .B1(new_n331), .B2(new_n393), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n394), .A2(new_n380), .ZN(new_n395));
  OR3_X1    g194(.A1(new_n395), .A2(new_n391), .A3(new_n382), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n392), .A2(KEYINPUT39), .A3(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(G1gat), .B(G29gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(new_n398), .B(KEYINPUT0), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n399), .B(G57gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n400), .B(new_n232), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT39), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n389), .A2(new_n402), .A3(new_n391), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n397), .A2(new_n401), .A3(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT40), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n391), .A2(KEYINPUT5), .ZN(new_n407));
  OAI211_X1 g206(.A(new_n366), .B(new_n407), .C1(new_n384), .C2(new_n388), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT84), .ZN(new_n409));
  AOI211_X1 g208(.A(new_n367), .B(new_n378), .C1(new_n385), .C2(new_n375), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n367), .B1(new_n346), .B2(new_n365), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n390), .B1(new_n411), .B2(new_n382), .ZN(new_n412));
  OAI21_X1  g211(.A(KEYINPUT83), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n364), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n353), .A2(new_n361), .A3(new_n362), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(KEYINPUT4), .B1(new_n394), .B2(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n391), .B1(new_n417), .B2(new_n381), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT83), .ZN(new_n419));
  OAI211_X1 g218(.A(KEYINPUT4), .B(new_n380), .C1(new_n374), .C2(new_n376), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n418), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n413), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n391), .B1(new_n395), .B2(new_n382), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT5), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n409), .B1(new_n422), .B2(new_n425), .ZN(new_n426));
  AOI211_X1 g225(.A(KEYINPUT84), .B(new_n424), .C1(new_n413), .C2(new_n421), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n408), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n401), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n397), .A2(KEYINPUT40), .A3(new_n401), .A4(new_n403), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT22), .ZN(new_n432));
  INV_X1    g231(.A(G218gat), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n432), .B1(new_n290), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT79), .ZN(new_n435));
  XNOR2_X1  g234(.A(G197gat), .B(G204gat), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT79), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n437), .B(new_n432), .C1(new_n290), .C2(new_n433), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n435), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  XNOR2_X1  g238(.A(G211gat), .B(G218gat), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n435), .A2(new_n440), .A3(new_n436), .A4(new_n438), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT80), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n442), .A2(KEYINPUT80), .A3(new_n443), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT29), .ZN(new_n450));
  NAND2_X1  g249(.A1(G226gat), .A2(G233gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(KEYINPUT27), .B(G183gat), .ZN(new_n452));
  INV_X1    g251(.A(G190gat), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n452), .A2(KEYINPUT28), .A3(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(G183gat), .ZN(new_n456));
  OAI21_X1  g255(.A(KEYINPUT27), .B1(new_n456), .B2(KEYINPUT67), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT67), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT27), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n458), .A2(new_n459), .A3(G183gat), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n457), .A2(new_n460), .A3(new_n453), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT68), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT28), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n457), .A2(new_n460), .A3(KEYINPUT68), .A4(new_n453), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT69), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n463), .A2(KEYINPUT69), .A3(new_n464), .A4(new_n465), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n455), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(G169gat), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n471), .A2(new_n294), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n294), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n473), .A2(KEYINPUT26), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(KEYINPUT26), .ZN(new_n475));
  OR2_X1    g274(.A1(new_n475), .A2(KEYINPUT70), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(KEYINPUT70), .ZN(new_n477));
  AOI211_X1 g276(.A(new_n472), .B(new_n474), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(G183gat), .A2(G190gat), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  NOR3_X1   g279(.A1(new_n470), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT23), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n473), .B1(new_n472), .B2(new_n482), .ZN(new_n483));
  XNOR2_X1  g282(.A(KEYINPUT65), .B(G169gat), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n484), .A2(KEYINPUT23), .A3(new_n294), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT64), .ZN(new_n486));
  OAI21_X1  g285(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(new_n479), .ZN(new_n488));
  NAND3_X1  g287(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n486), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  AND2_X1   g289(.A1(new_n489), .A2(new_n486), .ZN(new_n491));
  OAI211_X1 g290(.A(new_n483), .B(new_n485), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT25), .ZN(new_n493));
  AND3_X1   g292(.A1(new_n492), .A2(KEYINPUT66), .A3(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(KEYINPUT66), .B1(new_n492), .B2(new_n493), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n483), .B(KEYINPUT25), .C1(new_n482), .C2(new_n473), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n496), .B1(new_n489), .B2(new_n488), .ZN(new_n497));
  NOR3_X1   g296(.A1(new_n494), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n450), .B(new_n451), .C1(new_n481), .C2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n478), .ZN(new_n500));
  AND2_X1   g299(.A1(new_n468), .A2(new_n469), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n500), .B(new_n479), .C1(new_n501), .C2(new_n455), .ZN(new_n502));
  OR3_X1    g301(.A1(new_n494), .A2(new_n495), .A3(new_n497), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n502), .A2(new_n503), .A3(G226gat), .A4(G233gat), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n449), .B1(new_n499), .B2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT81), .ZN(new_n507));
  AND3_X1   g306(.A1(new_n442), .A2(KEYINPUT80), .A3(new_n443), .ZN(new_n508));
  AOI21_X1  g307(.A(KEYINPUT80), .B1(new_n442), .B2(new_n443), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n446), .A2(KEYINPUT81), .A3(new_n447), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n499), .A2(new_n504), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n506), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(G8gat), .B(G36gat), .ZN(new_n515));
  INV_X1    g314(.A(G64gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n515), .B(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n517), .B(new_n233), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(KEYINPUT30), .B1(new_n514), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n506), .A2(new_n518), .A3(new_n513), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n514), .A2(KEYINPUT30), .A3(new_n519), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n406), .A2(new_n430), .A3(new_n431), .A4(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(KEYINPUT31), .B(G50gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n526), .B(G106gat), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n415), .A2(new_n450), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n510), .A2(new_n511), .A3(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(G228gat), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n531), .A2(new_n298), .ZN(new_n532));
  AOI21_X1  g331(.A(KEYINPUT29), .B1(new_n442), .B2(new_n443), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n378), .B1(new_n533), .B2(KEYINPUT3), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n530), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT89), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT89), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n530), .A2(new_n537), .A3(new_n532), .A4(new_n534), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G22gat), .B(G78gat), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n448), .A2(new_n529), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(KEYINPUT88), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT88), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n448), .A2(new_n544), .A3(new_n529), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n543), .A2(new_n534), .A3(new_n545), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n546), .B1(new_n531), .B2(new_n298), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n539), .A2(new_n541), .A3(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n541), .B1(new_n539), .B2(new_n547), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n528), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n550), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n552), .A2(new_n527), .A3(new_n548), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  XOR2_X1   g353(.A(KEYINPUT86), .B(KEYINPUT6), .Z(new_n555));
  NAND3_X1  g354(.A1(new_n428), .A2(new_n429), .A3(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT87), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n555), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n401), .B(new_n408), .C1(new_n426), .C2(new_n427), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n430), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT37), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n519), .B1(new_n514), .B2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT38), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n499), .A2(new_n504), .ZN(new_n565));
  OR3_X1    g364(.A1(new_n565), .A2(KEYINPUT90), .A3(new_n449), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n512), .ZN(new_n567));
  OAI21_X1  g366(.A(KEYINPUT90), .B1(new_n565), .B2(new_n449), .ZN(new_n568));
  AND3_X1   g367(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n563), .B(new_n564), .C1(new_n569), .C2(new_n562), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n428), .A2(KEYINPUT87), .A3(new_n429), .A4(new_n555), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n558), .A2(new_n561), .A3(new_n570), .A4(new_n571), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n563), .B1(new_n562), .B2(new_n514), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(KEYINPUT38), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n514), .A2(new_n519), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  OAI211_X1 g375(.A(new_n525), .B(new_n554), .C1(new_n572), .C2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n558), .A2(new_n561), .A3(new_n571), .ZN(new_n578));
  AND3_X1   g377(.A1(new_n523), .A2(KEYINPUT82), .A3(new_n522), .ZN(new_n579));
  AOI21_X1  g378(.A(KEYINPUT82), .B1(new_n523), .B2(new_n522), .ZN(new_n580));
  NOR3_X1   g379(.A1(new_n579), .A2(new_n580), .A3(new_n520), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n554), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT36), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n385), .A2(new_n375), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n585), .B1(new_n481), .B2(new_n498), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n502), .A2(new_n377), .A3(new_n503), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(G227gat), .A2(G233gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(KEYINPUT78), .B1(new_n590), .B2(KEYINPUT34), .ZN(new_n591));
  INV_X1    g390(.A(new_n589), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n592), .B1(new_n586), .B2(new_n587), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT78), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT34), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n590), .A2(KEYINPUT77), .A3(KEYINPUT34), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT77), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n598), .B1(new_n593), .B2(new_n595), .ZN(new_n599));
  AOI22_X1  g398(.A1(new_n591), .A2(new_n596), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n586), .A2(new_n587), .A3(new_n592), .ZN(new_n601));
  XNOR2_X1  g400(.A(G15gat), .B(G43gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(G71gat), .ZN(new_n603));
  INV_X1    g402(.A(G99gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(KEYINPUT33), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n601), .A2(KEYINPUT32), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n601), .A2(KEYINPUT32), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT76), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT33), .ZN(new_n610));
  AND3_X1   g409(.A1(new_n601), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n609), .B1(new_n601), .B2(new_n610), .ZN(new_n612));
  OAI211_X1 g411(.A(new_n608), .B(new_n605), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n600), .A2(new_n607), .A3(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n600), .B1(new_n607), .B2(new_n613), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n584), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n613), .A2(new_n607), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n591), .A2(new_n596), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n597), .A2(new_n599), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n622), .A2(KEYINPUT36), .A3(new_n614), .ZN(new_n623));
  AOI22_X1  g422(.A1(new_n582), .A2(new_n583), .B1(new_n617), .B2(new_n623), .ZN(new_n624));
  AND3_X1   g423(.A1(new_n622), .A2(new_n554), .A3(new_n614), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n625), .A2(new_n578), .A3(new_n581), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(KEYINPUT35), .ZN(new_n627));
  INV_X1    g426(.A(new_n524), .ZN(new_n628));
  XNOR2_X1  g427(.A(KEYINPUT91), .B(KEYINPUT35), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n625), .A2(new_n578), .A3(new_n628), .A4(new_n629), .ZN(new_n630));
  AOI22_X1  g429(.A1(new_n577), .A2(new_n624), .B1(new_n627), .B2(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n222), .A2(new_n281), .A3(new_n223), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n282), .B1(new_n220), .B2(new_n221), .ZN(new_n633));
  NAND2_X1  g432(.A1(G229gat), .A2(G233gat), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT18), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  OR3_X1    g436(.A1(new_n220), .A2(new_n221), .A3(new_n282), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(new_n633), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n634), .B(KEYINPUT13), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n632), .A2(KEYINPUT18), .A3(new_n633), .A4(new_n634), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n637), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n645));
  XNOR2_X1  g444(.A(G113gat), .B(G141gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(G169gat), .B(G197gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(KEYINPUT93), .B(KEYINPUT12), .ZN(new_n650));
  XOR2_X1   g449(.A(new_n649), .B(new_n650), .Z(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n644), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n637), .A2(new_n651), .A3(new_n642), .A4(new_n643), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n320), .B1(new_n631), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n582), .A2(new_n583), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n617), .A2(new_n623), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n577), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n627), .A2(new_n630), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n662), .A2(KEYINPUT97), .A3(new_n655), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n319), .B1(new_n657), .B2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n578), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(G1gat), .ZN(G1324gat));
  INV_X1    g466(.A(new_n664), .ZN(new_n668));
  OAI21_X1  g467(.A(G8gat), .B1(new_n668), .B2(new_n628), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT42), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n277), .A2(new_n280), .ZN(new_n671));
  NAND2_X1  g470(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n664), .A2(new_n524), .A3(new_n671), .A4(new_n672), .ZN(new_n673));
  AND3_X1   g472(.A1(new_n673), .A2(KEYINPUT105), .A3(new_n670), .ZN(new_n674));
  AOI21_X1  g473(.A(KEYINPUT105), .B1(new_n673), .B2(new_n670), .ZN(new_n675));
  OAI221_X1 g474(.A(new_n669), .B1(new_n670), .B2(new_n673), .C1(new_n674), .C2(new_n675), .ZN(G1325gat));
  INV_X1    g475(.A(new_n659), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n664), .A2(G15gat), .A3(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n615), .A2(new_n616), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n668), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n678), .B1(new_n681), .B2(G15gat), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n682), .B(KEYINPUT106), .Z(G1326gat));
  NAND2_X1  g482(.A1(new_n664), .A2(new_n583), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT43), .B(G22gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1327gat));
  INV_X1    g485(.A(new_n318), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n292), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  AOI211_X1 g488(.A(new_n264), .B(new_n689), .C1(new_n657), .C2(new_n663), .ZN(new_n690));
  INV_X1    g489(.A(G29gat), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n690), .A2(new_n691), .A3(new_n665), .ZN(new_n692));
  XOR2_X1   g491(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  OR2_X1    g493(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n692), .A2(new_n694), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n689), .A2(new_n656), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  AND3_X1   g497(.A1(new_n262), .A2(KEYINPUT109), .A3(new_n263), .ZN(new_n699));
  AOI21_X1  g498(.A(KEYINPUT109), .B1(new_n262), .B2(new_n263), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n701), .A2(KEYINPUT44), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT108), .ZN(new_n703));
  AND3_X1   g502(.A1(new_n660), .A2(new_n661), .A3(new_n703), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n703), .B1(new_n660), .B2(new_n661), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n702), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n264), .B1(new_n660), .B2(new_n661), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708));
  OAI21_X1  g507(.A(KEYINPUT110), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  OAI211_X1 g509(.A(KEYINPUT110), .B(new_n702), .C1(new_n704), .C2(new_n705), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n698), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  AND2_X1   g511(.A1(new_n712), .A2(new_n665), .ZN(new_n713));
  OAI211_X1 g512(.A(new_n695), .B(new_n696), .C1(new_n691), .C2(new_n713), .ZN(G1328gat));
  INV_X1    g513(.A(G36gat), .ZN(new_n715));
  AND3_X1   g514(.A1(new_n690), .A2(new_n715), .A3(new_n524), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT46), .ZN(new_n717));
  OR2_X1    g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n716), .A2(new_n717), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n712), .A2(new_n524), .ZN(new_n720));
  OAI211_X1 g519(.A(new_n718), .B(new_n719), .C1(new_n715), .C2(new_n720), .ZN(G1329gat));
  AOI21_X1  g520(.A(new_n689), .B1(new_n657), .B2(new_n663), .ZN(new_n722));
  INV_X1    g521(.A(G43gat), .ZN(new_n723));
  INV_X1    g522(.A(new_n264), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n722), .A2(new_n723), .A3(new_n679), .A4(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(KEYINPUT111), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT111), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n690), .A2(new_n727), .A3(new_n723), .A4(new_n679), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT112), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT47), .ZN(new_n731));
  INV_X1    g530(.A(new_n702), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n662), .A2(KEYINPUT108), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n631), .A2(new_n703), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT110), .ZN(new_n736));
  AND3_X1   g535(.A1(new_n577), .A2(new_n658), .A3(new_n659), .ZN(new_n737));
  AND3_X1   g536(.A1(new_n578), .A2(new_n628), .A3(new_n629), .ZN(new_n738));
  AOI22_X1  g537(.A1(new_n738), .A2(new_n625), .B1(new_n626), .B2(KEYINPUT35), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n724), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n736), .B1(new_n740), .B2(KEYINPUT44), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n711), .B1(new_n735), .B2(new_n741), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n742), .A2(new_n677), .A3(new_n697), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(G43gat), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n729), .A2(new_n730), .A3(new_n731), .A4(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n730), .A2(new_n731), .ZN(new_n746));
  NAND2_X1  g545(.A1(KEYINPUT112), .A2(KEYINPUT47), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n726), .A2(new_n728), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n723), .B1(new_n712), .B2(new_n677), .ZN(new_n749));
  OAI211_X1 g548(.A(new_n746), .B(new_n747), .C1(new_n748), .C2(new_n749), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n745), .A2(new_n750), .ZN(G1330gat));
  INV_X1    g550(.A(KEYINPUT48), .ZN(new_n752));
  INV_X1    g551(.A(G50gat), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n753), .B1(new_n712), .B2(new_n583), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n690), .A2(new_n753), .A3(new_n583), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n752), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT113), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n752), .B1(new_n756), .B2(KEYINPUT114), .ZN(new_n760));
  INV_X1    g559(.A(new_n754), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT114), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n755), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n760), .A2(new_n761), .A3(new_n763), .ZN(new_n764));
  OAI211_X1 g563(.A(KEYINPUT113), .B(new_n752), .C1(new_n754), .C2(new_n756), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n759), .A2(new_n764), .A3(new_n765), .ZN(G1331gat));
  AOI21_X1  g565(.A(new_n655), .B1(new_n733), .B2(new_n734), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n264), .A2(new_n292), .A3(new_n687), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n665), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g572(.A1(new_n770), .A2(new_n628), .ZN(new_n774));
  NOR2_X1   g573(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n775));
  AND2_X1   g574(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n774), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n777), .B1(new_n774), .B2(new_n775), .ZN(G1333gat));
  NAND3_X1  g577(.A1(new_n771), .A2(G71gat), .A3(new_n677), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n770), .A2(new_n680), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n779), .B1(G71gat), .B2(new_n780), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g581(.A1(new_n771), .A2(new_n583), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g583(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n292), .A2(new_n655), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n785), .B1(new_n740), .B2(new_n787), .ZN(new_n788));
  XNOR2_X1  g587(.A(KEYINPUT115), .B(KEYINPUT51), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n707), .A2(new_n786), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n578), .A2(new_n318), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n791), .A2(new_n232), .A3(new_n792), .ZN(new_n793));
  AND3_X1   g592(.A1(new_n742), .A2(new_n792), .A3(new_n786), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n793), .B1(new_n794), .B2(new_n232), .ZN(G1336gat));
  INV_X1    g594(.A(KEYINPUT116), .ZN(new_n796));
  OR2_X1    g595(.A1(new_n796), .A2(KEYINPUT52), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n742), .A2(new_n524), .A3(new_n687), .A4(new_n786), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(G92gat), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n796), .A2(KEYINPUT52), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n628), .A2(G92gat), .ZN(new_n801));
  AND3_X1   g600(.A1(new_n791), .A2(new_n687), .A3(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  AND4_X1   g602(.A1(new_n797), .A2(new_n799), .A3(new_n800), .A4(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n802), .B1(new_n798), .B2(G92gat), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n797), .B1(new_n805), .B2(new_n800), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n804), .A2(new_n806), .ZN(G1337gat));
  AND4_X1   g606(.A1(new_n677), .A2(new_n742), .A3(new_n687), .A4(new_n786), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n791), .A2(new_n687), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n679), .A2(new_n604), .ZN(new_n810));
  OAI22_X1  g609(.A1(new_n808), .A2(new_n604), .B1(new_n809), .B2(new_n810), .ZN(G1338gat));
  OR2_X1    g610(.A1(new_n554), .A2(G106gat), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n742), .A2(new_n583), .A3(new_n687), .A4(new_n786), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n813), .B1(G106gat), .B2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT53), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n815), .B(new_n816), .ZN(G1339gat));
  INV_X1    g616(.A(new_n700), .ZN(new_n818));
  OAI211_X1 g617(.A(new_n299), .B(new_n307), .C1(new_n311), .C2(KEYINPUT10), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n309), .A2(new_n819), .A3(KEYINPUT54), .ZN(new_n820));
  XOR2_X1   g619(.A(KEYINPUT117), .B(KEYINPUT54), .Z(new_n821));
  OAI211_X1 g620(.A(new_n300), .B(new_n821), .C1(new_n306), .C2(new_n308), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n820), .A2(new_n296), .A3(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT55), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n309), .A2(new_n312), .A3(new_n316), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n820), .A2(KEYINPUT55), .A3(new_n296), .A4(new_n822), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n825), .A2(new_n826), .A3(new_n655), .A4(new_n827), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n639), .A2(new_n641), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n634), .B1(new_n632), .B2(new_n633), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n649), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n654), .A2(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n832), .B1(new_n315), .B2(new_n317), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n828), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n262), .A2(KEYINPUT109), .A3(new_n263), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n818), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  AND4_X1   g635(.A1(new_n826), .A2(new_n825), .A3(new_n827), .A4(new_n832), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n837), .B1(new_n699), .B2(new_n700), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n292), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n319), .A2(new_n655), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n578), .A2(new_n524), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n625), .ZN(new_n845));
  OAI21_X1  g644(.A(G113gat), .B1(new_n845), .B2(new_n656), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n655), .A2(new_n326), .ZN(new_n847));
  XOR2_X1   g646(.A(new_n847), .B(KEYINPUT118), .Z(new_n848));
  OAI21_X1  g647(.A(new_n846), .B1(new_n845), .B2(new_n848), .ZN(G1340gat));
  NOR2_X1   g648(.A1(new_n845), .A2(new_n318), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n850), .B(new_n327), .ZN(G1341gat));
  INV_X1    g650(.A(new_n292), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n845), .A2(new_n852), .ZN(new_n853));
  XOR2_X1   g652(.A(new_n853), .B(G127gat), .Z(G1342gat));
  NAND3_X1  g653(.A1(new_n844), .A2(new_n625), .A3(new_n724), .ZN(new_n855));
  NOR2_X1   g654(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n856));
  AND2_X1   g655(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n858), .B1(new_n855), .B2(new_n856), .ZN(G1343gat));
  OAI21_X1  g658(.A(new_n583), .B1(new_n839), .B2(new_n840), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT57), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT119), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n834), .A2(new_n264), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n292), .B1(new_n838), .B2(new_n865), .ZN(new_n866));
  OAI211_X1 g665(.A(KEYINPUT57), .B(new_n583), .C1(new_n866), .C2(new_n840), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n860), .A2(KEYINPUT119), .A3(new_n861), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n864), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n843), .A2(new_n677), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n869), .A2(new_n655), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(G141gat), .ZN(new_n872));
  INV_X1    g671(.A(new_n860), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n870), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n875), .A2(new_n354), .A3(new_n655), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(KEYINPUT58), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT58), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n872), .A2(new_n879), .A3(new_n876), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n878), .A2(new_n880), .ZN(G1344gat));
  NAND2_X1  g680(.A1(new_n724), .A2(new_n837), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n292), .B1(new_n865), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n861), .B1(new_n883), .B2(new_n840), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n884), .A2(new_n554), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n885), .B1(KEYINPUT57), .B2(new_n860), .ZN(new_n886));
  AND3_X1   g685(.A1(new_n886), .A2(new_n687), .A3(new_n870), .ZN(new_n887));
  OAI21_X1  g686(.A(KEYINPUT59), .B1(new_n887), .B2(new_n356), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT59), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n869), .A2(new_n870), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n889), .B1(new_n890), .B2(new_n318), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n888), .B1(new_n891), .B2(new_n356), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n875), .A2(new_n356), .A3(new_n687), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(G1345gat));
  AND3_X1   g693(.A1(new_n875), .A2(KEYINPUT120), .A3(new_n292), .ZN(new_n895));
  AOI21_X1  g694(.A(KEYINPUT120), .B1(new_n875), .B2(new_n292), .ZN(new_n896));
  NOR3_X1   g695(.A1(new_n895), .A2(new_n896), .A3(G155gat), .ZN(new_n897));
  INV_X1    g696(.A(new_n890), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n292), .A2(G155gat), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n897), .B1(new_n898), .B2(new_n899), .ZN(G1346gat));
  AOI21_X1  g699(.A(G162gat), .B1(new_n875), .B2(new_n724), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n701), .A2(new_n249), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n901), .B1(new_n898), .B2(new_n902), .ZN(G1347gat));
  OR2_X1    g702(.A1(new_n839), .A2(new_n840), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n665), .A2(new_n628), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n904), .A2(new_n625), .A3(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n907), .A2(new_n655), .A3(new_n484), .ZN(new_n908));
  XOR2_X1   g707(.A(new_n905), .B(KEYINPUT121), .Z(new_n909));
  NAND3_X1  g708(.A1(new_n904), .A2(new_n625), .A3(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT122), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n904), .A2(KEYINPUT122), .A3(new_n625), .A4(new_n909), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n914), .A2(new_n655), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n908), .B1(new_n915), .B2(new_n471), .ZN(G1348gat));
  AOI21_X1  g715(.A(G176gat), .B1(new_n907), .B2(new_n687), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n318), .A2(new_n294), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n917), .B1(new_n914), .B2(new_n918), .ZN(G1349gat));
  INV_X1    g718(.A(KEYINPUT123), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n920), .A2(KEYINPUT60), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n920), .A2(KEYINPUT60), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n912), .A2(new_n292), .A3(new_n913), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(G183gat), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n907), .A2(new_n452), .A3(new_n292), .ZN(new_n925));
  AOI211_X1 g724(.A(new_n921), .B(new_n922), .C1(new_n924), .C2(new_n925), .ZN(new_n926));
  AND4_X1   g725(.A1(new_n920), .A2(new_n924), .A3(KEYINPUT60), .A4(new_n925), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n926), .A2(new_n927), .ZN(G1350gat));
  INV_X1    g727(.A(new_n701), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n907), .A2(new_n453), .A3(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT61), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n914), .A2(new_n724), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n931), .B1(new_n932), .B2(G190gat), .ZN(new_n933));
  AOI211_X1 g732(.A(KEYINPUT61), .B(new_n453), .C1(new_n914), .C2(new_n724), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n930), .B1(new_n933), .B2(new_n934), .ZN(G1351gat));
  XNOR2_X1  g734(.A(KEYINPUT124), .B(G197gat), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n909), .A2(new_n659), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n886), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n936), .B1(new_n938), .B2(new_n656), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n905), .A2(new_n659), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n904), .A2(new_n583), .A3(new_n940), .ZN(new_n941));
  OR2_X1    g740(.A1(new_n656), .A2(new_n936), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n939), .B1(new_n941), .B2(new_n942), .ZN(G1352gat));
  INV_X1    g742(.A(new_n941), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(new_n687), .ZN(new_n945));
  XOR2_X1   g744(.A(KEYINPUT125), .B(G204gat), .Z(new_n946));
  OAI211_X1 g745(.A(KEYINPUT126), .B(KEYINPUT62), .C1(new_n945), .C2(new_n946), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n886), .A2(new_n687), .A3(new_n937), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(new_n946), .ZN(new_n949));
  NAND2_X1  g748(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n941), .A2(new_n318), .A3(new_n946), .ZN(new_n951));
  NOR2_X1   g750(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n950), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n947), .A2(new_n949), .A3(new_n953), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT127), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND4_X1  g755(.A1(new_n947), .A2(new_n949), .A3(new_n953), .A4(KEYINPUT127), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(G1353gat));
  NAND3_X1  g757(.A1(new_n944), .A2(new_n290), .A3(new_n292), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n886), .A2(new_n292), .A3(new_n937), .ZN(new_n960));
  AND3_X1   g759(.A1(new_n960), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n961));
  AOI21_X1  g760(.A(KEYINPUT63), .B1(new_n960), .B2(G211gat), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n959), .B1(new_n961), .B2(new_n962), .ZN(G1354gat));
  NOR3_X1   g762(.A1(new_n938), .A2(new_n433), .A3(new_n264), .ZN(new_n964));
  AOI21_X1  g763(.A(G218gat), .B1(new_n944), .B2(new_n929), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n964), .A2(new_n965), .ZN(G1355gat));
endmodule


