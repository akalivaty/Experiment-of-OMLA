//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 0 1 0 0 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 0 1 1 1 0 0 0 1 1 1 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:47 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n903, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966;
  INV_X1    g000(.A(G953), .ZN(new_n187));
  AND2_X1   g001(.A1(new_n187), .A2(G952), .ZN(new_n188));
  NAND2_X1  g002(.A1(G234), .A2(G237), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  XOR2_X1   g004(.A(new_n190), .B(KEYINPUT97), .Z(new_n191));
  AND3_X1   g005(.A1(new_n189), .A2(G902), .A3(G953), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT21), .B(G898), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  AND2_X1   g008(.A1(new_n191), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  NOR2_X1   g010(.A1(G475), .A2(G902), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  AOI21_X1  g012(.A(KEYINPUT20), .B1(new_n198), .B2(KEYINPUT93), .ZN(new_n199));
  OR2_X1    g013(.A1(new_n198), .A2(KEYINPUT93), .ZN(new_n200));
  AND2_X1   g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  XNOR2_X1  g016(.A(G113), .B(G122), .ZN(new_n203));
  INV_X1    g017(.A(G104), .ZN(new_n204));
  XNOR2_X1  g018(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G237), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(new_n187), .A3(G214), .ZN(new_n207));
  INV_X1    g021(.A(G143), .ZN(new_n208));
  XNOR2_X1  g022(.A(new_n207), .B(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(KEYINPUT18), .A2(G131), .ZN(new_n210));
  XNOR2_X1  g024(.A(new_n209), .B(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(G125), .A2(G140), .ZN(new_n212));
  XNOR2_X1  g026(.A(KEYINPUT79), .B(G125), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n212), .B1(new_n213), .B2(G140), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G146), .ZN(new_n215));
  XOR2_X1   g029(.A(G125), .B(G140), .Z(new_n216));
  OR2_X1    g030(.A1(new_n216), .A2(G146), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n211), .A2(new_n218), .ZN(new_n219));
  AND2_X1   g033(.A1(KEYINPUT66), .A2(G131), .ZN(new_n220));
  NOR2_X1   g034(.A1(KEYINPUT66), .A2(G131), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  XNOR2_X1  g037(.A(new_n209), .B(new_n223), .ZN(new_n224));
  OR2_X1    g038(.A1(new_n224), .A2(KEYINPUT17), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n209), .A2(KEYINPUT17), .A3(new_n223), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G146), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT16), .ZN(new_n229));
  AND2_X1   g043(.A1(KEYINPUT79), .A2(G125), .ZN(new_n230));
  NOR2_X1   g044(.A1(KEYINPUT79), .A2(G125), .ZN(new_n231));
  OAI21_X1  g045(.A(G140), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n212), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n229), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G140), .ZN(new_n235));
  AND3_X1   g049(.A1(new_n213), .A2(new_n229), .A3(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n228), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT80), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n213), .A2(new_n229), .A3(new_n235), .ZN(new_n239));
  OAI211_X1 g053(.A(G146), .B(new_n239), .C1(new_n214), .C2(new_n229), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n237), .A2(new_n238), .A3(new_n240), .ZN(new_n241));
  OAI211_X1 g055(.A(KEYINPUT80), .B(new_n228), .C1(new_n234), .C2(new_n236), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n227), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT92), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n225), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  AOI211_X1 g059(.A(KEYINPUT92), .B(new_n227), .C1(new_n241), .C2(new_n242), .ZN(new_n246));
  OAI211_X1 g060(.A(new_n205), .B(new_n219), .C1(new_n245), .C2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT19), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n216), .A2(new_n248), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n249), .B1(new_n214), .B2(new_n248), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(new_n228), .ZN(new_n251));
  XNOR2_X1  g065(.A(new_n251), .B(KEYINPUT91), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT81), .ZN(new_n253));
  OR2_X1    g067(.A1(new_n240), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n240), .A2(new_n253), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n254), .A2(new_n255), .A3(new_n224), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n219), .B1(new_n252), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n205), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n202), .B1(new_n247), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n247), .A2(new_n259), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(new_n197), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n260), .B1(new_n262), .B2(KEYINPUT20), .ZN(new_n263));
  INV_X1    g077(.A(G475), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n219), .B1(new_n245), .B2(new_n246), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(new_n258), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(new_n247), .ZN(new_n267));
  INV_X1    g081(.A(G902), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n264), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(KEYINPUT94), .B1(new_n263), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n241), .A2(new_n242), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(new_n226), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(KEYINPUT92), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n243), .A2(new_n244), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n273), .A2(new_n274), .A3(new_n225), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n205), .B1(new_n275), .B2(new_n219), .ZN(new_n276));
  INV_X1    g090(.A(new_n247), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n268), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G475), .ZN(new_n279));
  INV_X1    g093(.A(new_n261), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n198), .B1(new_n247), .B2(new_n259), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT20), .ZN(new_n282));
  OAI22_X1  g096(.A1(new_n280), .A2(new_n202), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT94), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n279), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(G128), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n286), .A2(G143), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n208), .A2(G128), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(G134), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(G134), .B1(new_n287), .B2(new_n288), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OR2_X1    g107(.A1(new_n293), .A2(KEYINPUT95), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(KEYINPUT95), .ZN(new_n295));
  INV_X1    g109(.A(G107), .ZN(new_n296));
  INV_X1    g110(.A(G116), .ZN(new_n297));
  OR2_X1    g111(.A1(new_n297), .A2(G122), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n296), .B1(new_n298), .B2(KEYINPUT14), .ZN(new_n299));
  XNOR2_X1  g113(.A(G116), .B(G122), .ZN(new_n300));
  XNOR2_X1  g114(.A(new_n299), .B(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n294), .A2(new_n295), .A3(new_n301), .ZN(new_n302));
  AOI22_X1  g116(.A1(new_n289), .A2(new_n290), .B1(G107), .B2(new_n300), .ZN(new_n303));
  AND2_X1   g117(.A1(new_n287), .A2(KEYINPUT13), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n287), .A2(KEYINPUT13), .ZN(new_n305));
  NOR3_X1   g119(.A1(new_n304), .A2(new_n305), .A3(new_n288), .ZN(new_n306));
  OAI221_X1 g120(.A(new_n303), .B1(G107), .B2(new_n300), .C1(new_n306), .C2(new_n290), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n302), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(KEYINPUT9), .B(G234), .ZN(new_n309));
  INV_X1    g123(.A(G217), .ZN(new_n310));
  NOR3_X1   g124(.A1(new_n309), .A2(new_n310), .A3(G953), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT96), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n302), .A2(new_n307), .A3(new_n311), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n308), .A2(KEYINPUT96), .A3(new_n312), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n316), .A2(new_n268), .A3(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G478), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n319), .A2(KEYINPUT15), .ZN(new_n320));
  OR2_X1    g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n318), .A2(new_n320), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  AND4_X1   g138(.A1(new_n196), .A2(new_n270), .A3(new_n285), .A4(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(G214), .B1(G237), .B2(G902), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT5), .ZN(new_n328));
  INV_X1    g142(.A(G119), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n328), .A2(new_n329), .A3(G116), .ZN(new_n330));
  XOR2_X1   g144(.A(G116), .B(G119), .Z(new_n331));
  OAI211_X1 g145(.A(G113), .B(new_n330), .C1(new_n331), .C2(new_n328), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT2), .B(G113), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n332), .B1(new_n333), .B2(new_n331), .ZN(new_n334));
  OAI21_X1  g148(.A(KEYINPUT3), .B1(new_n204), .B2(G107), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT3), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n336), .A2(new_n296), .A3(G104), .ZN(new_n337));
  INV_X1    g151(.A(G101), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n204), .A2(G107), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n335), .A2(new_n337), .A3(new_n338), .A4(new_n339), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n204), .A2(G107), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n296), .A2(G104), .ZN(new_n342));
  OAI21_X1  g156(.A(G101), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  OR2_X1    g158(.A1(new_n334), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n333), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT68), .ZN(new_n347));
  XNOR2_X1  g161(.A(G116), .B(G119), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n346), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n331), .A2(new_n333), .A3(KEYINPUT68), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n335), .A2(new_n337), .A3(new_n339), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(G101), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n353), .A2(KEYINPUT4), .A3(new_n340), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT4), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n352), .A2(new_n355), .A3(G101), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n351), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n345), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g172(.A(G110), .B(G122), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n345), .A2(new_n357), .A3(new_n359), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n361), .A2(KEYINPUT6), .A3(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(KEYINPUT1), .B1(new_n208), .B2(G146), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n208), .A2(G146), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n228), .A2(G143), .ZN(new_n366));
  OAI211_X1 g180(.A(G128), .B(new_n364), .C1(new_n365), .C2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n228), .A2(G143), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n208), .A2(G146), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n368), .B(new_n369), .C1(KEYINPUT1), .C2(new_n286), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n371), .A2(new_n213), .ZN(new_n372));
  XNOR2_X1  g186(.A(G143), .B(G146), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT65), .ZN(new_n374));
  OAI211_X1 g188(.A(KEYINPUT0), .B(G128), .C1(new_n373), .C2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n368), .A2(new_n369), .ZN(new_n376));
  NAND2_X1  g190(.A1(KEYINPUT0), .A2(G128), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n376), .A2(KEYINPUT65), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  NOR3_X1   g193(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n373), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n372), .B1(new_n384), .B2(new_n213), .ZN(new_n385));
  INV_X1    g199(.A(G224), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n386), .A2(G953), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n387), .B(KEYINPUT88), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n385), .B(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT6), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n358), .A2(new_n390), .A3(new_n360), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n363), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n334), .B(new_n344), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n359), .B(KEYINPUT8), .ZN(new_n394));
  OAI21_X1  g208(.A(KEYINPUT7), .B1(new_n386), .B2(G953), .ZN(new_n395));
  AOI22_X1  g209(.A1(new_n393), .A2(new_n394), .B1(new_n385), .B2(new_n395), .ZN(new_n396));
  OR2_X1    g210(.A1(new_n387), .A2(KEYINPUT89), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n387), .A2(KEYINPUT89), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n397), .A2(KEYINPUT7), .A3(new_n398), .ZN(new_n399));
  OR3_X1    g213(.A1(new_n385), .A2(KEYINPUT90), .A3(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(KEYINPUT90), .B1(new_n385), .B2(new_n399), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n396), .A2(new_n400), .A3(new_n362), .A4(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n392), .A2(new_n268), .A3(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(G210), .B1(G237), .B2(G902), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n392), .A2(new_n268), .A3(new_n404), .A4(new_n402), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n327), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(G469), .ZN(new_n409));
  XNOR2_X1  g223(.A(G110), .B(G140), .ZN(new_n410));
  AND2_X1   g224(.A1(new_n187), .A2(G227), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n410), .B(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n354), .A2(new_n356), .ZN(new_n414));
  AOI22_X1  g228(.A1(new_n375), .A2(new_n378), .B1(new_n381), .B2(new_n382), .ZN(new_n415));
  OAI21_X1  g229(.A(KEYINPUT86), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT86), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n384), .A2(new_n417), .A3(new_n356), .A4(new_n354), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n367), .A2(new_n340), .A3(new_n343), .A4(new_n370), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT10), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n420), .B(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n419), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT69), .ZN(new_n425));
  OAI21_X1  g239(.A(KEYINPUT11), .B1(new_n290), .B2(G137), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT11), .ZN(new_n427));
  INV_X1    g241(.A(G137), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(new_n428), .A3(G134), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n290), .A2(G137), .ZN(new_n431));
  AND3_X1   g245(.A1(new_n430), .A2(new_n431), .A3(new_n222), .ZN(new_n432));
  INV_X1    g246(.A(G131), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n433), .B1(new_n430), .B2(new_n431), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n425), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n430), .A2(new_n431), .A3(new_n222), .ZN(new_n436));
  AOI22_X1  g250(.A1(new_n426), .A2(new_n429), .B1(new_n290), .B2(G137), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n436), .B(KEYINPUT69), .C1(new_n433), .C2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n424), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n419), .A2(new_n439), .A3(new_n423), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n413), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n436), .B1(new_n433), .B2(new_n437), .ZN(new_n444));
  INV_X1    g258(.A(new_n420), .ZN(new_n445));
  AOI22_X1  g259(.A1(new_n370), .A2(new_n367), .B1(new_n340), .B2(new_n343), .ZN(new_n446));
  OAI211_X1 g260(.A(KEYINPUT12), .B(new_n444), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n445), .A2(new_n446), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n439), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n447), .B1(new_n449), .B2(KEYINPUT12), .ZN(new_n450));
  AND3_X1   g264(.A1(new_n442), .A2(new_n450), .A3(new_n413), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n409), .B(new_n268), .C1(new_n443), .C2(new_n451), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n409), .A2(new_n268), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n442), .A2(new_n450), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n412), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n422), .B1(new_n416), .B2(new_n418), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n412), .B1(new_n457), .B2(new_n439), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n441), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n456), .A2(new_n459), .A3(G469), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n452), .A2(new_n454), .A3(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT87), .ZN(new_n462));
  OAI21_X1  g276(.A(G221), .B1(new_n309), .B2(G902), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n462), .B1(new_n461), .B2(new_n463), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AND3_X1   g281(.A1(new_n325), .A2(new_n408), .A3(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT28), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n435), .A2(new_n384), .A3(new_n438), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT67), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n431), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n290), .A2(KEYINPUT67), .A3(G137), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n472), .B(new_n473), .C1(new_n290), .C2(G137), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(G131), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n475), .A2(new_n370), .A3(new_n367), .A4(new_n436), .ZN(new_n476));
  AND3_X1   g290(.A1(new_n349), .A2(new_n350), .A3(KEYINPUT71), .ZN(new_n477));
  AOI21_X1  g291(.A(KEYINPUT71), .B1(new_n349), .B2(new_n350), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n469), .B1(new_n470), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(KEYINPUT73), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT73), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n482), .B(new_n469), .C1(new_n470), .C2(new_n479), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n435), .A2(new_n384), .A3(new_n438), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(KEYINPUT70), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT70), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n435), .A2(new_n384), .A3(new_n487), .A4(new_n438), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT71), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n351), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n349), .A2(new_n350), .A3(KEYINPUT71), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n432), .A2(new_n371), .ZN(new_n492));
  AOI22_X1  g306(.A1(new_n490), .A2(new_n491), .B1(new_n492), .B2(new_n475), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n486), .A2(new_n488), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n384), .A2(new_n444), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n476), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n351), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n469), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n484), .A2(new_n498), .ZN(new_n499));
  XOR2_X1   g313(.A(KEYINPUT72), .B(KEYINPUT27), .Z(new_n500));
  NAND3_X1  g314(.A1(new_n206), .A2(new_n187), .A3(G210), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n500), .B(new_n501), .ZN(new_n502));
  XNOR2_X1  g316(.A(KEYINPUT26), .B(G101), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n502), .B(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(KEYINPUT29), .B1(new_n499), .B2(new_n504), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n486), .A2(KEYINPUT30), .A3(new_n476), .A4(new_n488), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT30), .ZN(new_n507));
  AOI22_X1  g321(.A1(new_n496), .A2(new_n507), .B1(new_n349), .B2(new_n350), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n504), .B1(new_n509), .B2(new_n494), .ZN(new_n510));
  OR2_X1    g324(.A1(new_n510), .A2(KEYINPUT75), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(KEYINPUT75), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n505), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n486), .A2(new_n476), .A3(new_n488), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n477), .A2(new_n478), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n494), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(KEYINPUT28), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n504), .A2(KEYINPUT29), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n518), .A2(new_n483), .A3(new_n481), .A4(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n521), .A2(KEYINPUT76), .A3(new_n268), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT76), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n469), .B1(new_n516), .B2(new_n494), .ZN(new_n524));
  NOR3_X1   g338(.A1(new_n524), .A2(new_n484), .A3(new_n519), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n523), .B1(new_n525), .B2(G902), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n513), .A2(new_n522), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(G472), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT32), .ZN(new_n529));
  AND2_X1   g343(.A1(new_n506), .A2(new_n508), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n494), .A2(new_n504), .ZN(new_n531));
  OAI21_X1  g345(.A(KEYINPUT31), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n504), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n533), .B1(new_n484), .B2(new_n498), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT31), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n509), .A2(new_n535), .A3(new_n494), .A4(new_n504), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n532), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT74), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n532), .A2(new_n534), .A3(KEYINPUT74), .A4(new_n536), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(G472), .A2(G902), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n529), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n542), .ZN(new_n544));
  AOI211_X1 g358(.A(KEYINPUT32), .B(new_n544), .C1(new_n539), .C2(new_n540), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n528), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT85), .ZN(new_n547));
  XNOR2_X1  g361(.A(G119), .B(G128), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n548), .B(KEYINPUT77), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  XNOR2_X1  g364(.A(KEYINPUT24), .B(G110), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(KEYINPUT23), .B1(new_n286), .B2(G119), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n553), .B(KEYINPUT78), .C1(new_n329), .C2(G128), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n329), .A2(G128), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT78), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n555), .B1(new_n556), .B2(KEYINPUT23), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  OAI22_X1  g372(.A1(new_n550), .A2(new_n552), .B1(G110), .B2(new_n558), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n254), .A2(new_n559), .A3(new_n255), .A4(new_n217), .ZN(new_n560));
  AOI22_X1  g374(.A1(new_n550), .A2(new_n552), .B1(G110), .B2(new_n558), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n561), .A2(new_n241), .A3(new_n242), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  XNOR2_X1  g377(.A(KEYINPUT22), .B(G137), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n187), .A2(G221), .A3(G234), .ZN(new_n565));
  XOR2_X1   g379(.A(new_n564), .B(new_n565), .Z(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n560), .A2(new_n562), .A3(new_n566), .ZN(new_n569));
  AND2_X1   g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n310), .B1(G234), .B2(new_n268), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n571), .A2(G902), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n572), .B(KEYINPUT83), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT84), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n570), .A2(KEYINPUT84), .A3(new_n573), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n568), .A2(new_n268), .A3(new_n569), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT25), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n568), .A2(KEYINPUT25), .A3(new_n268), .A4(new_n569), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n581), .A2(KEYINPUT82), .A3(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n571), .B1(new_n581), .B2(KEYINPUT82), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n578), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  AND3_X1   g400(.A1(new_n546), .A2(new_n547), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n547), .B1(new_n546), .B2(new_n586), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n468), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n589), .B(G101), .ZN(G3));
  INV_X1    g404(.A(new_n583), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n576), .B(new_n577), .C1(new_n591), .C2(new_n584), .ZN(new_n592));
  NOR3_X1   g406(.A1(new_n465), .A2(new_n592), .A3(new_n466), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n544), .B1(new_n539), .B2(new_n540), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n541), .A2(new_n268), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n594), .B1(new_n595), .B2(G472), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  XOR2_X1   g411(.A(new_n597), .B(KEYINPUT98), .Z(new_n598));
  INV_X1    g412(.A(KEYINPUT33), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n316), .A2(new_n599), .A3(new_n317), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n313), .A2(KEYINPUT33), .A3(new_n315), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n319), .A2(G902), .ZN(new_n604));
  XNOR2_X1  g418(.A(KEYINPUT99), .B(G478), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  AOI22_X1  g420(.A1(new_n603), .A2(new_n604), .B1(new_n318), .B2(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n607), .B1(new_n270), .B2(new_n285), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n408), .A2(new_n196), .ZN(new_n609));
  AND2_X1   g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n598), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(KEYINPUT100), .ZN(new_n612));
  XOR2_X1   g426(.A(KEYINPUT34), .B(G104), .Z(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(G6));
  NAND2_X1  g428(.A1(new_n281), .A2(new_n282), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n262), .A2(KEYINPUT20), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n269), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  AND3_X1   g431(.A1(new_n609), .A2(new_n323), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n598), .A2(new_n618), .ZN(new_n619));
  XOR2_X1   g433(.A(KEYINPUT35), .B(G107), .Z(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G9));
  AND3_X1   g435(.A1(new_n419), .A2(new_n439), .A3(new_n423), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n439), .B1(new_n419), .B2(new_n423), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n412), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n458), .A2(new_n450), .ZN(new_n625));
  AOI211_X1 g439(.A(G469), .B(G902), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n460), .A2(new_n454), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n463), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(KEYINPUT87), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n567), .A2(KEYINPUT36), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n563), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n573), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n632), .B1(new_n591), .B2(new_n584), .ZN(new_n633));
  AND4_X1   g447(.A1(new_n408), .A2(new_n629), .A3(new_n464), .A4(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n634), .A2(new_n325), .A3(new_n596), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT37), .B(G110), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G12));
  INV_X1    g451(.A(G900), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n192), .A2(new_n638), .ZN(new_n639));
  AND2_X1   g453(.A1(new_n191), .A2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  AND3_X1   g455(.A1(new_n617), .A2(new_n323), .A3(new_n641), .ZN(new_n642));
  AND3_X1   g456(.A1(new_n546), .A2(new_n634), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(new_n286), .ZN(G30));
  XOR2_X1   g458(.A(new_n640), .B(KEYINPUT39), .Z(new_n645));
  NAND2_X1  g459(.A1(new_n467), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(KEYINPUT103), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT103), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n467), .A2(new_n648), .A3(new_n645), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT40), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n647), .A2(KEYINPUT40), .A3(new_n649), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n324), .B1(new_n270), .B2(new_n285), .ZN(new_n655));
  INV_X1    g469(.A(new_n633), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n655), .A2(new_n326), .A3(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(new_n657), .B(KEYINPUT102), .Z(new_n658));
  NAND2_X1  g472(.A1(new_n541), .A2(new_n542), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(KEYINPUT32), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n594), .A2(new_n529), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n509), .A2(new_n494), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n504), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n268), .B1(new_n517), .B2(new_n504), .ZN(new_n666));
  OAI21_X1  g480(.A(G472), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n662), .A2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT101), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n662), .A2(KEYINPUT101), .A3(new_n667), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AND2_X1   g486(.A1(new_n406), .A2(new_n407), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(KEYINPUT38), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n654), .A2(new_n658), .A3(new_n672), .A4(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G143), .ZN(G45));
  AOI211_X1 g491(.A(new_n640), .B(new_n607), .C1(new_n270), .C2(new_n285), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n546), .A2(new_n634), .A3(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT104), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n546), .A2(new_n634), .A3(new_n678), .A4(KEYINPUT104), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G146), .ZN(G48));
  AOI21_X1  g498(.A(G902), .B1(new_n624), .B2(new_n625), .ZN(new_n685));
  NAND2_X1  g499(.A1(KEYINPUT105), .A2(G469), .ZN(new_n686));
  OR2_X1    g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n685), .A2(new_n686), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n463), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n610), .A2(new_n546), .A3(new_n691), .A4(new_n586), .ZN(new_n692));
  XNOR2_X1  g506(.A(KEYINPUT41), .B(G113), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G15));
  NAND4_X1  g508(.A1(new_n546), .A2(new_n618), .A3(new_n586), .A4(new_n691), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G116), .ZN(G18));
  NAND4_X1  g510(.A1(new_n408), .A2(new_n463), .A3(new_n687), .A4(new_n688), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n656), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n546), .A2(new_n325), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G119), .ZN(G21));
  XNOR2_X1  g514(.A(new_n655), .B(KEYINPUT108), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n697), .A2(new_n195), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n533), .B1(new_n524), .B2(new_n484), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT106), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n703), .A2(new_n704), .A3(new_n532), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n536), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n704), .B1(new_n703), .B2(new_n532), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n542), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(G472), .ZN(new_n709));
  AOI21_X1  g523(.A(G902), .B1(new_n539), .B2(new_n540), .ZN(new_n710));
  OAI211_X1 g524(.A(new_n708), .B(new_n586), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT107), .ZN(new_n712));
  AND2_X1   g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n711), .A2(new_n712), .ZN(new_n714));
  OAI211_X1 g528(.A(new_n701), .B(new_n702), .C1(new_n713), .C2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G122), .ZN(G24));
  INV_X1    g530(.A(new_n697), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n608), .A2(new_n717), .A3(new_n641), .ZN(new_n718));
  OAI211_X1 g532(.A(new_n708), .B(new_n633), .C1(new_n709), .C2(new_n710), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT109), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n595), .A2(G472), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n722), .A2(KEYINPUT109), .A3(new_n633), .A4(new_n708), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n718), .B1(new_n721), .B2(new_n723), .ZN(new_n724));
  XOR2_X1   g538(.A(new_n724), .B(G125), .Z(G27));
  AOI21_X1  g539(.A(new_n592), .B1(new_n662), .B2(new_n528), .ZN(new_n726));
  NOR2_X1   g540(.A1(KEYINPUT110), .A2(KEYINPUT42), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n673), .A2(new_n326), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n729), .A2(new_n628), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n726), .A2(new_n678), .A3(new_n728), .A4(new_n730), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n546), .A2(new_n678), .A3(new_n586), .A4(new_n730), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n727), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G131), .ZN(G33));
  AND4_X1   g549(.A1(new_n546), .A2(new_n586), .A3(new_n642), .A4(new_n730), .ZN(new_n736));
  XNOR2_X1  g550(.A(KEYINPUT111), .B(G134), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n736), .B(new_n737), .ZN(G36));
  NOR2_X1   g552(.A1(new_n596), .A2(new_n656), .ZN(new_n739));
  XOR2_X1   g553(.A(new_n739), .B(KEYINPUT115), .Z(new_n740));
  INV_X1    g554(.A(new_n607), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n270), .A2(new_n285), .A3(new_n741), .ZN(new_n742));
  XOR2_X1   g556(.A(KEYINPUT114), .B(KEYINPUT43), .Z(new_n743));
  OR2_X1    g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(KEYINPUT114), .A2(KEYINPUT43), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n740), .A2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT44), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n729), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n456), .A2(new_n459), .A3(KEYINPUT45), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT112), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n752), .B(new_n753), .ZN(new_n754));
  AOI21_X1  g568(.A(KEYINPUT45), .B1(new_n456), .B2(new_n459), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n755), .A2(new_n409), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT113), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n754), .A2(KEYINPUT113), .A3(new_n756), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n453), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n761), .A2(KEYINPUT46), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n452), .B1(new_n761), .B2(KEYINPUT46), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n463), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n645), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n740), .A2(KEYINPUT44), .A3(new_n747), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n750), .A2(new_n751), .A3(new_n766), .A4(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G137), .ZN(G39));
  INV_X1    g583(.A(KEYINPUT47), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n764), .A2(new_n770), .ZN(new_n771));
  OAI211_X1 g585(.A(KEYINPUT47), .B(new_n463), .C1(new_n762), .C2(new_n763), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI22_X1  g587(.A1(new_n660), .A2(new_n661), .B1(G472), .B2(new_n527), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n586), .A2(new_n729), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n773), .A2(new_n774), .A3(new_n678), .A4(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G140), .ZN(G42));
  NOR3_X1   g591(.A1(new_n592), .A2(new_n327), .A3(new_n690), .ZN(new_n778));
  OR2_X1    g592(.A1(new_n689), .A2(KEYINPUT49), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n689), .A2(KEYINPUT49), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n778), .A2(new_n674), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  OR3_X1    g595(.A1(new_n672), .A2(new_n742), .A3(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n711), .B(new_n712), .ZN(new_n783));
  INV_X1    g597(.A(new_n191), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n783), .A2(new_n784), .A3(new_n747), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n717), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n751), .A2(new_n691), .A3(KEYINPUT117), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT117), .ZN(new_n788));
  INV_X1    g602(.A(new_n691), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n788), .B1(new_n789), .B2(new_n729), .ZN(new_n790));
  AND4_X1   g604(.A1(new_n784), .A2(new_n747), .A3(new_n787), .A4(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT48), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n791), .A2(new_n792), .A3(new_n726), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n792), .B1(new_n791), .B2(new_n726), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n188), .B(new_n786), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT118), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n790), .A2(new_n586), .A3(new_n784), .A4(new_n787), .ZN(new_n797));
  OR3_X1    g611(.A1(new_n672), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n796), .B1(new_n672), .B2(new_n797), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n798), .A2(new_n799), .A3(new_n608), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  OAI21_X1  g615(.A(KEYINPUT119), .B1(new_n795), .B2(new_n801), .ZN(new_n802));
  OAI211_X1 g616(.A(new_n771), .B(new_n772), .C1(new_n463), .C2(new_n689), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n785), .A2(new_n751), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT51), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n675), .A2(new_n326), .A3(new_n789), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n785), .A2(KEYINPUT50), .A3(new_n807), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n783), .A2(new_n784), .A3(new_n747), .A4(new_n807), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT50), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n806), .B1(new_n808), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n721), .A2(new_n723), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n791), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n270), .A2(new_n285), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n815), .A2(new_n741), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n798), .A2(new_n799), .A3(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n805), .A2(new_n812), .A3(new_n814), .A4(new_n817), .ZN(new_n818));
  OR2_X1    g632(.A1(new_n793), .A2(new_n794), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n786), .A2(new_n188), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT119), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n819), .A2(new_n800), .A3(new_n820), .A4(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n802), .A2(new_n818), .A3(new_n822), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n817), .A2(new_n814), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT116), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n805), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n803), .A2(KEYINPUT116), .A3(new_n804), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n808), .A2(new_n811), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n824), .A2(new_n826), .A3(new_n827), .A4(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n823), .B1(new_n806), .B2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT53), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n724), .A2(new_n643), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n633), .A2(new_n628), .A3(new_n640), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n701), .A2(new_n408), .A3(new_n668), .A4(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n832), .A2(new_n683), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(KEYINPUT52), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT52), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n832), .A2(new_n683), .A3(new_n837), .A4(new_n834), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n589), .A2(new_n715), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n692), .A2(new_n695), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n593), .A2(new_n596), .A3(new_n609), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n815), .A2(new_n607), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n843), .B1(new_n815), .B2(new_n323), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n699), .A2(new_n635), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n841), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n736), .B1(new_n731), .B2(new_n733), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n608), .A2(new_n463), .A3(new_n461), .A4(new_n641), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n849), .B1(new_n721), .B2(new_n723), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n323), .A2(new_n640), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n467), .A2(new_n617), .A3(new_n633), .A4(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n852), .A2(new_n774), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n751), .B1(new_n850), .B2(new_n853), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n840), .A2(new_n847), .A3(new_n848), .A4(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n831), .B1(new_n839), .B2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(new_n736), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n734), .A2(new_n854), .A3(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n846), .A2(new_n845), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n726), .B(new_n691), .C1(new_n610), .C2(new_n618), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n859), .A2(new_n589), .A3(new_n715), .A4(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n831), .B1(new_n832), .B2(new_n837), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n862), .A2(new_n836), .A3(new_n838), .A4(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n856), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(KEYINPUT54), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n832), .A2(new_n837), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n867), .A2(new_n831), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n862), .A2(new_n836), .A3(new_n838), .A4(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT54), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n856), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n830), .A2(new_n866), .A3(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(G952), .A2(G953), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n782), .B1(new_n872), .B2(new_n873), .ZN(G75));
  AOI21_X1  g688(.A(new_n268), .B1(new_n856), .B2(new_n869), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n875), .A2(KEYINPUT120), .A3(G210), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT56), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n363), .A2(new_n391), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(new_n389), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(KEYINPUT55), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n876), .A2(new_n877), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(KEYINPUT120), .B1(new_n875), .B2(G210), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n187), .A2(G952), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(KEYINPUT56), .B1(new_n875), .B2(G210), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n885), .B1(new_n886), .B2(new_n880), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n883), .A2(new_n887), .ZN(G51));
  XNOR2_X1  g702(.A(new_n453), .B(KEYINPUT57), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n856), .A2(new_n870), .A3(new_n869), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n870), .B1(new_n856), .B2(new_n869), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT121), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n624), .A2(new_n625), .ZN(new_n895));
  OAI211_X1 g709(.A(KEYINPUT121), .B(new_n889), .C1(new_n890), .C2(new_n891), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n875), .A2(new_n759), .A3(new_n760), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n884), .B1(new_n897), .B2(new_n898), .ZN(G54));
  NAND3_X1  g713(.A1(new_n875), .A2(KEYINPUT58), .A3(G475), .ZN(new_n900));
  OR3_X1    g714(.A1(new_n900), .A2(KEYINPUT122), .A3(new_n280), .ZN(new_n901));
  OAI21_X1  g715(.A(KEYINPUT122), .B1(new_n900), .B2(new_n280), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n884), .B1(new_n900), .B2(new_n280), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(G60));
  NAND2_X1  g718(.A1(G478), .A2(G902), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(KEYINPUT59), .Z(new_n906));
  AOI21_X1  g720(.A(new_n906), .B1(new_n866), .B2(new_n871), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n885), .B1(new_n907), .B2(new_n603), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n602), .A2(new_n906), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n909), .B1(new_n890), .B2(new_n891), .ZN(new_n910));
  OR2_X1    g724(.A1(new_n910), .A2(KEYINPUT123), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(KEYINPUT123), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n908), .B1(new_n911), .B2(new_n912), .ZN(G63));
  NAND2_X1  g727(.A1(G217), .A2(G902), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT60), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n915), .B1(new_n856), .B2(new_n869), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n884), .B1(new_n916), .B2(new_n631), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n570), .B(KEYINPUT124), .Z(new_n918));
  OAI21_X1  g732(.A(new_n917), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  XNOR2_X1  g733(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n919), .B(new_n921), .ZN(G66));
  OAI21_X1  g736(.A(G953), .B1(new_n193), .B2(new_n386), .ZN(new_n923));
  INV_X1    g737(.A(new_n861), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n923), .B1(new_n924), .B2(G953), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n878), .B1(G898), .B2(new_n187), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n925), .B(new_n926), .ZN(G69));
  NAND2_X1  g741(.A1(new_n768), .A2(new_n776), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n766), .A2(new_n726), .A3(new_n408), .A4(new_n701), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n832), .A2(new_n683), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n929), .A2(new_n848), .A3(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n928), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(new_n187), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n496), .A2(new_n507), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n506), .A2(new_n934), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(new_n250), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n936), .B1(G900), .B2(G953), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT127), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n187), .B1(G227), .B2(G900), .ZN(new_n939));
  AOI22_X1  g753(.A1(new_n933), .A2(new_n937), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT62), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n676), .A2(new_n941), .A3(new_n930), .ZN(new_n942));
  NOR3_X1   g756(.A1(new_n650), .A2(new_n729), .A3(new_n844), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n943), .B1(new_n588), .B2(new_n587), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n768), .A2(new_n776), .A3(new_n942), .A4(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n676), .A2(new_n930), .ZN(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(KEYINPUT126), .B1(new_n947), .B2(new_n941), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT126), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n946), .A2(new_n949), .A3(KEYINPUT62), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n945), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n936), .B1(new_n951), .B2(G953), .ZN(new_n952));
  OR2_X1    g766(.A1(new_n939), .A2(new_n938), .ZN(new_n953));
  AND3_X1   g767(.A1(new_n940), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n953), .B1(new_n940), .B2(new_n952), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n954), .A2(new_n955), .ZN(G72));
  NAND2_X1  g770(.A1(new_n951), .A2(new_n924), .ZN(new_n957));
  NAND2_X1  g771(.A1(G472), .A2(G902), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT63), .Z(new_n959));
  AOI21_X1  g773(.A(new_n664), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n511), .B(new_n512), .C1(new_n530), .C2(new_n531), .ZN(new_n961));
  AND3_X1   g775(.A1(new_n865), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n959), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n963), .B1(new_n932), .B2(new_n924), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n509), .A2(new_n494), .A3(new_n533), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n885), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n960), .A2(new_n962), .A3(new_n966), .ZN(G57));
endmodule


