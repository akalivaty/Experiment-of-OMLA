//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 0 0 1 0 0 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 0 1 0 0 1 0 1 0 0 0 0 0 1 1 1 1 1 1 0 1 1 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:44 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1348, new_n1349;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  AOI22_X1  g0009(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n210));
  INV_X1    g0010(.A(G226), .ZN(new_n211));
  XOR2_X1   g0011(.A(KEYINPUT64), .B(G238), .Z(new_n212));
  INV_X1    g0012(.A(G68), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n210), .B1(new_n202), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n215));
  XOR2_X1   g0015(.A(new_n215), .B(KEYINPUT65), .Z(new_n216));
  NOR2_X1   g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G58), .A2(G232), .ZN(new_n218));
  INV_X1    g0018(.A(G107), .ZN(new_n219));
  INV_X1    g0019(.A(G264), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n217), .B(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(new_n206), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT1), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(new_n201), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(G50), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  AOI211_X1 g0029(.A(new_n209), .B(new_n223), .C1(new_n226), .C2(new_n229), .ZN(G361));
  XOR2_X1   g0030(.A(G226), .B(G232), .Z(new_n231));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G250), .B(G257), .Z(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n235), .B(new_n238), .Z(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  XNOR2_X1  g0046(.A(KEYINPUT3), .B(G33), .ZN(new_n247));
  XNOR2_X1  g0047(.A(KEYINPUT67), .B(G1698), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n247), .A2(new_n248), .A3(G232), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n247), .A2(G1698), .ZN(new_n250));
  OAI221_X1 g0050(.A(new_n249), .B1(new_n219), .B2(new_n247), .C1(new_n212), .C2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  INV_X1    g0052(.A(G41), .ZN(new_n253));
  OAI211_X1 g0053(.A(G1), .B(G13), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n251), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G1), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n257), .B1(G41), .B2(G45), .ZN(new_n258));
  INV_X1    g0058(.A(G274), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n254), .A2(new_n258), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G244), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n256), .A2(new_n261), .A3(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G179), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(KEYINPUT68), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT68), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G179), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n266), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G169), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n265), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G13), .ZN(new_n275));
  NOR3_X1   g0075(.A1(new_n275), .A2(new_n225), .A3(G1), .ZN(new_n276));
  INV_X1    g0076(.A(G77), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(new_n278), .B(KEYINPUT69), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n224), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n225), .A2(G1), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT8), .B(G58), .ZN(new_n285));
  NOR2_X1   g0085(.A1(G20), .A2(G33), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  OAI22_X1  g0087(.A1(new_n285), .A2(new_n287), .B1(new_n225), .B2(new_n277), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n252), .A2(G20), .ZN(new_n289));
  XOR2_X1   g0089(.A(KEYINPUT15), .B(G87), .Z(new_n290));
  AOI21_X1  g0090(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n281), .ZN(new_n292));
  OAI221_X1 g0092(.A(new_n279), .B1(new_n277), .B2(new_n284), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n272), .A2(new_n274), .A3(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n285), .A2(new_n282), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n295), .B(KEYINPUT77), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n276), .A2(new_n281), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n296), .A2(new_n297), .B1(new_n276), .B2(new_n285), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  XNOR2_X1  g0099(.A(G58), .B(G68), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n300), .A2(G20), .B1(G159), .B2(new_n286), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT3), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G33), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n306), .A2(KEYINPUT7), .A3(new_n225), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT76), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n304), .A2(G33), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n308), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n303), .A2(new_n305), .A3(KEYINPUT76), .ZN(new_n312));
  AOI21_X1  g0112(.A(G20), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n307), .B1(new_n313), .B2(KEYINPUT7), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n302), .B1(new_n314), .B2(G68), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n292), .B1(new_n315), .B2(KEYINPUT16), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT16), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT7), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n318), .B1(new_n247), .B2(G20), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n213), .B1(new_n319), .B2(new_n307), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n317), .B1(new_n320), .B2(new_n302), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n299), .B1(new_n316), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT78), .ZN(new_n323));
  AND2_X1   g0123(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n324));
  NOR2_X1   g0124(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n325));
  OAI21_X1  g0125(.A(G223), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n323), .B1(new_n326), .B2(new_n306), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n247), .A2(new_n248), .A3(KEYINPUT78), .A4(G223), .ZN(new_n328));
  NAND2_X1  g0128(.A1(G33), .A2(G87), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n247), .A2(G226), .A3(G1698), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n327), .A2(new_n328), .A3(new_n329), .A4(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n255), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n263), .A2(G232), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n332), .A2(G190), .A3(new_n261), .A4(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n332), .A2(new_n261), .A3(new_n333), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(G200), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n322), .A2(KEYINPUT17), .A3(new_n334), .A4(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n307), .ZN(new_n338));
  AND3_X1   g0138(.A1(new_n303), .A2(new_n305), .A3(KEYINPUT76), .ZN(new_n339));
  AOI21_X1  g0139(.A(KEYINPUT76), .B1(new_n303), .B2(new_n305), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n225), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n338), .B1(new_n341), .B2(new_n318), .ZN(new_n342));
  OAI211_X1 g0142(.A(KEYINPUT16), .B(new_n301), .C1(new_n342), .C2(new_n213), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n343), .A2(new_n281), .A3(new_n321), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n344), .A2(new_n336), .A3(new_n334), .A4(new_n298), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT17), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n344), .A2(new_n298), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n335), .A2(G169), .ZN(new_n349));
  INV_X1    g0149(.A(new_n271), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n332), .A2(new_n261), .A3(new_n350), .A4(new_n333), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  AND3_X1   g0152(.A1(new_n348), .A2(KEYINPUT18), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(KEYINPUT18), .B1(new_n348), .B2(new_n352), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n337), .B(new_n347), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(KEYINPUT79), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n289), .A2(G77), .ZN(new_n357));
  OAI221_X1 g0157(.A(new_n357), .B1(new_n225), .B2(G68), .C1(new_n202), .C2(new_n287), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n281), .ZN(new_n359));
  XOR2_X1   g0159(.A(new_n359), .B(KEYINPUT11), .Z(new_n360));
  NAND2_X1  g0160(.A1(new_n282), .A2(G13), .ZN(new_n361));
  NOR3_X1   g0161(.A1(new_n361), .A2(KEYINPUT12), .A3(G68), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT12), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n363), .B1(new_n276), .B2(new_n213), .ZN(new_n364));
  OAI22_X1  g0164(.A1(new_n362), .A2(new_n364), .B1(new_n284), .B2(new_n213), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n360), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT74), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT13), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n303), .A2(new_n305), .A3(G226), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n324), .A2(new_n325), .ZN(new_n371));
  OAI21_X1  g0171(.A(KEYINPUT70), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT70), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n247), .A2(new_n248), .A3(new_n373), .A4(G226), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT71), .ZN(new_n375));
  INV_X1    g0175(.A(G97), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n375), .B1(new_n252), .B2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(KEYINPUT71), .A2(G33), .A3(G97), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n247), .A2(G232), .A3(G1698), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n372), .A2(new_n374), .A3(new_n379), .A4(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(new_n255), .ZN(new_n382));
  INV_X1    g0182(.A(G238), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n261), .B1(new_n262), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n369), .B1(new_n382), .B2(new_n385), .ZN(new_n386));
  AOI211_X1 g0186(.A(KEYINPUT13), .B(new_n384), .C1(new_n381), .C2(new_n255), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n368), .B1(new_n388), .B2(G179), .ZN(new_n389));
  NOR4_X1   g0189(.A1(new_n386), .A2(new_n387), .A3(KEYINPUT74), .A4(new_n267), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n382), .A2(new_n385), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(KEYINPUT13), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT72), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n384), .B1(new_n381), .B2(new_n255), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n394), .B1(new_n395), .B2(new_n369), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n392), .A2(new_n394), .A3(KEYINPUT13), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n397), .A2(G169), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(KEYINPUT14), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT14), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n397), .A2(new_n401), .A3(G169), .A4(new_n398), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n391), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n397), .A2(G200), .A3(new_n398), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n388), .A2(G190), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n404), .A2(new_n405), .A3(new_n366), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT73), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n404), .A2(KEYINPUT73), .A3(new_n405), .A4(new_n366), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n367), .A2(new_n403), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT75), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n294), .B(new_n356), .C1(new_n410), .C2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n266), .A2(G190), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n293), .B1(new_n265), .B2(G200), .ZN(new_n414));
  AND2_X1   g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n403), .A2(new_n367), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n408), .A2(new_n409), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n416), .B1(new_n419), .B2(KEYINPUT75), .ZN(new_n420));
  XOR2_X1   g0220(.A(KEYINPUT8), .B(G58), .Z(new_n421));
  AOI22_X1  g0221(.A1(new_n421), .A2(new_n289), .B1(G150), .B2(new_n286), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n203), .A2(G20), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n424), .A2(new_n281), .B1(new_n202), .B2(new_n276), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n283), .A2(G50), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g0227(.A(new_n427), .B(KEYINPUT9), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n248), .A2(G222), .B1(G223), .B2(G1698), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n254), .B1(new_n429), .B2(new_n247), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n430), .B1(G77), .B2(new_n247), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n431), .B(new_n261), .C1(new_n211), .C2(new_n262), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(G200), .ZN(new_n433));
  INV_X1    g0233(.A(G190), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n428), .B(new_n433), .C1(new_n434), .C2(new_n432), .ZN(new_n435));
  XNOR2_X1  g0235(.A(new_n435), .B(KEYINPUT10), .ZN(new_n436));
  AND2_X1   g0236(.A1(new_n432), .A2(new_n273), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n427), .B1(new_n432), .B2(new_n350), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n436), .A2(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n355), .A2(KEYINPUT79), .ZN(new_n442));
  NOR4_X1   g0242(.A1(new_n412), .A2(new_n420), .A3(new_n441), .A4(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT4), .ZN(new_n444));
  OAI21_X1  g0244(.A(G244), .B1(new_n324), .B2(new_n325), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n444), .B1(new_n445), .B2(new_n306), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n247), .A2(new_n248), .A3(KEYINPUT4), .A4(G244), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n247), .A2(G250), .A3(G1698), .ZN(new_n448));
  NAND2_X1  g0248(.A1(G33), .A2(G283), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n446), .A2(new_n447), .A3(new_n448), .A4(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n255), .ZN(new_n451));
  OR2_X1    g0251(.A1(new_n253), .A2(KEYINPUT5), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n253), .A2(KEYINPUT5), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n452), .A2(new_n257), .A3(G45), .A4(new_n453), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n454), .A2(new_n254), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(G257), .ZN(new_n456));
  OR2_X1    g0256(.A1(new_n454), .A2(new_n259), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n451), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n273), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n361), .A2(G97), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n292), .B(new_n361), .C1(G1), .C2(new_n252), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n462), .A2(new_n376), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n219), .B1(new_n319), .B2(new_n307), .ZN(new_n465));
  XNOR2_X1  g0265(.A(KEYINPUT80), .B(G97), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n466), .A2(KEYINPUT6), .A3(new_n219), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT6), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n376), .A2(new_n219), .ZN(new_n469));
  NOR2_X1   g0269(.A1(G97), .A2(G107), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n225), .B1(new_n467), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n287), .A2(new_n277), .ZN(new_n473));
  NOR3_X1   g0273(.A1(new_n465), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n461), .B(new_n464), .C1(new_n474), .C2(new_n292), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n451), .A2(new_n271), .A3(new_n456), .A4(new_n457), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n459), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT81), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n458), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n451), .A2(KEYINPUT81), .A3(new_n456), .A4(new_n457), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n479), .A2(G200), .A3(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n475), .ZN(new_n482));
  AND3_X1   g0282(.A1(new_n451), .A2(new_n456), .A3(new_n457), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(G190), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n481), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n378), .ZN(new_n486));
  AOI21_X1  g0286(.A(KEYINPUT71), .B1(G33), .B2(G97), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT19), .ZN(new_n488));
  NOR3_X1   g0288(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  OAI21_X1  g0289(.A(KEYINPUT82), .B1(new_n489), .B2(G20), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT82), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n491), .B(new_n225), .C1(new_n379), .C2(new_n488), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n376), .A2(KEYINPUT80), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT80), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G97), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(G87), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n496), .A2(new_n497), .A3(new_n219), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n490), .A2(new_n492), .A3(new_n498), .ZN(new_n499));
  NOR3_X1   g0299(.A1(new_n306), .A2(G20), .A3(new_n213), .ZN(new_n500));
  AOI21_X1  g0300(.A(KEYINPUT19), .B1(new_n466), .B2(new_n289), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n281), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n290), .A2(new_n361), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n290), .ZN(new_n507));
  OR2_X1    g0307(.A1(new_n462), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n504), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(G45), .ZN(new_n510));
  NOR3_X1   g0310(.A1(new_n510), .A2(new_n259), .A3(G1), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n254), .B(G250), .C1(G1), .C2(new_n510), .ZN(new_n513));
  NAND2_X1  g0313(.A1(G33), .A2(G116), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(G244), .A2(G1698), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n516), .B1(new_n371), .B2(new_n383), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n515), .B1(new_n517), .B2(new_n247), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n512), .B(new_n513), .C1(new_n518), .C2(new_n254), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n271), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n273), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n509), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n505), .B1(new_n503), .B2(new_n281), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n462), .A2(new_n497), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n519), .A2(G200), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n248), .A2(G238), .B1(G244), .B2(G1698), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n514), .B1(new_n528), .B2(new_n306), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n511), .B1(new_n529), .B2(new_n255), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n530), .A2(G190), .A3(new_n513), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n524), .A2(new_n526), .A3(new_n527), .A4(new_n531), .ZN(new_n532));
  AND4_X1   g0332(.A1(new_n477), .A2(new_n485), .A3(new_n523), .A4(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n276), .A2(KEYINPUT25), .A3(new_n219), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(KEYINPUT25), .B1(new_n276), .B2(new_n219), .ZN(new_n536));
  OAI22_X1  g0336(.A1(new_n462), .A2(new_n219), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n303), .A2(new_n305), .A3(new_n225), .A4(G87), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT83), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(KEYINPUT22), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n247), .A2(new_n225), .A3(G87), .A4(new_n541), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n514), .A2(G20), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n225), .A2(G107), .ZN(new_n548));
  XNOR2_X1  g0348(.A(new_n548), .B(KEYINPUT23), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n545), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(KEYINPUT24), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n546), .B1(new_n543), .B2(new_n544), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT24), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n552), .A2(new_n553), .A3(new_n549), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(KEYINPUT84), .B1(new_n555), .B2(new_n281), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT84), .ZN(new_n557));
  AOI211_X1 g0357(.A(new_n557), .B(new_n292), .C1(new_n551), .C2(new_n554), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n538), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n454), .A2(G264), .A3(new_n254), .ZN(new_n560));
  INV_X1    g0360(.A(G294), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n252), .A2(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(G250), .B1(new_n324), .B2(new_n325), .ZN(new_n563));
  NAND2_X1  g0363(.A1(G257), .A2(G1698), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n562), .B1(new_n565), .B2(new_n247), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n457), .B(new_n560), .C1(new_n566), .C2(new_n254), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n273), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(G179), .B2(new_n567), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n559), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(G200), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n567), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(KEYINPUT85), .ZN(new_n574));
  OR2_X1    g0374(.A1(new_n567), .A2(G190), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT85), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n567), .A2(new_n576), .A3(new_n572), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n574), .A2(new_n575), .A3(new_n577), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n578), .B(new_n538), .C1(new_n556), .C2(new_n558), .ZN(new_n579));
  AND2_X1   g0379(.A1(new_n571), .A2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(G116), .ZN(new_n581));
  OR2_X1    g0381(.A1(new_n462), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n276), .A2(new_n581), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n225), .B(new_n449), .C1(new_n496), .C2(G33), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n280), .A2(new_n224), .B1(G20), .B2(new_n581), .ZN(new_n585));
  AND3_X1   g0385(.A1(new_n584), .A2(KEYINPUT20), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(KEYINPUT20), .B1(new_n584), .B2(new_n585), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n582), .B(new_n583), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n247), .A2(new_n248), .A3(G257), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n306), .A2(G303), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n589), .B(new_n590), .C1(new_n220), .C2(new_n250), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n255), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n455), .A2(G270), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n592), .A2(new_n457), .A3(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n588), .A2(new_n594), .A3(G169), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT21), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AND3_X1   g0397(.A1(new_n592), .A2(new_n457), .A3(new_n593), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n598), .A2(G179), .A3(new_n588), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n588), .A2(new_n594), .A3(KEYINPUT21), .A4(G169), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n597), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n588), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n594), .A2(new_n434), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n603), .B1(G200), .B2(new_n594), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n601), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  AND4_X1   g0405(.A1(new_n443), .A2(new_n533), .A3(new_n580), .A4(new_n605), .ZN(G372));
  INV_X1    g0406(.A(KEYINPUT87), .ZN(new_n607));
  AND3_X1   g0407(.A1(new_n552), .A2(new_n553), .A3(new_n549), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n553), .B1(new_n552), .B2(new_n549), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n281), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n557), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n555), .A2(KEYINPUT84), .A3(new_n281), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n537), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n607), .B1(new_n613), .B2(new_n569), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n559), .A2(KEYINPUT87), .A3(new_n570), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n597), .A2(new_n599), .A3(new_n600), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n523), .A2(new_n532), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(KEYINPUT86), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT86), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n523), .A2(new_n620), .A3(new_n532), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n579), .A2(new_n477), .A3(new_n485), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n617), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT88), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n523), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n509), .A2(new_n521), .A3(KEYINPUT88), .A4(new_n522), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT26), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n477), .A2(KEYINPUT89), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT89), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n459), .A2(new_n475), .A3(new_n631), .A4(new_n476), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n622), .A2(new_n629), .A3(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(KEYINPUT26), .B1(new_n618), .B2(new_n477), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n624), .A2(new_n628), .A3(new_n634), .A4(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n443), .A2(new_n636), .ZN(new_n637));
  OR2_X1    g0437(.A1(new_n353), .A2(new_n354), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n294), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n418), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n417), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n337), .A2(new_n347), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n639), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n436), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n440), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n637), .A2(new_n647), .ZN(G369));
  NOR2_X1   g0448(.A1(new_n275), .A2(G20), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n257), .ZN(new_n650));
  OR2_X1    g0450(.A1(new_n650), .A2(KEYINPUT27), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(KEYINPUT27), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n651), .A2(G213), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(G343), .ZN(new_n654));
  XNOR2_X1  g0454(.A(new_n654), .B(KEYINPUT90), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n655), .A2(new_n602), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n657), .A2(new_n601), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT91), .ZN(new_n659));
  XNOR2_X1  g0459(.A(new_n605), .B(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n658), .B1(new_n660), .B2(new_n657), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(G330), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n580), .B1(new_n613), .B2(new_n655), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n664), .B1(new_n571), .B2(new_n655), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n655), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n667), .B1(new_n614), .B2(new_n615), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n601), .A2(new_n655), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n668), .B1(new_n580), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n666), .A2(new_n671), .ZN(G399));
  NOR2_X1   g0472(.A1(new_n498), .A2(G116), .ZN(new_n673));
  INV_X1    g0473(.A(new_n207), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n674), .A2(G41), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n673), .A2(G1), .A3(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(new_n228), .B2(new_n676), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n678), .B(KEYINPUT28), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT29), .ZN(new_n680));
  INV_X1    g0480(.A(new_n477), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n681), .A2(new_n523), .A3(new_n629), .A4(new_n532), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n628), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n621), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n620), .B1(new_n523), .B2(new_n532), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n633), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n683), .B1(new_n686), .B2(KEYINPUT26), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT94), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n611), .A2(new_n612), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n569), .B1(new_n689), .B2(new_n538), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n688), .B1(new_n690), .B2(new_n601), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n571), .A2(KEYINPUT94), .A3(new_n616), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n622), .A2(new_n691), .A3(new_n623), .A4(new_n692), .ZN(new_n693));
  AOI211_X1 g0493(.A(new_n680), .B(new_n667), .C1(new_n687), .C2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n636), .A2(new_n655), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n694), .B1(new_n680), .B2(new_n695), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n580), .A2(new_n533), .A3(new_n605), .A4(new_n655), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT93), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT30), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n598), .A2(G179), .A3(new_n520), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n566), .A2(new_n254), .ZN(new_n701));
  INV_X1    g0501(.A(new_n560), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n703), .A2(new_n456), .A3(new_n451), .A4(new_n457), .ZN(new_n704));
  OAI211_X1 g0504(.A(new_n698), .B(new_n699), .C1(new_n700), .C2(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n483), .A2(new_n598), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n706), .A2(new_n271), .A3(new_n519), .A4(new_n567), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n594), .A2(new_n519), .A3(new_n267), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n708), .A2(KEYINPUT30), .A3(new_n483), .A4(new_n703), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n705), .A2(new_n707), .A3(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n708), .A2(new_n483), .A3(new_n703), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n698), .B1(new_n711), .B2(new_n699), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n667), .B1(new_n710), .B2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT31), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XOR2_X1   g0515(.A(KEYINPUT92), .B(KEYINPUT31), .Z(new_n716));
  NAND2_X1  g0516(.A1(new_n707), .A2(new_n709), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n711), .A2(new_n699), .ZN(new_n718));
  OAI211_X1 g0518(.A(new_n667), .B(new_n716), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n697), .A2(new_n715), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(G330), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(KEYINPUT95), .B1(new_n696), .B2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT95), .ZN(new_n724));
  AOI21_X1  g0524(.A(KEYINPUT29), .B1(new_n636), .B2(new_n655), .ZN(new_n725));
  OAI211_X1 g0525(.A(new_n724), .B(new_n721), .C1(new_n725), .C2(new_n694), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n679), .B1(new_n727), .B2(G1), .ZN(G364));
  NOR2_X1   g0528(.A1(G13), .A2(G33), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(G20), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n661), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n225), .A2(G179), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n734), .A2(new_n434), .A3(G200), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n306), .B1(new_n736), .B2(G107), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n271), .A2(new_n225), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n738), .A2(G190), .A3(G200), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(G200), .ZN(new_n740));
  OR3_X1    g0540(.A1(new_n740), .A2(KEYINPUT98), .A3(G190), .ZN(new_n741));
  OAI21_X1  g0541(.A(KEYINPUT98), .B1(new_n740), .B2(G190), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  OAI221_X1 g0544(.A(new_n737), .B1(new_n202), .B2(new_n739), .C1(new_n744), .C2(new_n213), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n734), .A2(G190), .A3(G200), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(new_n497), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n434), .A2(G200), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n738), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(G58), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G190), .A2(G200), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n738), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n749), .A2(new_n267), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G20), .ZN(new_n758));
  AOI22_X1  g0558(.A1(new_n756), .A2(G77), .B1(G97), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n734), .A2(new_n754), .ZN(new_n760));
  INV_X1    g0560(.A(G159), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g0562(.A(KEYINPUT97), .B(KEYINPUT32), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n762), .B(new_n763), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n748), .A2(new_n753), .A3(new_n759), .A4(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(G322), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n750), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(G283), .ZN(new_n768));
  INV_X1    g0568(.A(G326), .ZN(new_n769));
  OAI221_X1 g0569(.A(new_n306), .B1(new_n768), .B2(new_n735), .C1(new_n739), .C2(new_n769), .ZN(new_n770));
  AOI211_X1 g0570(.A(new_n767), .B(new_n770), .C1(G311), .C2(new_n756), .ZN(new_n771));
  INV_X1    g0571(.A(new_n760), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G329), .ZN(new_n773));
  XNOR2_X1  g0573(.A(KEYINPUT33), .B(G317), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n743), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n746), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(G303), .ZN(new_n777));
  NAND4_X1  g0577(.A1(new_n771), .A2(new_n773), .A3(new_n775), .A4(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n758), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n561), .ZN(new_n780));
  OR2_X1    g0580(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n765), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(KEYINPUT99), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n224), .B1(G20), .B2(new_n273), .ZN(new_n784));
  INV_X1    g0584(.A(KEYINPUT99), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n765), .A2(new_n781), .A3(new_n785), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n783), .A2(new_n784), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n649), .A2(G45), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n676), .A2(G1), .A3(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n311), .A2(new_n312), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n674), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n229), .A2(new_n510), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n793), .B(new_n794), .C1(new_n510), .C2(new_n245), .ZN(new_n795));
  INV_X1    g0595(.A(G355), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n247), .A2(new_n207), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n795), .B1(G116), .B2(new_n207), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n731), .A2(new_n784), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n787), .A2(new_n790), .A3(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n733), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(KEYINPUT96), .B1(new_n661), .B2(G330), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n661), .A2(KEYINPUT96), .A3(G330), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n661), .ZN(new_n807));
  INV_X1    g0607(.A(G330), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n790), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n802), .B1(new_n806), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n810), .A2(KEYINPUT100), .ZN(new_n811));
  INV_X1    g0611(.A(KEYINPUT100), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n812), .B(new_n802), .C1(new_n806), .C2(new_n809), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(G396));
  INV_X1    g0615(.A(KEYINPUT102), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n294), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g0617(.A1(new_n272), .A2(new_n274), .A3(KEYINPUT102), .A4(new_n293), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n415), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n667), .A2(new_n293), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n819), .A2(new_n820), .B1(new_n640), .B2(new_n667), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n695), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n636), .A2(new_n655), .A3(new_n819), .ZN(new_n823));
  AND2_X1   g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  OR2_X1    g0624(.A1(new_n824), .A2(new_n722), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(new_n722), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n825), .A2(new_n826), .A3(new_n789), .ZN(new_n827));
  INV_X1    g0627(.A(new_n739), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n743), .A2(G150), .B1(G137), .B2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(G143), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n829), .B1(new_n830), .B2(new_n750), .C1(new_n761), .C2(new_n755), .ZN(new_n831));
  XOR2_X1   g0631(.A(new_n831), .B(KEYINPUT101), .Z(new_n832));
  XNOR2_X1  g0632(.A(new_n832), .B(KEYINPUT34), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n779), .A2(new_n751), .B1(new_n746), .B2(new_n202), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n791), .B1(G132), .B2(new_n772), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n213), .B2(new_n735), .ZN(new_n836));
  NOR3_X1   g0636(.A1(new_n833), .A2(new_n834), .A3(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n750), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n838), .A2(G294), .B1(G311), .B2(new_n772), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n839), .B1(new_n581), .B2(new_n755), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n743), .A2(G283), .B1(G107), .B2(new_n776), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n247), .B1(new_n758), .B2(G97), .ZN(new_n842));
  INV_X1    g0642(.A(G303), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n841), .B(new_n842), .C1(new_n843), .C2(new_n739), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n840), .B(new_n844), .C1(G87), .C2(new_n736), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n784), .B1(new_n837), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n821), .A2(new_n729), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n784), .A2(new_n729), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(new_n277), .ZN(new_n849));
  NAND4_X1  g0649(.A1(new_n846), .A2(new_n790), .A3(new_n847), .A4(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n827), .A2(new_n850), .ZN(G384));
  XOR2_X1   g0651(.A(KEYINPUT106), .B(KEYINPUT40), .Z(new_n852));
  NAND2_X1  g0652(.A1(new_n343), .A2(new_n281), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n314), .A2(G68), .ZN(new_n854));
  AOI21_X1  g0654(.A(KEYINPUT16), .B1(new_n854), .B2(new_n301), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n298), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(KEYINPUT103), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT103), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n858), .B(new_n298), .C1(new_n853), .C2(new_n855), .ZN(new_n859));
  INV_X1    g0659(.A(new_n653), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n349), .A2(new_n351), .A3(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n857), .A2(new_n859), .A3(new_n861), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n862), .A2(new_n345), .ZN(new_n863));
  AND3_X1   g0663(.A1(new_n857), .A2(new_n653), .A3(new_n859), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n863), .A2(KEYINPUT37), .B1(new_n355), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n348), .B1(new_n352), .B2(new_n653), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n345), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT37), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(KEYINPUT38), .B1(new_n865), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n355), .A2(new_n864), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n862), .A2(KEYINPUT37), .A3(new_n345), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n871), .A2(KEYINPUT38), .A3(new_n869), .A4(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n870), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n716), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n713), .A2(new_n876), .ZN(new_n877));
  OAI211_X1 g0677(.A(KEYINPUT31), .B(new_n667), .C1(new_n710), .C2(new_n712), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n697), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n821), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n367), .A2(new_n667), .ZN(new_n881));
  AND3_X1   g0681(.A1(new_n417), .A2(new_n418), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n881), .B1(new_n417), .B2(new_n418), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n879), .B(new_n880), .C1(new_n882), .C2(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n852), .B1(new_n875), .B2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT40), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT38), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n860), .B1(new_n344), .B2(new_n298), .ZN(new_n888));
  AND2_X1   g0688(.A1(new_n355), .A2(new_n888), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n344), .A2(new_n298), .B1(new_n349), .B2(new_n351), .ZN(new_n890));
  NOR3_X1   g0690(.A1(new_n890), .A2(new_n888), .A3(KEYINPUT104), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n867), .B1(new_n891), .B2(new_n868), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n866), .A2(KEYINPUT104), .A3(KEYINPUT37), .A4(new_n345), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n887), .B1(new_n889), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n886), .B1(new_n895), .B2(new_n873), .ZN(new_n896));
  INV_X1    g0696(.A(new_n881), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n419), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n410), .A2(new_n881), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n821), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n896), .A2(new_n879), .A3(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n885), .A2(G330), .A3(new_n901), .ZN(new_n902));
  NOR3_X1   g0702(.A1(new_n412), .A2(new_n420), .A3(new_n442), .ZN(new_n903));
  INV_X1    g0703(.A(new_n441), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n903), .A2(G330), .A3(new_n904), .A4(new_n879), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n871), .A2(new_n869), .A3(new_n872), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n887), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n873), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n909), .A2(new_n900), .A3(new_n879), .ZN(new_n910));
  INV_X1    g0710(.A(new_n884), .ZN(new_n911));
  AOI22_X1  g0711(.A1(new_n910), .A2(new_n852), .B1(new_n911), .B2(new_n896), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n912), .A2(new_n443), .A3(new_n879), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n906), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT39), .ZN(new_n915));
  AND3_X1   g0715(.A1(new_n895), .A2(new_n915), .A3(new_n873), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n915), .B1(new_n908), .B2(new_n873), .ZN(new_n917));
  OAI21_X1  g0717(.A(KEYINPUT105), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(KEYINPUT39), .B1(new_n870), .B2(new_n874), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT105), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n895), .A2(new_n915), .A3(new_n873), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n417), .A2(new_n667), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n918), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n882), .A2(new_n883), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n817), .A2(new_n655), .A3(new_n818), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n925), .B1(new_n823), .B2(new_n926), .ZN(new_n927));
  AOI22_X1  g0727(.A1(new_n927), .A2(new_n909), .B1(new_n639), .B2(new_n860), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n924), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n914), .B(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n646), .B1(new_n696), .B2(new_n443), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n930), .B(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n257), .B2(new_n649), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n467), .A2(new_n471), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n581), .B1(new_n934), .B2(KEYINPUT35), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n935), .B(new_n226), .C1(KEYINPUT35), .C2(new_n934), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(KEYINPUT36), .ZN(new_n937));
  OAI21_X1  g0737(.A(G77), .B1(new_n751), .B2(new_n213), .ZN(new_n938));
  OAI22_X1  g0738(.A1(new_n228), .A2(new_n938), .B1(G50), .B2(new_n213), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n939), .A2(G1), .A3(new_n275), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n933), .A2(new_n937), .A3(new_n940), .ZN(G367));
  NAND2_X1  g0741(.A1(new_n580), .A2(new_n670), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n485), .B(new_n477), .C1(new_n482), .C2(new_n655), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT42), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n477), .B1(new_n943), .B2(new_n571), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n655), .ZN(new_n947));
  INV_X1    g0747(.A(new_n622), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n655), .B1(new_n524), .B2(new_n526), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n626), .A2(new_n627), .A3(new_n949), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AOI22_X1  g0752(.A1(new_n945), .A2(new_n947), .B1(KEYINPUT43), .B2(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n952), .A2(KEYINPUT43), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n953), .B(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n666), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n681), .A2(new_n667), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n943), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n955), .B(new_n959), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n675), .B(KEYINPUT41), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n942), .B1(new_n665), .B2(new_n670), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n662), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(new_n806), .B2(new_n963), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT45), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT107), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n671), .A2(new_n967), .A3(new_n958), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n967), .B1(new_n671), .B2(new_n958), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n966), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n970), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n972), .A2(KEYINPUT45), .A3(new_n968), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT44), .ZN(new_n974));
  OR3_X1    g0774(.A1(new_n671), .A2(new_n974), .A3(new_n958), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n974), .B1(new_n671), .B2(new_n958), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n971), .A2(new_n973), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n956), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n666), .A2(new_n977), .A3(new_n973), .A4(new_n971), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n727), .A2(new_n965), .A3(new_n979), .A4(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n962), .B1(new_n981), .B2(new_n727), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n788), .A2(G1), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n960), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(G317), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n760), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(G311), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n739), .A2(new_n987), .B1(new_n496), .B2(new_n735), .ZN(new_n988));
  AOI211_X1 g0788(.A(new_n986), .B(new_n988), .C1(new_n743), .C2(G294), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n791), .B1(new_n779), .B2(new_n219), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n746), .A2(new_n581), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT46), .ZN(new_n992));
  AOI211_X1 g0792(.A(new_n990), .B(new_n992), .C1(G283), .C2(new_n756), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n989), .B(new_n993), .C1(new_n843), .C2(new_n750), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT108), .Z(new_n995));
  INV_X1    g0795(.A(G150), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n750), .A2(new_n996), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n744), .A2(new_n761), .B1(new_n202), .B2(new_n755), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n306), .B1(new_n736), .B2(G77), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n998), .B1(KEYINPUT109), .B2(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(KEYINPUT109), .B2(new_n999), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n997), .B(new_n1001), .C1(G143), .C2(new_n828), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n772), .A2(G137), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n1002), .B(new_n1003), .C1(new_n751), .C2(new_n746), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n779), .A2(new_n213), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n995), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT47), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n784), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n950), .A2(new_n731), .A3(new_n951), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n793), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n799), .B1(new_n207), .B2(new_n507), .C1(new_n1010), .C2(new_n238), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n1008), .A2(new_n790), .A3(new_n1009), .A4(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n984), .A2(new_n1012), .ZN(G387));
  AND2_X1   g0813(.A1(new_n806), .A2(new_n963), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n726), .B(new_n723), .C1(new_n1014), .C2(new_n964), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n727), .A2(new_n965), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1015), .A2(new_n675), .A3(new_n1016), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n791), .B1(new_n581), .B2(new_n735), .C1(new_n769), .C2(new_n760), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT113), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n743), .A2(G311), .B1(G322), .B2(new_n828), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT112), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(G303), .A2(new_n756), .B1(new_n838), .B2(G317), .ZN(new_n1022));
  AND2_X1   g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT48), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  AND3_X1   g0825(.A1(new_n1021), .A2(new_n1024), .A3(new_n1022), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT49), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n758), .A2(G283), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n776), .A2(G294), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1029), .B(new_n1030), .C1(new_n1025), .C2(new_n1026), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(KEYINPUT49), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1019), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n743), .A2(new_n421), .B1(G97), .B2(new_n736), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT111), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n776), .A2(G77), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n996), .B2(new_n760), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1035), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n739), .A2(new_n761), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n779), .A2(new_n507), .ZN(new_n1041));
  AND2_X1   g0841(.A1(new_n1038), .A2(new_n1036), .ZN(new_n1042));
  NOR4_X1   g0842(.A1(new_n1039), .A2(new_n1040), .A3(new_n1041), .A4(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n756), .A2(G68), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1043), .A2(new_n792), .A3(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(G50), .B2(new_n838), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n784), .B1(new_n1034), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n235), .A2(G45), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n673), .B(new_n510), .C1(new_n213), .C2(new_n277), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT110), .Z(new_n1050));
  NOR2_X1   g0850(.A1(new_n285), .A2(G50), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(KEYINPUT50), .Z(new_n1052));
  OAI211_X1 g0852(.A(new_n793), .B(new_n1048), .C1(new_n1050), .C2(new_n1052), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1053), .B1(G107), .B2(new_n207), .C1(new_n673), .C2(new_n797), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n789), .B1(new_n1054), .B2(new_n799), .ZN(new_n1055));
  AND2_X1   g0855(.A1(new_n1047), .A2(new_n1055), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n665), .A2(new_n732), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n1056), .A2(new_n1057), .B1(new_n965), .B2(new_n983), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1017), .A2(new_n1058), .ZN(G393));
  NAND3_X1  g0859(.A1(new_n979), .A2(new_n980), .A3(KEYINPUT114), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT114), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n978), .A2(new_n1061), .A3(new_n956), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1016), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n675), .B(new_n981), .C1(new_n1063), .C2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1063), .A2(new_n983), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n739), .A2(new_n996), .B1(new_n750), .B2(new_n761), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1067), .B(KEYINPUT51), .Z(new_n1068));
  OAI21_X1  g0868(.A(new_n792), .B1(new_n755), .B2(new_n285), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n779), .A2(new_n277), .ZN(new_n1070));
  NOR3_X1   g0870(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n743), .A2(G50), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n776), .A2(G68), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n735), .A2(new_n497), .B1(new_n760), .B2(new_n830), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .A4(new_n1075), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n743), .A2(G303), .B1(G116), .B2(new_n758), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT115), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n739), .A2(new_n985), .B1(new_n750), .B2(new_n987), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT52), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n306), .B1(new_n760), .B2(new_n766), .C1(new_n768), .C2(new_n746), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(G107), .B2(new_n736), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1078), .A2(new_n1080), .A3(new_n1082), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n755), .A2(new_n561), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1076), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n784), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n799), .B1(new_n207), .B2(new_n496), .C1(new_n1010), .C2(new_n242), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n943), .A2(new_n731), .A3(new_n957), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1086), .A2(new_n790), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(KEYINPUT116), .B1(new_n1066), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n983), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1091), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT116), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1089), .ZN(new_n1094));
  NOR3_X1   g0894(.A1(new_n1092), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1065), .B1(new_n1090), .B2(new_n1095), .ZN(G390));
  NOR2_X1   g0896(.A1(new_n821), .A2(new_n808), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n879), .B(new_n1097), .C1(new_n882), .C2(new_n883), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  AND4_X1   g0899(.A1(new_n622), .A2(new_n691), .A3(new_n623), .A4(new_n692), .ZN(new_n1100));
  AND2_X1   g0900(.A1(new_n628), .A2(new_n682), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n630), .A2(new_n632), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(new_n619), .B2(new_n621), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1101), .B1(new_n1103), .B2(new_n629), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n655), .B(new_n819), .C1(new_n1100), .C2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n925), .B1(new_n1105), .B2(new_n926), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n895), .A2(new_n873), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n923), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(KEYINPUT117), .B1(new_n1106), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT117), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n923), .B1(new_n895), .B2(new_n873), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n926), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n667), .B1(new_n687), .B2(new_n693), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1113), .B1(new_n1114), .B2(new_n819), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1111), .B(new_n1112), .C1(new_n1115), .C2(new_n925), .ZN(new_n1116));
  AND2_X1   g0916(.A1(new_n1110), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n823), .A2(new_n926), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n898), .A2(new_n899), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n918), .A2(new_n922), .B1(new_n1120), .B2(new_n1108), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1099), .B1(new_n1117), .B2(new_n1121), .ZN(new_n1122));
  NOR3_X1   g0922(.A1(new_n916), .A2(new_n917), .A3(KEYINPUT105), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n920), .B1(new_n919), .B2(new_n921), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n1123), .A2(new_n1124), .B1(new_n923), .B2(new_n927), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1110), .A2(new_n1116), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n722), .A2(new_n900), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1122), .A2(new_n983), .A3(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n729), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n848), .A2(new_n285), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n247), .B(new_n1070), .C1(new_n838), .C2(G116), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n743), .A2(G107), .B1(new_n466), .B2(new_n756), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1132), .B1(new_n1133), .B2(KEYINPUT118), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n1133), .A2(KEYINPUT118), .B1(G68), .B2(new_n736), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n1135), .B1(new_n497), .B2(new_n746), .C1(new_n768), .C2(new_n739), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n1134), .B(new_n1136), .C1(G294), .C2(new_n772), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n772), .A2(G125), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1138), .B1(new_n779), .B2(new_n761), .ZN(new_n1139));
  XOR2_X1   g0939(.A(KEYINPUT54), .B(G143), .Z(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n776), .A2(G150), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n755), .A2(new_n1141), .B1(new_n1142), .B2(KEYINPUT53), .ZN(new_n1143));
  AOI211_X1 g0943(.A(new_n1139), .B(new_n1143), .C1(G132), .C2(new_n838), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n306), .B1(new_n743), .B2(G137), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n1142), .A2(KEYINPUT53), .B1(G50), .B2(new_n736), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1144), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(G128), .B2(new_n828), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1137), .A2(new_n1148), .ZN(new_n1149));
  XOR2_X1   g0949(.A(new_n1149), .B(KEYINPUT119), .Z(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n784), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1130), .A2(new_n790), .A3(new_n1131), .A4(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1129), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n696), .A2(new_n443), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1154), .A2(new_n647), .A3(new_n905), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n879), .A2(new_n1097), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n722), .A2(new_n900), .B1(new_n1156), .B2(new_n925), .ZN(new_n1157));
  AND2_X1   g0957(.A1(new_n720), .A2(new_n1097), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1098), .B1(new_n1158), .B2(new_n1119), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n1157), .A2(new_n1115), .B1(new_n1159), .B2(new_n1118), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1155), .A2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1122), .A2(new_n1128), .A3(new_n1161), .ZN(new_n1162));
  AND2_X1   g0962(.A1(new_n1162), .A2(new_n675), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1159), .A2(new_n1118), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1156), .A2(new_n925), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1127), .A2(new_n1115), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1167), .A2(new_n931), .A3(new_n905), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1128), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1098), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1168), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1153), .B1(new_n1163), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(G378));
  NAND2_X1  g0973(.A1(new_n848), .A2(new_n202), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n427), .A2(new_n653), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n436), .A2(new_n440), .A3(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1177), .B1(new_n436), .B2(new_n440), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1176), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1177), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n441), .A2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1183), .A2(new_n1178), .A3(new_n1175), .ZN(new_n1184));
  AND2_X1   g0984(.A1(new_n1181), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1174), .B1(new_n1186), .B2(new_n730), .ZN(new_n1187));
  INV_X1    g0987(.A(G124), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n252), .B1(new_n760), .B2(new_n1188), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1141), .A2(new_n746), .ZN(new_n1190));
  INV_X1    g0990(.A(G128), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n1190), .A2(KEYINPUT120), .B1(new_n750), .B2(new_n1191), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n828), .A2(G125), .B1(new_n756), .B2(G137), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1193), .B1(new_n996), .B2(new_n779), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n1192), .B(new_n1194), .C1(KEYINPUT120), .C2(new_n1190), .ZN(new_n1195));
  INV_X1    g0995(.A(G132), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1195), .B1(new_n1196), .B2(new_n744), .ZN(new_n1197));
  AOI211_X1 g0997(.A(G41), .B(new_n1189), .C1(new_n1197), .C2(KEYINPUT59), .ZN(new_n1198));
  OAI221_X1 g0998(.A(new_n1198), .B1(KEYINPUT59), .B2(new_n1197), .C1(new_n761), .C2(new_n735), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1005), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n253), .B(new_n791), .C1(new_n739), .C2(new_n581), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(new_n743), .B2(G97), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n735), .A2(new_n751), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1202), .B(new_n1204), .C1(new_n507), .C2(new_n755), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(G107), .B2(new_n838), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n772), .A2(G283), .ZN(new_n1207));
  AND4_X1   g1007(.A1(new_n1200), .A2(new_n1206), .A3(new_n1037), .A4(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(KEYINPUT58), .ZN(new_n1209));
  OR2_X1    g1009(.A1(new_n1208), .A2(KEYINPUT58), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n253), .B1(new_n791), .B2(new_n252), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(new_n202), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1199), .A2(new_n1209), .A3(new_n1210), .A4(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1187), .B1(new_n784), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(new_n790), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1185), .B1(new_n912), .B2(G330), .ZN(new_n1216));
  AND4_X1   g1016(.A1(G330), .A2(new_n885), .A3(new_n901), .A4(new_n1185), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n929), .A2(KEYINPUT121), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  OAI211_X1 g1020(.A(KEYINPUT121), .B(new_n929), .C1(new_n1216), .C2(new_n1217), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1215), .B1(new_n1222), .B2(new_n1091), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1155), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1162), .A2(new_n1225), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n929), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n902), .A2(new_n1186), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n885), .A2(new_n1185), .A3(G330), .A4(new_n901), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1228), .A2(new_n924), .A3(new_n928), .A4(new_n1229), .ZN(new_n1230));
  AND3_X1   g1030(.A1(new_n1227), .A2(KEYINPUT57), .A3(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1226), .A2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(new_n675), .ZN(new_n1233));
  AND2_X1   g1033(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1234));
  AOI21_X1  g1034(.A(KEYINPUT57), .B1(new_n1234), .B2(new_n1226), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1224), .B1(new_n1233), .B2(new_n1235), .ZN(G375));
  NAND2_X1  g1036(.A1(new_n1155), .A2(new_n1160), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1237), .A2(new_n1168), .A3(new_n961), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n925), .A2(new_n729), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n743), .A2(G116), .B1(G303), .B2(new_n772), .ZN(new_n1240));
  OAI221_X1 g1040(.A(new_n1240), .B1(new_n376), .B2(new_n746), .C1(new_n768), .C2(new_n750), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n739), .A2(new_n561), .ZN(new_n1242));
  OAI221_X1 g1042(.A(new_n306), .B1(new_n277), .B2(new_n735), .C1(new_n755), .C2(new_n219), .ZN(new_n1243));
  NOR4_X1   g1043(.A1(new_n1241), .A2(new_n1041), .A3(new_n1242), .A4(new_n1243), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n743), .A2(new_n1140), .B1(G128), .B2(new_n772), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n756), .A2(G150), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n838), .A2(G137), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1245), .A2(new_n1204), .A3(new_n1246), .A4(new_n1247), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n779), .A2(new_n202), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n739), .A2(new_n1196), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n792), .B1(new_n761), .B2(new_n746), .ZN(new_n1251));
  NOR4_X1   g1051(.A1(new_n1248), .A2(new_n1249), .A3(new_n1250), .A4(new_n1251), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n784), .B1(new_n1244), .B2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n848), .A2(new_n213), .ZN(new_n1254));
  AND4_X1   g1054(.A1(new_n790), .A2(new_n1239), .A3(new_n1253), .A4(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1255), .B1(new_n1167), .B2(new_n983), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1238), .A2(new_n1256), .ZN(G381));
  INV_X1    g1057(.A(KEYINPUT57), .ZN(new_n1258));
  AND2_X1   g1058(.A1(new_n1162), .A2(new_n1225), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1258), .B1(new_n1259), .B2(new_n1222), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n676), .B1(new_n1226), .B2(new_n1231), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1223), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n1172), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1066), .A2(KEYINPUT116), .A3(new_n1089), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1093), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1266), .A2(new_n984), .A3(new_n1012), .A4(new_n1065), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n675), .B1(new_n727), .B2(new_n965), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n814), .B(new_n1058), .C1(new_n1064), .C2(new_n1268), .ZN(new_n1269));
  NOR4_X1   g1069(.A1(new_n1267), .A2(G384), .A3(G381), .A4(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT122), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1263), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1272), .B1(new_n1271), .B2(new_n1270), .ZN(G407));
  OAI211_X1 g1073(.A(G407), .B(G213), .C1(G343), .C2(new_n1263), .ZN(G409));
  INV_X1    g1074(.A(G213), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1275), .A2(G343), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1234), .A2(new_n1226), .A3(new_n961), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1227), .A2(new_n1230), .A3(new_n983), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1172), .A2(new_n1215), .A3(new_n1278), .A4(new_n1279), .ZN(new_n1280));
  OAI211_X1 g1080(.A(new_n1277), .B(new_n1280), .C1(new_n1262), .C2(new_n1172), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1155), .A2(KEYINPUT60), .A3(new_n1160), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1282), .A2(new_n1168), .A3(new_n675), .ZN(new_n1283));
  AOI21_X1  g1083(.A(KEYINPUT60), .B1(new_n1155), .B2(new_n1160), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1256), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(G384), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  OAI211_X1 g1087(.A(G384), .B(new_n1256), .C1(new_n1283), .C2(new_n1284), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  OAI21_X1  g1089(.A(KEYINPUT62), .B1(new_n1281), .B2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT61), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1276), .A2(G2897), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1293), .B1(new_n1289), .B2(KEYINPUT123), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT123), .ZN(new_n1295));
  AOI211_X1 g1095(.A(new_n1295), .B(new_n1292), .C1(new_n1287), .C2(new_n1288), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1294), .A2(new_n1296), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1289), .A2(KEYINPUT123), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1172), .B1(new_n1300), .B2(new_n1224), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1171), .A2(new_n675), .A3(new_n1162), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1153), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1303), .A2(new_n1304), .A3(new_n1215), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1277), .B1(new_n1302), .B2(new_n1305), .ZN(new_n1306));
  OAI211_X1 g1106(.A(new_n1297), .B(new_n1299), .C1(new_n1301), .C2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(G375), .A2(G378), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1279), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1222), .B1(new_n1225), .B2(new_n1162), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1309), .B1(new_n1310), .B2(new_n961), .ZN(new_n1311));
  AND3_X1   g1111(.A1(new_n1303), .A2(new_n1304), .A3(new_n1215), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1276), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT62), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1289), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1308), .A2(new_n1313), .A3(new_n1314), .A4(new_n1315), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1290), .A2(new_n1291), .A3(new_n1307), .A4(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT126), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n814), .B1(new_n1017), .B2(new_n1058), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1320), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1321), .A2(KEYINPUT124), .A3(new_n1269), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT124), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1269), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1323), .B1(new_n1324), .B2(new_n1320), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1322), .A2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(G390), .A2(G387), .ZN(new_n1327));
  AND3_X1   g1127(.A1(new_n1326), .A2(new_n1327), .A3(new_n1267), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1322), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1329), .B1(new_n1327), .B2(new_n1267), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1328), .A2(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT127), .ZN(new_n1332));
  XNOR2_X1  g1132(.A(new_n1331), .B(new_n1332), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1298), .B1(new_n1308), .B2(new_n1313), .ZN(new_n1334));
  AOI21_X1  g1134(.A(KEYINPUT61), .B1(new_n1334), .B2(new_n1297), .ZN(new_n1335));
  NAND4_X1  g1135(.A1(new_n1335), .A2(KEYINPUT126), .A3(new_n1316), .A4(new_n1290), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1319), .A2(new_n1333), .A3(new_n1336), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1291), .B1(new_n1328), .B2(new_n1330), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT125), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1338), .A2(new_n1339), .ZN(new_n1340));
  OAI211_X1 g1140(.A(KEYINPUT125), .B(new_n1291), .C1(new_n1328), .C2(new_n1330), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1340), .A2(new_n1341), .ZN(new_n1342));
  NOR2_X1   g1142(.A1(new_n1281), .A2(new_n1289), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1343), .A2(KEYINPUT63), .ZN(new_n1344));
  AND2_X1   g1144(.A1(new_n1307), .A2(KEYINPUT63), .ZN(new_n1345));
  OAI211_X1 g1145(.A(new_n1342), .B(new_n1344), .C1(new_n1343), .C2(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1337), .A2(new_n1346), .ZN(G405));
  NAND2_X1  g1147(.A1(new_n1263), .A2(new_n1308), .ZN(new_n1348));
  XNOR2_X1  g1148(.A(new_n1348), .B(new_n1289), .ZN(new_n1349));
  XNOR2_X1  g1149(.A(new_n1349), .B(new_n1331), .ZN(G402));
endmodule


