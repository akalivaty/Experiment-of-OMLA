

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783;

  OR2_X1 U376 ( .A1(n579), .A2(n578), .ZN(n581) );
  XNOR2_X1 U377 ( .A(n464), .B(G469), .ZN(n602) );
  NAND2_X2 U378 ( .A1(n387), .A2(n390), .ZN(n726) );
  XNOR2_X1 U379 ( .A(n497), .B(n452), .ZN(n517) );
  XNOR2_X1 U380 ( .A(n469), .B(n456), .ZN(n771) );
  XNOR2_X1 U381 ( .A(n552), .B(KEYINPUT97), .ZN(n728) );
  INV_X1 U382 ( .A(G953), .ZN(n509) );
  BUF_X1 U383 ( .A(n715), .Z(n355) );
  XNOR2_X1 U384 ( .A(n563), .B(KEYINPUT35), .ZN(n593) );
  XNOR2_X1 U385 ( .A(n574), .B(KEYINPUT106), .ZN(n781) );
  XNOR2_X1 U386 ( .A(n602), .B(n540), .ZN(n715) );
  NOR2_X2 U387 ( .A1(n610), .A2(n550), .ZN(n551) );
  INV_X1 U388 ( .A(G146), .ZN(n417) );
  INV_X1 U389 ( .A(KEYINPUT88), .ZN(n435) );
  XNOR2_X1 U390 ( .A(n642), .B(n641), .ZN(n372) );
  AND2_X1 U391 ( .A1(n781), .A2(n584), .ZN(n596) );
  XNOR2_X1 U392 ( .A(n436), .B(n435), .ZN(n573) );
  NOR2_X1 U393 ( .A1(n633), .A2(n637), .ZN(n539) );
  XNOR2_X1 U394 ( .A(n451), .B(KEYINPUT69), .ZN(n716) );
  AND2_X1 U395 ( .A1(n377), .A2(n389), .ZN(n387) );
  XNOR2_X1 U396 ( .A(n471), .B(n470), .ZN(n655) );
  XNOR2_X1 U397 ( .A(n415), .B(n412), .ZN(n687) );
  XNOR2_X1 U398 ( .A(n517), .B(n454), .ZN(n469) );
  INV_X1 U399 ( .A(n505), .ZN(n506) );
  XNOR2_X1 U400 ( .A(n417), .B(G125), .ZN(n519) );
  INV_X2 U401 ( .A(G107), .ZN(n367) );
  XNOR2_X1 U402 ( .A(G137), .B(G113), .ZN(n465) );
  XNOR2_X1 U403 ( .A(KEYINPUT72), .B(G110), .ZN(n518) );
  OR2_X2 U404 ( .A1(n591), .A2(n586), .ZN(n587) );
  AND2_X2 U405 ( .A1(n570), .A2(n569), .ZN(n572) );
  AND2_X2 U406 ( .A1(n716), .A2(n715), .ZN(n559) );
  OR2_X2 U407 ( .A1(n591), .A2(n437), .ZN(n436) );
  XNOR2_X2 U408 ( .A(n572), .B(n571), .ZN(n591) );
  OR2_X1 U409 ( .A1(n390), .A2(n360), .ZN(n385) );
  NOR2_X1 U410 ( .A1(n382), .A2(n381), .ZN(n380) );
  NOR2_X1 U411 ( .A1(n387), .A2(n360), .ZN(n381) );
  NAND2_X1 U412 ( .A1(n385), .A2(n383), .ZN(n382) );
  NAND2_X1 U413 ( .A1(n384), .A2(n473), .ZN(n383) );
  NAND2_X1 U414 ( .A1(n379), .A2(n387), .ZN(n378) );
  XNOR2_X1 U415 ( .A(KEYINPUT3), .B(G119), .ZN(n467) );
  XOR2_X1 U416 ( .A(G116), .B(G101), .Z(n468) );
  XNOR2_X1 U417 ( .A(n442), .B(n430), .ZN(n493) );
  INV_X1 U418 ( .A(KEYINPUT8), .ZN(n430) );
  XNOR2_X1 U419 ( .A(n515), .B(n516), .ZN(n434) );
  INV_X1 U420 ( .A(KEYINPUT77), .ZN(n516) );
  NOR2_X1 U421 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U422 ( .A(n502), .B(n501), .ZN(n566) );
  OR2_X1 U423 ( .A1(n662), .A2(G902), .ZN(n464) );
  XNOR2_X1 U424 ( .A(G140), .B(G137), .ZN(n455) );
  XNOR2_X1 U425 ( .A(n357), .B(n441), .ZN(n414) );
  XNOR2_X1 U426 ( .A(G119), .B(G128), .ZN(n441) );
  XNOR2_X1 U427 ( .A(n519), .B(n416), .ZN(n769) );
  XNOR2_X1 U428 ( .A(KEYINPUT10), .B(KEYINPUT70), .ZN(n416) );
  INV_X1 U429 ( .A(n777), .ZN(n706) );
  NAND2_X1 U430 ( .A1(n372), .A2(n643), .ZN(n777) );
  NAND2_X1 U431 ( .A1(n396), .A2(n395), .ZN(n393) );
  XNOR2_X1 U432 ( .A(n448), .B(n447), .ZN(n588) );
  XNOR2_X1 U433 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U434 ( .A(n491), .B(n411), .ZN(n567) );
  XNOR2_X1 U435 ( .A(n490), .B(n492), .ZN(n411) );
  NOR2_X1 U436 ( .A1(n756), .A2(G953), .ZN(n420) );
  AND2_X1 U437 ( .A1(n400), .A2(n403), .ZN(n402) );
  INV_X1 U438 ( .A(n473), .ZN(n386) );
  INV_X1 U439 ( .A(n734), .ZN(n384) );
  AND2_X1 U440 ( .A1(n509), .A2(n376), .ZN(n486) );
  INV_X1 U441 ( .A(G237), .ZN(n376) );
  INV_X1 U442 ( .A(KEYINPUT17), .ZN(n511) );
  XNOR2_X1 U443 ( .A(n612), .B(KEYINPUT81), .ZN(n621) );
  NAND2_X1 U444 ( .A1(G234), .A2(G237), .ZN(n474) );
  XNOR2_X1 U445 ( .A(n374), .B(n373), .ZN(n466) );
  XNOR2_X1 U446 ( .A(G146), .B(KEYINPUT96), .ZN(n373) );
  XNOR2_X1 U447 ( .A(n375), .B(KEYINPUT5), .ZN(n374) );
  NAND2_X1 U448 ( .A1(n486), .A2(G210), .ZN(n375) );
  XOR2_X1 U449 ( .A(KEYINPUT75), .B(KEYINPUT16), .Z(n504) );
  XOR2_X1 U450 ( .A(G113), .B(G104), .Z(n505) );
  XNOR2_X1 U451 ( .A(G131), .B(KEYINPUT11), .ZN(n484) );
  XNOR2_X1 U452 ( .A(G143), .B(G122), .ZN(n483) );
  XNOR2_X1 U453 ( .A(n505), .B(n485), .ZN(n406) );
  XOR2_X1 U454 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n485) );
  OR2_X1 U455 ( .A1(n588), .A2(n568), .ZN(n451) );
  OR2_X1 U456 ( .A1(n655), .A2(n391), .ZN(n390) );
  NAND2_X1 U457 ( .A1(n472), .A2(G902), .ZN(n389) );
  NAND2_X1 U458 ( .A1(n493), .A2(G217), .ZN(n429) );
  XNOR2_X1 U459 ( .A(n494), .B(KEYINPUT7), .ZN(n428) );
  XNOR2_X1 U460 ( .A(n407), .B(n405), .ZN(n677) );
  XNOR2_X1 U461 ( .A(n769), .B(n408), .ZN(n407) );
  XNOR2_X1 U462 ( .A(n489), .B(n406), .ZN(n405) );
  XNOR2_X1 U463 ( .A(n483), .B(n484), .ZN(n408) );
  XNOR2_X1 U464 ( .A(G101), .B(G146), .ZN(n459) );
  XNOR2_X1 U465 ( .A(G107), .B(G104), .ZN(n460) );
  XNOR2_X1 U466 ( .A(n433), .B(n432), .ZN(n521) );
  XNOR2_X1 U467 ( .A(n517), .B(n514), .ZN(n432) );
  XNOR2_X1 U468 ( .A(n520), .B(n434), .ZN(n433) );
  XNOR2_X1 U469 ( .A(n423), .B(n422), .ZN(n752) );
  INV_X1 U470 ( .A(KEYINPUT41), .ZN(n422) );
  NOR2_X1 U471 ( .A1(n738), .A2(n737), .ZN(n423) );
  NAND2_X1 U472 ( .A1(n392), .A2(n427), .ZN(n633) );
  NOR2_X1 U473 ( .A1(n538), .A2(n600), .ZN(n427) );
  INV_X1 U474 ( .A(KEYINPUT34), .ZN(n371) );
  XNOR2_X1 U475 ( .A(n545), .B(n544), .ZN(n610) );
  XNOR2_X1 U476 ( .A(n425), .B(KEYINPUT28), .ZN(n424) );
  NOR2_X1 U477 ( .A1(n600), .A2(n601), .ZN(n425) );
  OR2_X1 U478 ( .A1(n585), .A2(n355), .ZN(n437) );
  XNOR2_X1 U479 ( .A(n414), .B(n413), .ZN(n412) );
  XNOR2_X1 U480 ( .A(n443), .B(n769), .ZN(n415) );
  XNOR2_X1 U481 ( .A(n455), .B(KEYINPUT24), .ZN(n413) );
  AND2_X1 U482 ( .A1(n398), .A2(n397), .ZN(n394) );
  XNOR2_X1 U483 ( .A(n399), .B(KEYINPUT40), .ZN(n606) );
  XNOR2_X1 U484 ( .A(n410), .B(n409), .ZN(n702) );
  INV_X1 U485 ( .A(KEYINPUT104), .ZN(n409) );
  NOR2_X1 U486 ( .A1(n567), .A2(n536), .ZN(n410) );
  INV_X1 U487 ( .A(KEYINPUT53), .ZN(n418) );
  NAND2_X1 U488 ( .A1(n421), .A2(n420), .ZN(n419) );
  NAND2_X1 U489 ( .A1(n361), .A2(n714), .ZN(n421) );
  INV_X1 U490 ( .A(G122), .ZN(n564) );
  AND2_X1 U491 ( .A1(n397), .A2(n392), .ZN(n356) );
  XOR2_X1 U492 ( .A(KEYINPUT23), .B(G110), .Z(n357) );
  XOR2_X1 U493 ( .A(n429), .B(n428), .Z(n358) );
  AND2_X1 U494 ( .A1(n424), .A2(n602), .ZN(n359) );
  NAND2_X1 U495 ( .A1(n386), .A2(n734), .ZN(n360) );
  OR2_X1 U496 ( .A1(n713), .A2(n712), .ZN(n361) );
  AND2_X1 U497 ( .A1(n398), .A2(n356), .ZN(n362) );
  AND2_X1 U498 ( .A1(n643), .A2(KEYINPUT2), .ZN(n363) );
  XOR2_X1 U499 ( .A(n532), .B(KEYINPUT73), .Z(n364) );
  OR2_X1 U500 ( .A1(n622), .A2(KEYINPUT47), .ZN(n365) );
  INV_X1 U501 ( .A(n702), .ZN(n392) );
  XNOR2_X2 U502 ( .A(n366), .B(n506), .ZN(n508) );
  XNOR2_X2 U503 ( .A(n504), .B(n503), .ZN(n366) );
  XNOR2_X2 U504 ( .A(n587), .B(KEYINPUT32), .ZN(n782) );
  XNOR2_X2 U505 ( .A(n367), .B(G122), .ZN(n503) );
  NOR2_X2 U506 ( .A1(n368), .A2(n593), .ZN(n594) );
  NAND2_X1 U507 ( .A1(n782), .A2(n592), .ZN(n368) );
  XNOR2_X2 U508 ( .A(n369), .B(KEYINPUT45), .ZN(n598) );
  NAND2_X1 U509 ( .A1(n595), .A2(n596), .ZN(n369) );
  NAND2_X1 U510 ( .A1(n370), .A2(n439), .ZN(n563) );
  XNOR2_X1 U511 ( .A(n561), .B(n371), .ZN(n370) );
  NAND2_X1 U512 ( .A1(n372), .A2(n363), .ZN(n426) );
  NAND2_X1 U513 ( .A1(n655), .A2(n388), .ZN(n377) );
  NAND2_X1 U514 ( .A1(n380), .A2(n378), .ZN(n480) );
  AND2_X1 U515 ( .A1(n390), .A2(n473), .ZN(n379) );
  NOR2_X1 U516 ( .A1(n472), .A2(G902), .ZN(n388) );
  INV_X1 U517 ( .A(n472), .ZN(n391) );
  NAND2_X1 U518 ( .A1(n362), .A2(n393), .ZN(n399) );
  NAND2_X1 U519 ( .A1(n394), .A2(n393), .ZN(n565) );
  NOR2_X1 U520 ( .A1(n530), .A2(n364), .ZN(n395) );
  INV_X1 U521 ( .A(n531), .ZN(n396) );
  NAND2_X1 U522 ( .A1(n530), .A2(n364), .ZN(n397) );
  NAND2_X1 U523 ( .A1(n531), .A2(n364), .ZN(n398) );
  NAND2_X1 U524 ( .A1(n621), .A2(n622), .ZN(n400) );
  NAND2_X1 U525 ( .A1(n402), .A2(n401), .ZN(n624) );
  OR2_X1 U526 ( .A1(n621), .A2(n365), .ZN(n401) );
  AND2_X1 U527 ( .A1(n404), .A2(KEYINPUT80), .ZN(n403) );
  NAND2_X1 U528 ( .A1(n622), .A2(KEYINPUT47), .ZN(n404) );
  XNOR2_X1 U529 ( .A(n419), .B(n418), .ZN(G75) );
  NAND2_X1 U530 ( .A1(n359), .A2(n752), .ZN(n605) );
  NAND2_X1 U531 ( .A1(n735), .A2(n734), .ZN(n738) );
  XNOR2_X1 U532 ( .A(n426), .B(KEYINPUT85), .ZN(n648) );
  INV_X1 U533 ( .A(n598), .ZN(n647) );
  XNOR2_X1 U534 ( .A(n431), .B(n599), .ZN(n644) );
  NAND2_X1 U535 ( .A1(n598), .A2(n597), .ZN(n431) );
  NAND2_X1 U536 ( .A1(n597), .A2(KEYINPUT2), .ZN(n438) );
  XOR2_X1 U537 ( .A(n562), .B(KEYINPUT78), .Z(n439) );
  NOR2_X1 U538 ( .A1(n720), .A2(n585), .ZN(n440) );
  INV_X1 U539 ( .A(KEYINPUT76), .ZN(n622) );
  INV_X1 U540 ( .A(n645), .ZN(n597) );
  INV_X1 U541 ( .A(KEYINPUT84), .ZN(n599) );
  XNOR2_X1 U542 ( .A(n469), .B(n507), .ZN(n470) );
  INV_X1 U543 ( .A(KEYINPUT19), .ZN(n544) );
  INV_X1 U544 ( .A(n719), .ZN(n568) );
  NOR2_X1 U545 ( .A1(n737), .A2(n568), .ZN(n569) );
  INV_X1 U546 ( .A(KEYINPUT22), .ZN(n571) );
  NAND2_X1 U547 ( .A1(G234), .A2(n509), .ZN(n442) );
  NAND2_X1 U548 ( .A1(G221), .A2(n493), .ZN(n443) );
  NOR2_X1 U549 ( .A1(G902), .A2(n687), .ZN(n448) );
  XNOR2_X1 U550 ( .A(G902), .B(KEYINPUT15), .ZN(n645) );
  NAND2_X1 U551 ( .A1(G234), .A2(n645), .ZN(n444) );
  XNOR2_X1 U552 ( .A(KEYINPUT20), .B(n444), .ZN(n449) );
  NAND2_X1 U553 ( .A1(n449), .A2(G217), .ZN(n446) );
  XNOR2_X1 U554 ( .A(KEYINPUT95), .B(KEYINPUT25), .ZN(n445) );
  NAND2_X1 U555 ( .A1(n449), .A2(G221), .ZN(n450) );
  XOR2_X1 U556 ( .A(KEYINPUT21), .B(n450), .Z(n719) );
  XNOR2_X2 U557 ( .A(G143), .B(G128), .ZN(n497) );
  INV_X1 U558 ( .A(KEYINPUT4), .ZN(n452) );
  INV_X1 U559 ( .A(G134), .ZN(n453) );
  XNOR2_X1 U560 ( .A(n453), .B(G131), .ZN(n454) );
  XNOR2_X1 U561 ( .A(n455), .B(KEYINPUT93), .ZN(n456) );
  NAND2_X1 U562 ( .A1(n509), .A2(G227), .ZN(n457) );
  XNOR2_X1 U563 ( .A(n457), .B(KEYINPUT94), .ZN(n458) );
  XNOR2_X1 U564 ( .A(n458), .B(n518), .ZN(n462) );
  XNOR2_X1 U565 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U566 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U567 ( .A(n771), .B(n463), .ZN(n662) );
  NAND2_X1 U568 ( .A1(n716), .A2(n602), .ZN(n575) );
  INV_X1 U569 ( .A(n575), .ZN(n482) );
  XNOR2_X1 U570 ( .A(n466), .B(n465), .ZN(n471) );
  XNOR2_X1 U571 ( .A(n468), .B(n467), .ZN(n507) );
  INV_X1 U572 ( .A(G902), .ZN(n500) );
  XNOR2_X1 U573 ( .A(G472), .B(KEYINPUT74), .ZN(n472) );
  OR2_X1 U574 ( .A1(G237), .A2(G902), .ZN(n522) );
  NAND2_X1 U575 ( .A1(G214), .A2(n522), .ZN(n734) );
  XNOR2_X1 U576 ( .A(KEYINPUT108), .B(KEYINPUT30), .ZN(n473) );
  XOR2_X1 U577 ( .A(KEYINPUT14), .B(KEYINPUT91), .Z(n475) );
  XNOR2_X1 U578 ( .A(n475), .B(n474), .ZN(n476) );
  NAND2_X1 U579 ( .A1(G952), .A2(n476), .ZN(n749) );
  NOR2_X1 U580 ( .A1(G953), .A2(n749), .ZN(n548) );
  AND2_X1 U581 ( .A1(G953), .A2(n476), .ZN(n477) );
  NAND2_X1 U582 ( .A1(G902), .A2(n477), .ZN(n546) );
  NOR2_X1 U583 ( .A1(G900), .A2(n546), .ZN(n478) );
  OR2_X1 U584 ( .A1(n548), .A2(n478), .ZN(n479) );
  XNOR2_X1 U585 ( .A(n479), .B(KEYINPUT79), .ZN(n533) );
  NOR2_X1 U586 ( .A1(n480), .A2(n533), .ZN(n481) );
  NAND2_X1 U587 ( .A1(n482), .A2(n481), .ZN(n531) );
  XOR2_X1 U588 ( .A(G140), .B(KEYINPUT12), .Z(n488) );
  NAND2_X1 U589 ( .A1(G214), .A2(n486), .ZN(n487) );
  XNOR2_X1 U590 ( .A(n488), .B(n487), .ZN(n489) );
  NOR2_X1 U591 ( .A1(G902), .A2(n677), .ZN(n491) );
  XNOR2_X1 U592 ( .A(KEYINPUT102), .B(KEYINPUT13), .ZN(n490) );
  INV_X1 U593 ( .A(G475), .ZN(n492) );
  XOR2_X1 U594 ( .A(G134), .B(KEYINPUT9), .Z(n494) );
  INV_X1 U595 ( .A(KEYINPUT103), .ZN(n495) );
  XNOR2_X1 U596 ( .A(n495), .B(G116), .ZN(n496) );
  XNOR2_X1 U597 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U598 ( .A(n498), .B(n503), .ZN(n499) );
  XNOR2_X1 U599 ( .A(n358), .B(n499), .ZN(n652) );
  NAND2_X1 U600 ( .A1(n652), .A2(n500), .ZN(n502) );
  INV_X1 U601 ( .A(G478), .ZN(n501) );
  OR2_X1 U602 ( .A1(n567), .A2(n566), .ZN(n562) );
  INV_X1 U603 ( .A(n562), .ZN(n527) );
  XNOR2_X2 U604 ( .A(n508), .B(n507), .ZN(n763) );
  NAND2_X1 U605 ( .A1(G224), .A2(n509), .ZN(n515) );
  INV_X1 U606 ( .A(KEYINPUT18), .ZN(n510) );
  NAND2_X1 U607 ( .A1(n510), .A2(KEYINPUT17), .ZN(n513) );
  NAND2_X1 U608 ( .A1(n511), .A2(KEYINPUT18), .ZN(n512) );
  NAND2_X1 U609 ( .A1(n513), .A2(n512), .ZN(n514) );
  XNOR2_X1 U610 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U611 ( .A(n521), .B(n763), .ZN(n667) );
  NAND2_X1 U612 ( .A1(n667), .A2(n645), .ZN(n526) );
  INV_X1 U613 ( .A(n522), .ZN(n524) );
  INV_X1 U614 ( .A(G210), .ZN(n523) );
  NOR2_X1 U615 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X2 U616 ( .A(n526), .B(n525), .ZN(n543) );
  AND2_X1 U617 ( .A1(n543), .A2(n527), .ZN(n528) );
  NAND2_X1 U618 ( .A1(n396), .A2(n528), .ZN(n618) );
  XNOR2_X1 U619 ( .A(n618), .B(G143), .ZN(G45) );
  INV_X1 U620 ( .A(KEYINPUT38), .ZN(n529) );
  XNOR2_X1 U621 ( .A(n543), .B(n529), .ZN(n735) );
  INV_X1 U622 ( .A(n735), .ZN(n530) );
  XNOR2_X1 U623 ( .A(KEYINPUT87), .B(KEYINPUT39), .ZN(n532) );
  INV_X1 U624 ( .A(n566), .ZN(n536) );
  NAND2_X1 U625 ( .A1(n567), .A2(n536), .ZN(n698) );
  OR2_X1 U626 ( .A1(n565), .A2(n698), .ZN(n643) );
  XNOR2_X1 U627 ( .A(n643), .B(G134), .ZN(G36) );
  NOR2_X1 U628 ( .A1(n568), .A2(n533), .ZN(n534) );
  NAND2_X1 U629 ( .A1(n588), .A2(n534), .ZN(n535) );
  XOR2_X1 U630 ( .A(KEYINPUT71), .B(n535), .Z(n600) );
  INV_X1 U631 ( .A(KEYINPUT6), .ZN(n537) );
  XNOR2_X1 U632 ( .A(n726), .B(n537), .ZN(n585) );
  NAND2_X1 U633 ( .A1(n734), .A2(n585), .ZN(n538) );
  INV_X1 U634 ( .A(n543), .ZN(n637) );
  XNOR2_X1 U635 ( .A(n539), .B(KEYINPUT36), .ZN(n541) );
  XNOR2_X1 U636 ( .A(KEYINPUT66), .B(KEYINPUT1), .ZN(n540) );
  NAND2_X1 U637 ( .A1(n541), .A2(n355), .ZN(n625) );
  XOR2_X1 U638 ( .A(G125), .B(KEYINPUT37), .Z(n542) );
  XNOR2_X1 U639 ( .A(n625), .B(n542), .ZN(G27) );
  NAND2_X1 U640 ( .A1(n543), .A2(n734), .ZN(n545) );
  NOR2_X1 U641 ( .A1(G898), .A2(n546), .ZN(n547) );
  NOR2_X1 U642 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U643 ( .A(n549), .B(KEYINPUT92), .ZN(n550) );
  XNOR2_X1 U644 ( .A(n551), .B(KEYINPUT0), .ZN(n570) );
  BUF_X1 U645 ( .A(n570), .Z(n577) );
  NAND2_X1 U646 ( .A1(n559), .A2(n726), .ZN(n552) );
  NAND2_X1 U647 ( .A1(n577), .A2(n728), .ZN(n554) );
  XNOR2_X1 U648 ( .A(KEYINPUT98), .B(KEYINPUT31), .ZN(n553) );
  XNOR2_X1 U649 ( .A(n554), .B(n553), .ZN(n579) );
  INV_X1 U650 ( .A(n698), .ZN(n555) );
  NAND2_X1 U651 ( .A1(n579), .A2(n555), .ZN(n556) );
  XNOR2_X1 U652 ( .A(n556), .B(G116), .ZN(G18) );
  XNOR2_X1 U653 ( .A(G113), .B(KEYINPUT113), .ZN(n558) );
  NAND2_X1 U654 ( .A1(n579), .A2(n392), .ZN(n557) );
  XOR2_X1 U655 ( .A(n558), .B(n557), .Z(G15) );
  NAND2_X1 U656 ( .A1(n559), .A2(n585), .ZN(n560) );
  XNOR2_X2 U657 ( .A(n560), .B(KEYINPUT33), .ZN(n751) );
  NAND2_X1 U658 ( .A1(n577), .A2(n751), .ZN(n561) );
  XNOR2_X1 U659 ( .A(n564), .B(n593), .ZN(G24) );
  XNOR2_X1 U660 ( .A(n606), .B(G131), .ZN(G33) );
  NAND2_X1 U661 ( .A1(n567), .A2(n566), .ZN(n737) );
  XNOR2_X1 U662 ( .A(n588), .B(KEYINPUT105), .ZN(n720) );
  NAND2_X1 U663 ( .A1(n573), .A2(n720), .ZN(n574) );
  NOR2_X1 U664 ( .A1(n575), .A2(n726), .ZN(n576) );
  NAND2_X1 U665 ( .A1(n577), .A2(n576), .ZN(n692) );
  INV_X1 U666 ( .A(n692), .ZN(n578) );
  INV_X1 U667 ( .A(KEYINPUT99), .ZN(n580) );
  XNOR2_X1 U668 ( .A(n581), .B(n580), .ZN(n583) );
  NAND2_X1 U669 ( .A1(n702), .A2(n698), .ZN(n612) );
  INV_X1 U670 ( .A(n621), .ZN(n582) );
  NAND2_X1 U671 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U672 ( .A1(n440), .A2(n355), .ZN(n586) );
  INV_X1 U673 ( .A(n726), .ZN(n601) );
  NAND2_X1 U674 ( .A1(n601), .A2(n588), .ZN(n589) );
  OR2_X1 U675 ( .A1(n355), .A2(n589), .ZN(n590) );
  NOR2_X1 U676 ( .A1(n591), .A2(n590), .ZN(n697) );
  INV_X1 U677 ( .A(n697), .ZN(n592) );
  XNOR2_X1 U678 ( .A(n594), .B(KEYINPUT44), .ZN(n595) );
  INV_X1 U679 ( .A(KEYINPUT109), .ZN(n603) );
  XNOR2_X1 U680 ( .A(n603), .B(KEYINPUT42), .ZN(n604) );
  XNOR2_X1 U681 ( .A(n605), .B(n604), .ZN(n783) );
  NAND2_X1 U682 ( .A1(n606), .A2(n783), .ZN(n609) );
  INV_X1 U683 ( .A(KEYINPUT64), .ZN(n607) );
  XNOR2_X1 U684 ( .A(n607), .B(KEYINPUT46), .ZN(n608) );
  XNOR2_X1 U685 ( .A(n609), .B(n608), .ZN(n630) );
  INV_X1 U686 ( .A(n610), .ZN(n611) );
  NAND2_X1 U687 ( .A1(n359), .A2(n611), .ZN(n701) );
  NAND2_X1 U688 ( .A1(n701), .A2(KEYINPUT80), .ZN(n614) );
  AND2_X1 U689 ( .A1(n612), .A2(KEYINPUT47), .ZN(n613) );
  NAND2_X1 U690 ( .A1(n614), .A2(n613), .ZN(n617) );
  INV_X1 U691 ( .A(KEYINPUT47), .ZN(n615) );
  NAND2_X1 U692 ( .A1(n615), .A2(KEYINPUT80), .ZN(n616) );
  NAND2_X1 U693 ( .A1(n617), .A2(n616), .ZN(n620) );
  XNOR2_X1 U694 ( .A(n618), .B(KEYINPUT82), .ZN(n619) );
  NAND2_X1 U695 ( .A1(n620), .A2(n619), .ZN(n628) );
  INV_X1 U696 ( .A(n701), .ZN(n623) );
  NAND2_X1 U697 ( .A1(n624), .A2(n623), .ZN(n626) );
  NAND2_X1 U698 ( .A1(n626), .A2(n625), .ZN(n627) );
  NAND2_X1 U699 ( .A1(n630), .A2(n629), .ZN(n632) );
  INV_X1 U700 ( .A(KEYINPUT48), .ZN(n631) );
  XNOR2_X1 U701 ( .A(n632), .B(n631), .ZN(n640) );
  XOR2_X1 U702 ( .A(KEYINPUT107), .B(n633), .Z(n634) );
  NOR2_X1 U703 ( .A1(n634), .A2(n355), .ZN(n636) );
  INV_X1 U704 ( .A(KEYINPUT43), .ZN(n635) );
  XNOR2_X1 U705 ( .A(n636), .B(n635), .ZN(n638) );
  AND2_X1 U706 ( .A1(n638), .A2(n637), .ZN(n705) );
  INV_X1 U707 ( .A(n705), .ZN(n639) );
  NAND2_X1 U708 ( .A1(n640), .A2(n639), .ZN(n642) );
  INV_X1 U709 ( .A(KEYINPUT86), .ZN(n641) );
  NAND2_X1 U710 ( .A1(n644), .A2(n706), .ZN(n646) );
  NAND2_X1 U711 ( .A1(n646), .A2(n438), .ZN(n649) );
  NAND2_X1 U712 ( .A1(n648), .A2(n598), .ZN(n714) );
  NAND2_X1 U713 ( .A1(n649), .A2(n714), .ZN(n650) );
  XNOR2_X2 U714 ( .A(n650), .B(KEYINPUT65), .ZN(n684) );
  NAND2_X1 U715 ( .A1(n684), .A2(G478), .ZN(n651) );
  XOR2_X1 U716 ( .A(n652), .B(n651), .Z(n654) );
  INV_X1 U717 ( .A(G952), .ZN(n653) );
  NAND2_X1 U718 ( .A1(n653), .A2(G953), .ZN(n680) );
  INV_X1 U719 ( .A(n680), .ZN(n688) );
  NOR2_X1 U720 ( .A1(n654), .A2(n688), .ZN(G63) );
  NAND2_X1 U721 ( .A1(n684), .A2(G472), .ZN(n657) );
  XNOR2_X1 U722 ( .A(n655), .B(KEYINPUT62), .ZN(n656) );
  XNOR2_X1 U723 ( .A(n657), .B(n656), .ZN(n658) );
  NAND2_X1 U724 ( .A1(n658), .A2(n680), .ZN(n660) );
  XNOR2_X1 U725 ( .A(KEYINPUT90), .B(KEYINPUT63), .ZN(n659) );
  XNOR2_X1 U726 ( .A(n660), .B(n659), .ZN(G57) );
  NAND2_X1 U727 ( .A1(n684), .A2(G469), .ZN(n664) );
  XNOR2_X1 U728 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n661) );
  XNOR2_X1 U729 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U730 ( .A(n664), .B(n663), .ZN(n665) );
  NAND2_X1 U731 ( .A1(n665), .A2(n680), .ZN(n666) );
  XNOR2_X1 U732 ( .A(n666), .B(KEYINPUT121), .ZN(G54) );
  INV_X1 U733 ( .A(KEYINPUT56), .ZN(n674) );
  NAND2_X1 U734 ( .A1(n684), .A2(G210), .ZN(n671) );
  BUF_X1 U735 ( .A(n667), .Z(n669) );
  XOR2_X1 U736 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n668) );
  XNOR2_X1 U737 ( .A(n669), .B(n668), .ZN(n670) );
  XNOR2_X1 U738 ( .A(n671), .B(n670), .ZN(n672) );
  NAND2_X1 U739 ( .A1(n672), .A2(n680), .ZN(n673) );
  XNOR2_X1 U740 ( .A(n674), .B(n673), .ZN(G51) );
  NAND2_X1 U741 ( .A1(n684), .A2(G475), .ZN(n679) );
  XNOR2_X1 U742 ( .A(KEYINPUT67), .B(KEYINPUT89), .ZN(n675) );
  XNOR2_X1 U743 ( .A(n675), .B(KEYINPUT59), .ZN(n676) );
  XNOR2_X1 U744 ( .A(n677), .B(n676), .ZN(n678) );
  XNOR2_X1 U745 ( .A(n679), .B(n678), .ZN(n681) );
  NAND2_X1 U746 ( .A1(n681), .A2(n680), .ZN(n683) );
  XOR2_X1 U747 ( .A(KEYINPUT68), .B(KEYINPUT60), .Z(n682) );
  XNOR2_X1 U748 ( .A(n683), .B(n682), .ZN(G60) );
  BUF_X1 U749 ( .A(n684), .Z(n685) );
  NAND2_X1 U750 ( .A1(n685), .A2(G217), .ZN(n686) );
  XNOR2_X1 U751 ( .A(n687), .B(n686), .ZN(n689) );
  NOR2_X1 U752 ( .A1(n689), .A2(n688), .ZN(G66) );
  NOR2_X1 U753 ( .A1(n702), .A2(n692), .ZN(n690) );
  XOR2_X1 U754 ( .A(KEYINPUT110), .B(n690), .Z(n691) );
  XNOR2_X1 U755 ( .A(G104), .B(n691), .ZN(G6) );
  NOR2_X1 U756 ( .A1(n692), .A2(n698), .ZN(n696) );
  XOR2_X1 U757 ( .A(KEYINPUT111), .B(KEYINPUT27), .Z(n694) );
  XNOR2_X1 U758 ( .A(G107), .B(KEYINPUT26), .ZN(n693) );
  XNOR2_X1 U759 ( .A(n694), .B(n693), .ZN(n695) );
  XNOR2_X1 U760 ( .A(n696), .B(n695), .ZN(G9) );
  XOR2_X1 U761 ( .A(G110), .B(n697), .Z(G12) );
  NOR2_X1 U762 ( .A1(n698), .A2(n701), .ZN(n700) );
  XNOR2_X1 U763 ( .A(G128), .B(KEYINPUT29), .ZN(n699) );
  XNOR2_X1 U764 ( .A(n700), .B(n699), .ZN(G30) );
  OR2_X1 U765 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U766 ( .A(n703), .B(KEYINPUT112), .ZN(n704) );
  XNOR2_X1 U767 ( .A(G146), .B(n704), .ZN(G48) );
  XOR2_X1 U768 ( .A(G140), .B(n705), .Z(G42) );
  NOR2_X1 U769 ( .A1(n647), .A2(n777), .ZN(n707) );
  NOR2_X1 U770 ( .A1(n707), .A2(KEYINPUT2), .ZN(n708) );
  NOR2_X1 U771 ( .A1(n708), .A2(KEYINPUT83), .ZN(n713) );
  INV_X1 U772 ( .A(KEYINPUT83), .ZN(n709) );
  NOR2_X1 U773 ( .A1(n709), .A2(KEYINPUT2), .ZN(n710) );
  NAND2_X1 U774 ( .A1(n777), .A2(n710), .ZN(n711) );
  NOR2_X1 U775 ( .A1(n647), .A2(n711), .ZN(n712) );
  INV_X1 U776 ( .A(n752), .ZN(n733) );
  XOR2_X1 U777 ( .A(KEYINPUT115), .B(KEYINPUT50), .Z(n718) );
  NOR2_X1 U778 ( .A1(n716), .A2(n355), .ZN(n717) );
  XOR2_X1 U779 ( .A(n718), .B(n717), .Z(n724) );
  NOR2_X1 U780 ( .A1(n720), .A2(n719), .ZN(n722) );
  XNOR2_X1 U781 ( .A(KEYINPUT114), .B(KEYINPUT49), .ZN(n721) );
  XNOR2_X1 U782 ( .A(n722), .B(n721), .ZN(n723) );
  NAND2_X1 U783 ( .A1(n724), .A2(n723), .ZN(n725) );
  NOR2_X1 U784 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U785 ( .A(n727), .B(KEYINPUT116), .ZN(n729) );
  NOR2_X1 U786 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U787 ( .A(n730), .B(KEYINPUT117), .ZN(n731) );
  XNOR2_X1 U788 ( .A(KEYINPUT51), .B(n731), .ZN(n732) );
  NOR2_X1 U789 ( .A1(n733), .A2(n732), .ZN(n746) );
  NOR2_X1 U790 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U791 ( .A1(n737), .A2(n736), .ZN(n742) );
  INV_X1 U792 ( .A(n612), .ZN(n739) );
  NOR2_X1 U793 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U794 ( .A(n740), .B(KEYINPUT118), .ZN(n741) );
  NOR2_X1 U795 ( .A1(n742), .A2(n741), .ZN(n744) );
  INV_X1 U796 ( .A(n751), .ZN(n743) );
  NOR2_X1 U797 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U798 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U799 ( .A(n747), .B(KEYINPUT52), .ZN(n748) );
  NOR2_X1 U800 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U801 ( .A(n750), .B(KEYINPUT119), .ZN(n754) );
  NAND2_X1 U802 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U803 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U804 ( .A(n755), .B(KEYINPUT120), .ZN(n756) );
  NOR2_X1 U805 ( .A1(n647), .A2(G953), .ZN(n762) );
  NAND2_X1 U806 ( .A1(G224), .A2(G953), .ZN(n757) );
  XNOR2_X1 U807 ( .A(n757), .B(KEYINPUT122), .ZN(n758) );
  XNOR2_X1 U808 ( .A(KEYINPUT61), .B(n758), .ZN(n759) );
  NAND2_X1 U809 ( .A1(n759), .A2(G898), .ZN(n760) );
  XNOR2_X1 U810 ( .A(n760), .B(KEYINPUT123), .ZN(n761) );
  NOR2_X1 U811 ( .A1(n762), .A2(n761), .ZN(n768) );
  XNOR2_X1 U812 ( .A(n763), .B(G110), .ZN(n764) );
  XNOR2_X1 U813 ( .A(n764), .B(KEYINPUT124), .ZN(n766) );
  NOR2_X1 U814 ( .A1(G898), .A2(n509), .ZN(n765) );
  NOR2_X1 U815 ( .A1(n766), .A2(n765), .ZN(n767) );
  XOR2_X1 U816 ( .A(n768), .B(n767), .Z(G69) );
  XNOR2_X1 U817 ( .A(n769), .B(KEYINPUT125), .ZN(n770) );
  XOR2_X1 U818 ( .A(n771), .B(n770), .Z(n775) );
  XOR2_X1 U819 ( .A(G227), .B(n775), .Z(n772) );
  NAND2_X1 U820 ( .A1(n772), .A2(G900), .ZN(n773) );
  NAND2_X1 U821 ( .A1(G953), .A2(n773), .ZN(n774) );
  XOR2_X1 U822 ( .A(KEYINPUT127), .B(n774), .Z(n780) );
  XOR2_X1 U823 ( .A(n775), .B(KEYINPUT126), .Z(n776) );
  XNOR2_X1 U824 ( .A(n777), .B(n776), .ZN(n778) );
  NAND2_X1 U825 ( .A1(n778), .A2(n509), .ZN(n779) );
  NAND2_X1 U826 ( .A1(n780), .A2(n779), .ZN(G72) );
  XNOR2_X1 U827 ( .A(n781), .B(G101), .ZN(G3) );
  XNOR2_X1 U828 ( .A(n782), .B(G119), .ZN(G21) );
  XNOR2_X1 U829 ( .A(G137), .B(n783), .ZN(G39) );
endmodule

