//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 0 0 0 0 0 1 0 1 1 0 1 0 1 1 0 1 0 1 0 1 1 1 0 1 0 1 0 1 0 0 1 1 0 1 0 0 1 0 1 0 0 1 1 0 0 1 0 1 0 0 1 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n611, new_n612, new_n613, new_n614, new_n616, new_n617,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n646, new_n647,
    new_n649, new_n650, new_n651, new_n652, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n766, new_n767, new_n768, new_n770, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n848, new_n849, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n858, new_n859, new_n861, new_n862, new_n863, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906;
  NAND2_X1  g000(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n202));
  MUX2_X1   g001(.A(G183gat), .B(new_n202), .S(G190gat), .Z(new_n203));
  INV_X1    g002(.A(KEYINPUT24), .ZN(new_n204));
  INV_X1    g003(.A(G183gat), .ZN(new_n205));
  INV_X1    g004(.A(G190gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n203), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G169gat), .ZN(new_n209));
  INV_X1    g008(.A(G176gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n209), .A2(new_n210), .A3(KEYINPUT23), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT23), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n212), .B1(G169gat), .B2(G176gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n211), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  AOI21_X1  g015(.A(KEYINPUT25), .B1(new_n208), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT65), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n207), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(new_n203), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n207), .A2(new_n218), .ZN(new_n221));
  OAI211_X1 g020(.A(KEYINPUT25), .B(new_n216), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  OR2_X1    g021(.A1(new_n222), .A2(KEYINPUT66), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(KEYINPUT66), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n217), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  XOR2_X1   g024(.A(G127gat), .B(G134gat), .Z(new_n226));
  XNOR2_X1  g025(.A(G113gat), .B(G120gat), .ZN(new_n227));
  AND2_X1   g026(.A1(new_n227), .A2(KEYINPUT68), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT1), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n229), .B1(new_n227), .B2(KEYINPUT68), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n226), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(G120gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(G113gat), .ZN(new_n233));
  XOR2_X1   g032(.A(KEYINPUT69), .B(G113gat), .Z(new_n234));
  OAI21_X1  g033(.A(new_n233), .B1(new_n234), .B2(new_n232), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n226), .A2(KEYINPUT1), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  AND2_X1   g036(.A1(new_n231), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(KEYINPUT27), .B(G183gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(new_n206), .ZN(new_n240));
  OR2_X1    g039(.A1(new_n240), .A2(KEYINPUT28), .ZN(new_n241));
  AOI22_X1  g040(.A1(new_n240), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n209), .A2(new_n210), .A3(KEYINPUT67), .ZN(new_n243));
  OR2_X1    g042(.A1(new_n243), .A2(KEYINPUT26), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(KEYINPUT26), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n244), .A2(new_n214), .A3(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n241), .A2(new_n242), .A3(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  OR3_X1    g047(.A1(new_n225), .A2(new_n238), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(G227gat), .A2(G233gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(KEYINPUT64), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n238), .B1(new_n225), .B2(new_n248), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n249), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(KEYINPUT32), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n251), .B1(new_n249), .B2(new_n252), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT34), .ZN(new_n257));
  AND2_X1   g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(G15gat), .B(G43gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(G71gat), .B(G99gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n259), .B(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT33), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n261), .B1(new_n253), .B2(new_n262), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n256), .A2(new_n257), .ZN(new_n264));
  NOR3_X1   g063(.A1(new_n258), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n263), .B1(new_n258), .B2(new_n264), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n255), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n266), .A2(new_n255), .A3(new_n267), .ZN(new_n270));
  AOI21_X1  g069(.A(KEYINPUT36), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n267), .ZN(new_n272));
  NOR3_X1   g071(.A1(new_n272), .A2(new_n265), .A3(new_n254), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT36), .ZN(new_n274));
  NOR3_X1   g073(.A1(new_n268), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n271), .A2(new_n275), .ZN(new_n276));
  XOR2_X1   g075(.A(G1gat), .B(G29gat), .Z(new_n277));
  XNOR2_X1  g076(.A(G57gat), .B(G85gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(KEYINPUT75), .B(KEYINPUT0), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n283));
  NAND2_X1  g082(.A1(G155gat), .A2(G162gat), .ZN(new_n284));
  INV_X1    g083(.A(G155gat), .ZN(new_n285));
  INV_X1    g084(.A(G162gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n284), .B1(new_n287), .B2(KEYINPUT2), .ZN(new_n288));
  INV_X1    g087(.A(G141gat), .ZN(new_n289));
  OAI21_X1  g088(.A(KEYINPUT70), .B1(new_n289), .B2(G148gat), .ZN(new_n290));
  INV_X1    g089(.A(G148gat), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n290), .B1(G141gat), .B2(new_n291), .ZN(new_n292));
  NOR3_X1   g091(.A1(new_n289), .A2(KEYINPUT70), .A3(G148gat), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n288), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(G141gat), .B(G148gat), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n284), .B(new_n287), .C1(new_n295), .C2(KEYINPUT2), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n238), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT73), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n299), .B(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n238), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(new_n297), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(G225gat), .A2(G233gat), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n305), .B(KEYINPUT71), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n283), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT3), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n298), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n297), .A2(KEYINPUT3), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n302), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n306), .ZN(new_n313));
  AND2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n301), .A2(KEYINPUT4), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n299), .A2(KEYINPUT4), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n316), .B(KEYINPUT72), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n314), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT74), .ZN(new_n319));
  OR2_X1    g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n318), .A2(new_n319), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n308), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n299), .ZN(new_n323));
  MUX2_X1   g122(.A(new_n323), .B(new_n301), .S(KEYINPUT4), .Z(new_n324));
  NAND3_X1  g123(.A1(new_n324), .A2(new_n283), .A3(new_n314), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n282), .B1(new_n322), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT6), .ZN(new_n328));
  OAI21_X1  g127(.A(KEYINPUT76), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n320), .A2(new_n321), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(new_n307), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n331), .A2(new_n281), .A3(new_n325), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n332), .A2(new_n327), .A3(new_n328), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n331), .A2(new_n325), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT76), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n334), .A2(new_n335), .A3(KEYINPUT6), .A4(new_n282), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n329), .A2(new_n333), .A3(new_n336), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n225), .A2(new_n248), .ZN(new_n338));
  NAND2_X1  g137(.A1(G226gat), .A2(G233gat), .ZN(new_n339));
  OR2_X1    g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(G197gat), .B(G204gat), .ZN(new_n341));
  AND2_X1   g140(.A1(G211gat), .A2(G218gat), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n341), .B1(KEYINPUT22), .B2(new_n342), .ZN(new_n343));
  NOR2_X1   g142(.A1(G211gat), .A2(G218gat), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n343), .B(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n339), .B1(new_n338), .B2(KEYINPUT29), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n340), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n346), .B1(new_n340), .B2(new_n347), .ZN(new_n350));
  XNOR2_X1  g149(.A(G8gat), .B(G36gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(G64gat), .B(G92gat), .ZN(new_n352));
  XOR2_X1   g151(.A(new_n351), .B(new_n352), .Z(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  OR4_X1    g153(.A1(KEYINPUT30), .A2(new_n349), .A3(new_n350), .A4(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n354), .B1(new_n349), .B2(new_n350), .ZN(new_n356));
  INV_X1    g155(.A(new_n350), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n357), .A2(new_n348), .A3(new_n353), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n356), .A2(new_n358), .A3(KEYINPUT30), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n355), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n337), .A2(new_n360), .ZN(new_n361));
  XOR2_X1   g160(.A(G78gat), .B(G106gat), .Z(new_n362));
  XNOR2_X1  g161(.A(KEYINPUT31), .B(G50gat), .ZN(new_n363));
  XOR2_X1   g162(.A(new_n362), .B(new_n363), .Z(new_n364));
  INV_X1    g163(.A(KEYINPUT29), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n346), .B1(new_n310), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n346), .A2(new_n365), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n298), .B1(new_n367), .B2(new_n309), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(G228gat), .A2(G233gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n369), .B(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(G22gat), .ZN(new_n372));
  AND2_X1   g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n364), .B1(new_n373), .B2(KEYINPUT77), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n371), .B(new_n372), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n374), .B(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n276), .B1(new_n361), .B2(new_n377), .ZN(new_n378));
  OR3_X1    g177(.A1(new_n349), .A2(KEYINPUT37), .A3(new_n350), .ZN(new_n379));
  OAI21_X1  g178(.A(KEYINPUT37), .B1(new_n349), .B2(new_n350), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n379), .A2(new_n354), .A3(new_n380), .ZN(new_n381));
  OR2_X1    g180(.A1(new_n381), .A2(KEYINPUT38), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(KEYINPUT38), .ZN(new_n383));
  AND3_X1   g182(.A1(new_n382), .A2(new_n358), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT79), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n334), .A2(new_n385), .A3(new_n282), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n327), .A2(KEYINPUT79), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n386), .A2(new_n387), .A3(new_n328), .A4(new_n332), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n384), .A2(new_n388), .A3(new_n336), .A4(new_n329), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n327), .B(new_n385), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n313), .B1(new_n324), .B2(new_n312), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT39), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n301), .A2(new_n313), .A3(new_n303), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n394), .B(KEYINPUT78), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n282), .B1(new_n391), .B2(new_n392), .ZN(new_n397));
  AND3_X1   g196(.A1(new_n396), .A2(KEYINPUT40), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT40), .B1(new_n396), .B2(new_n397), .ZN(new_n399));
  NOR3_X1   g198(.A1(new_n398), .A2(new_n399), .A3(new_n360), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n377), .B1(new_n390), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n389), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n337), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n269), .A2(new_n376), .A3(new_n360), .A4(new_n270), .ZN(new_n404));
  OAI21_X1  g203(.A(KEYINPUT35), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n388), .A2(new_n336), .A3(new_n329), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n404), .A2(KEYINPUT35), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AOI22_X1  g207(.A1(new_n378), .A2(new_n402), .B1(new_n405), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(G50gat), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(G43gat), .ZN(new_n411));
  INV_X1    g210(.A(G43gat), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(G50gat), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT15), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  OR3_X1    g215(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n417));
  OAI21_X1  g216(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n411), .A2(new_n413), .A3(KEYINPUT15), .ZN(new_n420));
  NAND2_X1  g219(.A1(G29gat), .A2(G36gat), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n416), .A2(new_n419), .A3(new_n420), .A4(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n418), .A2(KEYINPUT81), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT81), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n424), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n423), .A2(new_n417), .A3(new_n425), .ZN(new_n426));
  AND2_X1   g225(.A1(new_n426), .A2(new_n421), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n422), .B1(new_n427), .B2(new_n420), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(G1gat), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(KEYINPUT16), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n372), .A2(G15gat), .ZN(new_n432));
  INV_X1    g231(.A(G15gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(G22gat), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n431), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  XNOR2_X1  g234(.A(G15gat), .B(G22gat), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n435), .B1(G1gat), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(G8gat), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT83), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n439), .B1(new_n436), .B2(G1gat), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n437), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  OAI221_X1 g240(.A(new_n435), .B1(new_n439), .B2(G8gat), .C1(G1gat), .C2(new_n436), .ZN(new_n442));
  AND3_X1   g241(.A1(new_n441), .A2(KEYINPUT84), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT84), .B1(new_n441), .B2(new_n442), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n429), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n441), .A2(new_n442), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT84), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n441), .A2(KEYINPUT84), .A3(new_n442), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n448), .A2(new_n428), .A3(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n445), .A2(new_n450), .A3(KEYINPUT85), .ZN(new_n451));
  NAND2_X1  g250(.A1(G229gat), .A2(G233gat), .ZN(new_n452));
  XOR2_X1   g251(.A(new_n452), .B(KEYINPUT13), .Z(new_n453));
  INV_X1    g252(.A(KEYINPUT85), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n448), .A2(new_n454), .A3(new_n428), .A4(new_n449), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n451), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  OAI211_X1 g255(.A(KEYINPUT17), .B(new_n422), .C1(new_n427), .C2(new_n420), .ZN(new_n457));
  XOR2_X1   g256(.A(KEYINPUT82), .B(KEYINPUT17), .Z(new_n458));
  XNOR2_X1  g257(.A(G43gat), .B(G50gat), .ZN(new_n459));
  INV_X1    g258(.A(new_n418), .ZN(new_n460));
  NOR3_X1   g259(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n461));
  OAI22_X1  g260(.A1(new_n459), .A2(KEYINPUT15), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n420), .A2(new_n421), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n420), .B1(new_n426), .B2(new_n421), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n458), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n457), .A2(new_n466), .A3(new_n446), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n450), .A2(KEYINPUT18), .A3(new_n452), .A4(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n450), .A2(new_n452), .A3(new_n467), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT18), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n456), .A2(new_n468), .A3(new_n471), .ZN(new_n472));
  XNOR2_X1  g271(.A(G113gat), .B(G141gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(KEYINPUT80), .B(KEYINPUT11), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n473), .B(new_n474), .ZN(new_n475));
  XOR2_X1   g274(.A(G169gat), .B(G197gat), .Z(new_n476));
  XNOR2_X1  g275(.A(new_n475), .B(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n477), .B(KEYINPUT12), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n472), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT87), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n456), .A2(new_n468), .A3(new_n478), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT86), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n469), .A2(new_n484), .A3(new_n470), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n484), .B1(new_n469), .B2(new_n470), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n481), .B1(new_n483), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n471), .A2(KEYINPUT86), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(new_n485), .ZN(new_n491));
  NOR3_X1   g290(.A1(new_n491), .A2(new_n482), .A3(KEYINPUT87), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n480), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n409), .A2(new_n494), .ZN(new_n495));
  AND2_X1   g294(.A1(G71gat), .A2(G78gat), .ZN(new_n496));
  NOR2_X1   g295(.A1(G71gat), .A2(G78gat), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  XNOR2_X1  g297(.A(G57gat), .B(G64gat), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT9), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(G57gat), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n502), .A2(G64gat), .ZN(new_n503));
  XNOR2_X1  g302(.A(KEYINPUT88), .B(G57gat), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n503), .B1(new_n504), .B2(G64gat), .ZN(new_n505));
  NOR3_X1   g304(.A1(new_n500), .A2(G71gat), .A3(G78gat), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n506), .A2(new_n496), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n501), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT21), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(G231gat), .A2(G233gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n510), .B(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(G127gat), .B(G155gat), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n513), .B(KEYINPUT20), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n512), .B(new_n514), .ZN(new_n515));
  XOR2_X1   g314(.A(G183gat), .B(G211gat), .Z(new_n516));
  XNOR2_X1  g315(.A(new_n515), .B(new_n516), .ZN(new_n517));
  OAI22_X1  g316(.A1(new_n443), .A2(new_n444), .B1(new_n509), .B2(new_n508), .ZN(new_n518));
  XNOR2_X1  g317(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n519));
  XNOR2_X1  g318(.A(KEYINPUT89), .B(KEYINPUT90), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n518), .B(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n517), .B(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(G99gat), .B(G106gat), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(G85gat), .A2(G92gat), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT93), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT7), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(KEYINPUT93), .ZN(new_n531));
  AND3_X1   g330(.A1(new_n527), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n526), .A2(KEYINPUT93), .A3(new_n530), .ZN(new_n533));
  NOR2_X1   g332(.A1(G85gat), .A2(G92gat), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(G99gat), .A2(G106gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT8), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n533), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n525), .B1(new_n532), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n534), .B1(new_n540), .B2(new_n526), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n527), .A2(new_n529), .A3(new_n531), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n541), .A2(new_n542), .A3(new_n524), .A4(new_n537), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n539), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  AND2_X1   g344(.A1(G232gat), .A2(G233gat), .ZN(new_n546));
  AOI22_X1  g345(.A1(new_n428), .A2(new_n545), .B1(KEYINPUT41), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n457), .A2(new_n466), .A3(new_n544), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  XOR2_X1   g348(.A(G190gat), .B(G218gat), .Z(new_n550));
  AND2_X1   g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n546), .A2(KEYINPUT41), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(KEYINPUT92), .ZN(new_n553));
  XNOR2_X1  g352(.A(G134gat), .B(G162gat), .ZN(new_n554));
  XOR2_X1   g353(.A(new_n553), .B(new_n554), .Z(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n549), .A2(new_n550), .ZN(new_n557));
  OR4_X1    g356(.A1(KEYINPUT94), .A2(new_n551), .A3(new_n556), .A4(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n555), .B(KEYINPUT94), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n559), .B1(new_n551), .B2(new_n557), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n523), .A2(new_n561), .ZN(new_n562));
  XOR2_X1   g361(.A(G120gat), .B(G148gat), .Z(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(KEYINPUT96), .ZN(new_n564));
  XNOR2_X1  g363(.A(G176gat), .B(G204gat), .ZN(new_n565));
  XOR2_X1   g364(.A(new_n564), .B(new_n565), .Z(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT10), .ZN(new_n568));
  NOR3_X1   g367(.A1(new_n544), .A2(new_n568), .A3(new_n508), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n502), .A2(KEYINPUT88), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT88), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(G57gat), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n570), .A2(new_n572), .A3(G64gat), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n573), .B1(new_n502), .B2(G64gat), .ZN(new_n574));
  INV_X1    g373(.A(new_n507), .ZN(new_n575));
  AND2_X1   g374(.A1(new_n502), .A2(G64gat), .ZN(new_n576));
  OAI21_X1  g375(.A(KEYINPUT9), .B1(new_n576), .B2(new_n503), .ZN(new_n577));
  AOI22_X1  g376(.A1(new_n574), .A2(new_n575), .B1(new_n577), .B2(new_n498), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT95), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n543), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n544), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  OAI211_X1 g380(.A(new_n543), .B(new_n539), .C1(new_n508), .C2(new_n579), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n569), .B1(new_n583), .B2(new_n568), .ZN(new_n584));
  NAND2_X1  g383(.A1(G230gat), .A2(G233gat), .ZN(new_n585));
  XOR2_X1   g384(.A(new_n585), .B(KEYINPUT97), .Z(new_n586));
  OAI21_X1  g385(.A(KEYINPUT98), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT98), .ZN(new_n588));
  INV_X1    g387(.A(new_n586), .ZN(new_n589));
  AOI21_X1  g388(.A(KEYINPUT10), .B1(new_n581), .B2(new_n582), .ZN(new_n590));
  OAI211_X1 g389(.A(new_n588), .B(new_n589), .C1(new_n590), .C2(new_n569), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n583), .A2(new_n585), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n567), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n585), .B1(new_n590), .B2(new_n569), .ZN(new_n595));
  INV_X1    g394(.A(new_n593), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n595), .A2(new_n596), .A3(new_n566), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n562), .A2(new_n598), .ZN(new_n599));
  AND2_X1   g398(.A1(new_n495), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(new_n403), .ZN(new_n601));
  XOR2_X1   g400(.A(KEYINPUT99), .B(G1gat), .Z(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(G1324gat));
  INV_X1    g402(.A(new_n360), .ZN(new_n604));
  XOR2_X1   g403(.A(KEYINPUT16), .B(G8gat), .Z(new_n605));
  NAND3_X1  g404(.A1(new_n600), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n600), .ZN(new_n607));
  OAI21_X1  g406(.A(G8gat), .B1(new_n607), .B2(new_n360), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(new_n606), .ZN(new_n609));
  MUX2_X1   g408(.A(new_n606), .B(new_n609), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g409(.A(new_n276), .ZN(new_n611));
  OAI21_X1  g410(.A(G15gat), .B1(new_n607), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n268), .A2(new_n273), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n600), .A2(new_n433), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n614), .ZN(G1326gat));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n377), .ZN(new_n616));
  XNOR2_X1  g415(.A(KEYINPUT43), .B(G22gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(G1327gat));
  INV_X1    g417(.A(KEYINPUT45), .ZN(new_n619));
  INV_X1    g418(.A(new_n523), .ZN(new_n620));
  INV_X1    g419(.A(new_n598), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n622), .A2(new_n561), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n495), .A2(new_n623), .ZN(new_n624));
  OR3_X1    g423(.A1(new_n624), .A2(G29gat), .A3(new_n337), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(KEYINPUT100), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n625), .A2(KEYINPUT100), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n619), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n628), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n630), .A2(KEYINPUT45), .A3(new_n626), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n378), .A2(new_n402), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n405), .A2(new_n408), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n561), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n634), .A2(KEYINPUT44), .A3(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT44), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n637), .B1(new_n409), .B2(new_n561), .ZN(new_n638));
  AND2_X1   g437(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n622), .A2(new_n494), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  OAI21_X1  g440(.A(G29gat), .B1(new_n641), .B2(new_n337), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n629), .A2(new_n631), .A3(new_n642), .ZN(G1328gat));
  NOR3_X1   g442(.A1(new_n624), .A2(G36gat), .A3(new_n360), .ZN(new_n644));
  XNOR2_X1  g443(.A(KEYINPUT101), .B(KEYINPUT46), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(G36gat), .B1(new_n641), .B2(new_n360), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(G1329gat));
  INV_X1    g447(.A(new_n613), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n412), .B1(new_n624), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n276), .A2(G43gat), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n650), .B1(new_n641), .B2(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g452(.A1(new_n377), .A2(new_n410), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT102), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n495), .A2(new_n623), .A3(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n641), .A2(new_n376), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n656), .B1(new_n657), .B2(new_n410), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT48), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  OAI211_X1 g459(.A(KEYINPUT48), .B(new_n656), .C1(new_n657), .C2(new_n410), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(G1331gat));
  INV_X1    g461(.A(KEYINPUT103), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n562), .A2(new_n621), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n634), .A2(new_n663), .A3(new_n494), .A4(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n494), .ZN(new_n666));
  OAI21_X1  g465(.A(KEYINPUT103), .B1(new_n409), .B2(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n665), .A2(new_n667), .A3(new_n403), .ZN(new_n668));
  XOR2_X1   g467(.A(new_n668), .B(new_n504), .Z(G1332gat));
  AND3_X1   g468(.A1(new_n665), .A2(new_n667), .A3(KEYINPUT104), .ZN(new_n670));
  AOI21_X1  g469(.A(KEYINPUT104), .B1(new_n665), .B2(new_n667), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(new_n604), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n673), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n674));
  XOR2_X1   g473(.A(KEYINPUT49), .B(G64gat), .Z(new_n675));
  OAI21_X1  g474(.A(new_n674), .B1(new_n673), .B2(new_n675), .ZN(G1333gat));
  INV_X1    g475(.A(G71gat), .ZN(new_n677));
  NAND4_X1  g476(.A1(new_n665), .A2(new_n667), .A3(new_n677), .A4(new_n613), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n670), .A2(new_n671), .A3(new_n611), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n678), .B1(new_n679), .B2(new_n677), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT50), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  OAI211_X1 g481(.A(KEYINPUT50), .B(new_n678), .C1(new_n679), .C2(new_n677), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(G1334gat));
  NAND2_X1  g483(.A1(new_n672), .A2(new_n377), .ZN(new_n685));
  XOR2_X1   g484(.A(KEYINPUT105), .B(G78gat), .Z(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(G1335gat));
  NOR2_X1   g486(.A1(new_n523), .A2(new_n493), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n634), .A2(new_n635), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(KEYINPUT51), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT51), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n634), .A2(new_n691), .A3(new_n635), .A4(new_n688), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n690), .A2(new_n598), .A3(new_n692), .ZN(new_n693));
  OR3_X1    g492(.A1(new_n693), .A2(G85gat), .A3(new_n337), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n523), .A2(new_n493), .A3(new_n621), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n639), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(G85gat), .B1(new_n696), .B2(new_n337), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n694), .A2(new_n697), .ZN(G1336gat));
  NAND4_X1  g497(.A1(new_n636), .A2(new_n638), .A3(new_n604), .A4(new_n695), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(G92gat), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n360), .A2(G92gat), .ZN(new_n701));
  NAND4_X1  g500(.A1(new_n690), .A2(new_n598), .A3(new_n692), .A4(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT107), .ZN(new_n703));
  AND3_X1   g502(.A1(new_n700), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n703), .B1(new_n700), .B2(new_n702), .ZN(new_n705));
  AOI21_X1  g504(.A(KEYINPUT106), .B1(new_n699), .B2(G92gat), .ZN(new_n706));
  OAI22_X1  g505(.A1(new_n704), .A2(new_n705), .B1(KEYINPUT52), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n700), .A2(new_n702), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(KEYINPUT107), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n706), .A2(KEYINPUT52), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n700), .A2(new_n702), .A3(new_n703), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  AND2_X1   g511(.A1(new_n707), .A2(new_n712), .ZN(G1337gat));
  OAI21_X1  g512(.A(G99gat), .B1(new_n696), .B2(new_n611), .ZN(new_n714));
  OR2_X1    g513(.A1(new_n649), .A2(G99gat), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n714), .B1(new_n693), .B2(new_n715), .ZN(G1338gat));
  OAI21_X1  g515(.A(G106gat), .B1(new_n696), .B2(new_n376), .ZN(new_n717));
  OR2_X1    g516(.A1(new_n376), .A2(G106gat), .ZN(new_n718));
  OR2_X1    g517(.A1(new_n693), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT108), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n720), .A2(new_n722), .A3(KEYINPUT53), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT53), .ZN(new_n724));
  OAI211_X1 g523(.A(new_n717), .B(new_n719), .C1(new_n721), .C2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n723), .A2(new_n725), .ZN(G1339gat));
  NAND2_X1  g525(.A1(new_n599), .A2(new_n494), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n597), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n584), .A2(new_n586), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n730), .A2(KEYINPUT54), .A3(new_n595), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT54), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n592), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT109), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n734), .A2(new_n735), .A3(new_n567), .ZN(new_n736));
  AOI21_X1  g535(.A(KEYINPUT54), .B1(new_n587), .B2(new_n591), .ZN(new_n737));
  OAI21_X1  g536(.A(KEYINPUT109), .B1(new_n737), .B2(new_n566), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n732), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n729), .B1(new_n739), .B2(KEYINPUT55), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n735), .B1(new_n734), .B2(new_n567), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n737), .A2(KEYINPUT109), .A3(new_n566), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n731), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT55), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n740), .A2(new_n635), .A3(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n492), .ZN(new_n747));
  OAI21_X1  g546(.A(KEYINPUT87), .B1(new_n491), .B2(new_n482), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n453), .B1(new_n451), .B2(new_n455), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n452), .B1(new_n450), .B2(new_n467), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n477), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  XOR2_X1   g551(.A(new_n752), .B(KEYINPUT110), .Z(new_n753));
  NAND2_X1  g552(.A1(new_n749), .A2(new_n753), .ZN(new_n754));
  OR2_X1    g553(.A1(new_n746), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n740), .A2(new_n493), .A3(new_n745), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n749), .A2(new_n753), .A3(new_n598), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n755), .B1(new_n758), .B2(new_n635), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n728), .B1(new_n759), .B2(new_n620), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n760), .A2(new_n337), .A3(new_n404), .ZN(new_n761));
  INV_X1    g560(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n762), .A2(new_n494), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n763), .A2(G113gat), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n764), .B1(new_n763), .B2(new_n234), .ZN(G1340gat));
  OAI21_X1  g564(.A(G120gat), .B1(new_n762), .B2(new_n621), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n598), .A2(new_n232), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(KEYINPUT111), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n766), .B1(new_n762), .B2(new_n768), .ZN(G1341gat));
  NAND2_X1  g568(.A1(new_n761), .A2(new_n523), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(G127gat), .ZN(G1342gat));
  INV_X1    g570(.A(new_n760), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n649), .A2(new_n377), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n774), .A2(G134gat), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n604), .A2(new_n561), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n772), .A2(new_n775), .A3(new_n403), .A4(new_n776), .ZN(new_n777));
  XOR2_X1   g576(.A(new_n777), .B(KEYINPUT56), .Z(new_n778));
  OAI21_X1  g577(.A(G134gat), .B1(new_n762), .B2(new_n561), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(G1343gat));
  NOR3_X1   g579(.A1(new_n276), .A2(new_n337), .A3(new_n604), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n760), .A2(new_n376), .ZN(new_n782));
  OAI211_X1 g581(.A(KEYINPUT55), .B(new_n731), .C1(new_n741), .C2(new_n742), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n783), .A2(new_n493), .A3(new_n597), .ZN(new_n784));
  XNOR2_X1  g583(.A(KEYINPUT112), .B(KEYINPUT55), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n739), .A2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n757), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(new_n561), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n523), .B1(new_n755), .B2(new_n788), .ZN(new_n789));
  OAI211_X1 g588(.A(KEYINPUT57), .B(new_n377), .C1(new_n789), .C2(new_n728), .ZN(new_n790));
  OAI22_X1  g589(.A1(new_n782), .A2(KEYINPUT57), .B1(KEYINPUT113), .B2(new_n790), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n790), .A2(KEYINPUT113), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n781), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OR2_X1    g592(.A1(new_n793), .A2(new_n494), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(G141gat), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT58), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT115), .ZN(new_n797));
  NOR4_X1   g596(.A1(new_n760), .A2(new_n337), .A3(new_n376), .A4(new_n276), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n360), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n494), .A2(G141gat), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n797), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n799), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n803), .A2(KEYINPUT115), .A3(new_n800), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n795), .A2(new_n796), .A3(new_n802), .A4(new_n804), .ZN(new_n805));
  OR3_X1    g604(.A1(new_n799), .A2(KEYINPUT114), .A3(new_n801), .ZN(new_n806));
  OAI21_X1  g605(.A(KEYINPUT114), .B1(new_n799), .B2(new_n801), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n808), .B1(G141gat), .B2(new_n794), .ZN(new_n809));
  OAI211_X1 g608(.A(new_n805), .B(KEYINPUT116), .C1(new_n809), .C2(new_n796), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT116), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n806), .A2(new_n807), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n796), .B1(new_n795), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n804), .A2(new_n796), .A3(new_n802), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n814), .B1(G141gat), .B2(new_n794), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n811), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n810), .A2(new_n816), .ZN(G1344gat));
  INV_X1    g616(.A(KEYINPUT59), .ZN(new_n818));
  OAI211_X1 g617(.A(new_n818), .B(G148gat), .C1(new_n793), .C2(new_n621), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT57), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n760), .A2(new_n820), .A3(new_n376), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT119), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT118), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n754), .B1(new_n746), .B2(new_n823), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n740), .A2(new_n745), .A3(KEYINPUT118), .A4(new_n635), .ZN(new_n825));
  AOI22_X1  g624(.A1(new_n824), .A2(new_n825), .B1(new_n561), .B2(new_n787), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n822), .B(new_n727), .C1(new_n826), .C2(new_n523), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n635), .B1(new_n739), .B2(KEYINPUT55), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n783), .A2(new_n597), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n823), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(new_n754), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n830), .A2(new_n831), .A3(new_n825), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n523), .B1(new_n832), .B2(new_n788), .ZN(new_n833));
  OAI21_X1  g632(.A(KEYINPUT119), .B1(new_n833), .B2(new_n728), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n827), .A2(new_n834), .A3(new_n377), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n820), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT120), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n821), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n835), .A2(KEYINPUT120), .A3(new_n820), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT117), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n598), .B1(new_n781), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n842), .B1(new_n841), .B2(new_n781), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n291), .B1(new_n840), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n819), .B1(new_n844), .B2(new_n818), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n803), .A2(new_n291), .A3(new_n598), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(G1345gat));
  OAI21_X1  g646(.A(G155gat), .B1(new_n793), .B2(new_n620), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n803), .A2(new_n285), .A3(new_n523), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(G1346gat));
  OAI21_X1  g649(.A(G162gat), .B1(new_n793), .B2(new_n561), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n798), .A2(new_n286), .A3(new_n776), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(G1347gat));
  NOR3_X1   g652(.A1(new_n774), .A2(new_n403), .A3(new_n360), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(new_n772), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n855), .A2(new_n494), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n856), .B(new_n209), .ZN(G1348gat));
  NOR2_X1   g656(.A1(new_n855), .A2(new_n621), .ZN(new_n858));
  XNOR2_X1  g657(.A(KEYINPUT121), .B(G176gat), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n858), .B(new_n859), .ZN(G1349gat));
  NOR2_X1   g659(.A1(new_n855), .A2(new_n620), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n861), .A2(new_n205), .ZN(new_n862));
  AOI211_X1 g661(.A(KEYINPUT122), .B(new_n862), .C1(new_n239), .C2(new_n861), .ZN(new_n863));
  XOR2_X1   g662(.A(new_n863), .B(KEYINPUT60), .Z(G1350gat));
  NAND3_X1  g663(.A1(new_n854), .A2(new_n772), .A3(new_n635), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n865), .A2(G190gat), .ZN(new_n866));
  XNOR2_X1  g665(.A(new_n866), .B(KEYINPUT123), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(G190gat), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n868), .B(KEYINPUT61), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n867), .A2(new_n869), .ZN(G1351gat));
  INV_X1    g669(.A(new_n782), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n276), .A2(new_n403), .A3(new_n360), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(G197gat), .B1(new_n874), .B2(new_n493), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n840), .B(KEYINPUT124), .ZN(new_n876));
  AND3_X1   g675(.A1(new_n872), .A2(G197gat), .A3(new_n493), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(G1352gat));
  NAND2_X1  g677(.A1(new_n876), .A2(new_n872), .ZN(new_n879));
  OAI21_X1  g678(.A(G204gat), .B1(new_n879), .B2(new_n621), .ZN(new_n880));
  NOR4_X1   g679(.A1(new_n871), .A2(new_n873), .A3(G204gat), .A4(new_n621), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(KEYINPUT62), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(new_n882), .ZN(G1353gat));
  INV_X1    g682(.A(KEYINPUT63), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n872), .A2(new_n523), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n885), .B1(new_n838), .B2(new_n839), .ZN(new_n886));
  INV_X1    g685(.A(G211gat), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n884), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AND3_X1   g687(.A1(new_n835), .A2(KEYINPUT120), .A3(new_n820), .ZN(new_n889));
  AOI21_X1  g688(.A(KEYINPUT120), .B1(new_n835), .B2(new_n820), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n889), .A2(new_n890), .A3(new_n821), .ZN(new_n891));
  OAI211_X1 g690(.A(KEYINPUT63), .B(G211gat), .C1(new_n891), .C2(new_n885), .ZN(new_n892));
  AND3_X1   g691(.A1(new_n888), .A2(KEYINPUT125), .A3(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT125), .ZN(new_n894));
  OAI211_X1 g693(.A(new_n894), .B(new_n884), .C1(new_n886), .C2(new_n887), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n782), .A2(new_n887), .A3(new_n523), .A4(new_n872), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(KEYINPUT126), .B1(new_n893), .B2(new_n897), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n888), .A2(new_n892), .A3(KEYINPUT125), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT126), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n899), .A2(new_n900), .A3(new_n895), .A4(new_n896), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n898), .A2(new_n901), .ZN(G1354gat));
  AOI21_X1  g701(.A(G218gat), .B1(new_n874), .B2(new_n635), .ZN(new_n903));
  INV_X1    g702(.A(new_n879), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n635), .A2(G218gat), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(KEYINPUT127), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n903), .B1(new_n904), .B2(new_n906), .ZN(G1355gat));
endmodule


