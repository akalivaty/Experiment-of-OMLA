

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762;

  AND2_X1 U374 ( .A1(n388), .A2(n390), .ZN(n352) );
  INV_X1 U375 ( .A(n641), .ZN(n400) );
  XNOR2_X1 U376 ( .A(n749), .B(n436), .ZN(n504) );
  INV_X1 U377 ( .A(G953), .ZN(n580) );
  NOR2_X1 U378 ( .A1(G953), .A2(G237), .ZN(n523) );
  NAND2_X1 U379 ( .A1(n352), .A2(n386), .ZN(G75) );
  NAND2_X1 U380 ( .A1(n391), .A2(n380), .ZN(n389) );
  NAND2_X1 U381 ( .A1(n658), .A2(n404), .ZN(n391) );
  XNOR2_X2 U382 ( .A(n431), .B(n430), .ZN(n761) );
  NOR2_X1 U383 ( .A1(n693), .A2(n691), .ZN(n633) );
  XNOR2_X1 U384 ( .A(n441), .B(n512), .ZN(n733) );
  INV_X1 U385 ( .A(G146), .ZN(n436) );
  AND2_X2 U386 ( .A1(n395), .A2(n418), .ZN(n394) );
  INV_X2 U387 ( .A(n426), .ZN(n513) );
  XNOR2_X1 U388 ( .A(n442), .B(KEYINPUT48), .ZN(n396) );
  XNOR2_X1 U389 ( .A(n467), .B(KEYINPUT0), .ZN(n607) );
  INV_X1 U390 ( .A(n638), .ZN(n466) );
  XNOR2_X1 U391 ( .A(KEYINPUT38), .B(n578), .ZN(n628) );
  BUF_X1 U392 ( .A(n559), .Z(n647) );
  XNOR2_X1 U393 ( .A(n504), .B(n353), .ZN(n668) );
  XNOR2_X2 U394 ( .A(G137), .B(G128), .ZN(n472) );
  INV_X2 U395 ( .A(G128), .ZN(n398) );
  NOR2_X1 U396 ( .A1(n547), .A2(n507), .ZN(n508) );
  XNOR2_X2 U397 ( .A(KEYINPUT3), .B(G119), .ZN(n500) );
  XOR2_X2 U398 ( .A(G101), .B(G113), .Z(n501) );
  XNOR2_X1 U399 ( .A(n397), .B(n489), .ZN(n749) );
  XNOR2_X1 U400 ( .A(G137), .B(G134), .ZN(n489) );
  XOR2_X1 U401 ( .A(G131), .B(G140), .Z(n529) );
  XNOR2_X1 U402 ( .A(KEYINPUT70), .B(G110), .ZN(n518) );
  XNOR2_X1 U403 ( .A(n586), .B(n585), .ZN(n637) );
  XNOR2_X1 U404 ( .A(n511), .B(KEYINPUT16), .ZN(n441) );
  NOR2_X1 U405 ( .A1(n637), .A2(n612), .ZN(n371) );
  XNOR2_X1 U406 ( .A(n545), .B(G478), .ZN(n557) );
  XNOR2_X1 U407 ( .A(n399), .B(KEYINPUT88), .ZN(n599) );
  XNOR2_X1 U408 ( .A(n366), .B(n365), .ZN(n364) );
  INV_X1 U409 ( .A(KEYINPUT114), .ZN(n365) );
  NOR2_X1 U410 ( .A1(n651), .A2(n652), .ZN(n366) );
  XNOR2_X1 U411 ( .A(KEYINPUT5), .B(KEYINPUT96), .ZN(n454) );
  XNOR2_X1 U412 ( .A(G116), .B(G131), .ZN(n502) );
  XNOR2_X1 U413 ( .A(n456), .B(KEYINPUT95), .ZN(n455) );
  AND2_X1 U414 ( .A1(n419), .A2(n700), .ZN(n418) );
  NAND2_X1 U415 ( .A1(n421), .A2(n420), .ZN(n419) );
  INV_X1 U416 ( .A(n701), .ZN(n421) );
  INV_X1 U417 ( .A(n396), .ZN(n393) );
  XNOR2_X1 U418 ( .A(n375), .B(n437), .ZN(n374) );
  INV_X1 U419 ( .A(KEYINPUT87), .ZN(n437) );
  XNOR2_X1 U420 ( .A(KEYINPUT4), .B(KEYINPUT67), .ZN(n468) );
  XNOR2_X1 U421 ( .A(n518), .B(KEYINPUT18), .ZN(n440) );
  XNOR2_X1 U422 ( .A(n564), .B(KEYINPUT19), .ZN(n373) );
  INV_X1 U423 ( .A(G472), .ZN(n452) );
  INV_X1 U424 ( .A(KEYINPUT66), .ZN(n405) );
  XNOR2_X1 U425 ( .A(n478), .B(n477), .ZN(n539) );
  XOR2_X1 U426 ( .A(KEYINPUT68), .B(KEYINPUT8), .Z(n478) );
  XOR2_X1 U427 ( .A(KEYINPUT7), .B(KEYINPUT100), .Z(n536) );
  XNOR2_X1 U428 ( .A(G134), .B(KEYINPUT9), .ZN(n535) );
  XNOR2_X1 U429 ( .A(G122), .B(KEYINPUT98), .ZN(n534) );
  XNOR2_X1 U430 ( .A(n522), .B(n459), .ZN(n527) );
  AND2_X1 U431 ( .A1(n368), .A2(n656), .ZN(n657) );
  NOR2_X1 U432 ( .A1(n654), .A2(n655), .ZN(n369) );
  INV_X1 U433 ( .A(KEYINPUT28), .ZN(n449) );
  NAND2_X1 U434 ( .A1(n554), .A2(n627), .ZN(n564) );
  AND2_X1 U435 ( .A1(n609), .A2(n466), .ZN(n465) );
  OR2_X1 U436 ( .A1(n641), .A2(n598), .ZN(n412) );
  XNOR2_X1 U437 ( .A(n462), .B(n461), .ZN(n561) );
  INV_X1 U438 ( .A(KEYINPUT101), .ZN(n461) );
  XNOR2_X1 U439 ( .A(n607), .B(n372), .ZN(n612) );
  NOR2_X1 U440 ( .A1(n607), .A2(n594), .ZN(n595) );
  BUF_X1 U441 ( .A(n515), .Z(n751) );
  XNOR2_X1 U442 ( .A(n408), .B(n493), .ZN(n495) );
  XNOR2_X1 U443 ( .A(n492), .B(n494), .ZN(n408) );
  XNOR2_X1 U444 ( .A(n706), .B(n705), .ZN(n707) );
  NOR2_X1 U445 ( .A1(n751), .A2(G952), .ZN(n732) );
  XNOR2_X1 U446 ( .A(n428), .B(n427), .ZN(n572) );
  INV_X1 U447 ( .A(KEYINPUT78), .ZN(n427) );
  INV_X1 U448 ( .A(KEYINPUT85), .ZN(n420) );
  XNOR2_X1 U449 ( .A(n483), .B(n482), .ZN(n484) );
  INV_X1 U450 ( .A(KEYINPUT25), .ZN(n482) );
  AND2_X1 U451 ( .A1(n619), .A2(n377), .ZN(n376) );
  XOR2_X1 U452 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n525) );
  XNOR2_X1 U453 ( .A(n460), .B(G104), .ZN(n522) );
  INV_X1 U454 ( .A(G122), .ZN(n460) );
  XNOR2_X1 U455 ( .A(G113), .B(G143), .ZN(n459) );
  XOR2_X1 U456 ( .A(G902), .B(KEYINPUT15), .Z(n662) );
  XNOR2_X1 U457 ( .A(n363), .B(n362), .ZN(n653) );
  INV_X1 U458 ( .A(KEYINPUT52), .ZN(n362) );
  NAND2_X1 U459 ( .A1(n400), .A2(n434), .ZN(n608) );
  OR2_X1 U460 ( .A1(G902), .A2(G237), .ZN(n519) );
  INV_X1 U461 ( .A(n662), .ZN(n664) );
  INV_X1 U462 ( .A(n647), .ZN(n609) );
  INV_X1 U463 ( .A(G469), .ZN(n422) );
  OR2_X1 U464 ( .A1(n713), .A2(G902), .ZN(n423) );
  XOR2_X1 U465 ( .A(n559), .B(KEYINPUT6), .Z(n590) );
  INV_X1 U466 ( .A(n606), .ZN(n638) );
  XNOR2_X1 U467 ( .A(KEYINPUT94), .B(KEYINPUT21), .ZN(n407) );
  XNOR2_X1 U468 ( .A(n455), .B(n453), .ZN(n503) );
  XNOR2_X1 U469 ( .A(n502), .B(n454), .ZN(n453) );
  NAND2_X1 U470 ( .A1(n393), .A2(n355), .ZN(n392) );
  XNOR2_X1 U471 ( .A(G119), .B(G110), .ZN(n473) );
  XNOR2_X1 U472 ( .A(n417), .B(n416), .ZN(n433) );
  XNOR2_X1 U473 ( .A(KEYINPUT81), .B(KEYINPUT23), .ZN(n417) );
  XNOR2_X1 U474 ( .A(G140), .B(KEYINPUT24), .ZN(n416) );
  XNOR2_X1 U475 ( .A(n491), .B(n490), .ZN(n492) );
  INV_X1 U476 ( .A(n529), .ZN(n490) );
  XNOR2_X1 U477 ( .A(G101), .B(G107), .ZN(n494) );
  XNOR2_X1 U478 ( .A(n733), .B(n379), .ZN(n704) );
  XNOR2_X1 U479 ( .A(n440), .B(n516), .ZN(n439) );
  NAND2_X1 U480 ( .A1(n367), .A2(KEYINPUT118), .ZN(n403) );
  INV_X1 U481 ( .A(n657), .ZN(n367) );
  INV_X1 U482 ( .A(n555), .ZN(n429) );
  XNOR2_X1 U483 ( .A(n532), .B(n432), .ZN(n558) );
  XNOR2_X1 U484 ( .A(n531), .B(n463), .ZN(n432) );
  INV_X1 U485 ( .A(G475), .ZN(n463) );
  XNOR2_X1 U486 ( .A(n541), .B(n425), .ZN(n726) );
  XNOR2_X1 U487 ( .A(n540), .B(n544), .ZN(n425) );
  XNOR2_X1 U488 ( .A(n718), .B(n717), .ZN(n719) );
  NAND2_X1 U489 ( .A1(n385), .A2(KEYINPUT118), .ZN(n381) );
  XNOR2_X1 U490 ( .A(KEYINPUT42), .B(n551), .ZN(n762) );
  INV_X1 U491 ( .A(KEYINPUT40), .ZN(n430) );
  XNOR2_X1 U492 ( .A(n371), .B(n587), .ZN(n370) );
  AND2_X1 U493 ( .A1(n588), .A2(n554), .ZN(n446) );
  NAND2_X2 U494 ( .A1(n411), .A2(n409), .ZN(n684) );
  NAND2_X1 U495 ( .A1(n410), .A2(KEYINPUT102), .ZN(n409) );
  AND2_X1 U496 ( .A1(n413), .A2(n359), .ZN(n411) );
  INV_X1 U497 ( .A(n561), .ZN(n691) );
  XNOR2_X1 U498 ( .A(n713), .B(n712), .ZN(n714) );
  NOR2_X1 U499 ( .A1(n732), .A2(n709), .ZN(n711) );
  XOR2_X1 U500 ( .A(n511), .B(n503), .Z(n353) );
  XNOR2_X1 U501 ( .A(n487), .B(n407), .ZN(n593) );
  OR2_X1 U502 ( .A1(n637), .A2(n636), .ZN(n354) );
  AND2_X1 U503 ( .A1(n701), .A2(KEYINPUT85), .ZN(n355) );
  AND2_X1 U504 ( .A1(n698), .A2(n571), .ZN(n356) );
  XOR2_X1 U505 ( .A(n520), .B(KEYINPUT76), .Z(n357) );
  AND2_X1 U506 ( .A1(n583), .A2(n626), .ZN(n358) );
  AND2_X1 U507 ( .A1(n465), .A2(n412), .ZN(n359) );
  AND2_X1 U508 ( .A1(n633), .A2(KEYINPUT47), .ZN(n360) );
  XOR2_X1 U509 ( .A(KEYINPUT1), .B(KEYINPUT65), .Z(n361) );
  NAND2_X1 U510 ( .A1(n364), .A2(n354), .ZN(n363) );
  XNOR2_X1 U511 ( .A(n369), .B(KEYINPUT117), .ZN(n368) );
  NAND2_X1 U512 ( .A1(n370), .A2(n588), .ZN(n589) );
  INV_X1 U513 ( .A(KEYINPUT93), .ZN(n372) );
  NAND2_X1 U514 ( .A1(n373), .A2(n358), .ZN(n467) );
  NAND2_X1 U515 ( .A1(n429), .A2(n373), .ZN(n568) );
  AND2_X1 U516 ( .A1(n376), .A2(n374), .ZN(n435) );
  NAND2_X1 U517 ( .A1(n758), .A2(KEYINPUT44), .ZN(n375) );
  NAND2_X1 U518 ( .A1(n599), .A2(KEYINPUT44), .ZN(n377) );
  XNOR2_X2 U519 ( .A(n378), .B(n357), .ZN(n554) );
  NAND2_X1 U520 ( .A1(n704), .A2(n664), .ZN(n378) );
  XNOR2_X1 U521 ( .A(n438), .B(n439), .ZN(n379) );
  INV_X1 U522 ( .A(n402), .ZN(n380) );
  NAND2_X1 U523 ( .A1(n382), .A2(n381), .ZN(n386) );
  INV_X1 U524 ( .A(n658), .ZN(n385) );
  AND2_X1 U525 ( .A1(n383), .A2(n391), .ZN(n382) );
  NOR2_X1 U526 ( .A1(n402), .A2(n661), .ZN(n383) );
  NAND2_X1 U527 ( .A1(n385), .A2(n384), .ZN(n390) );
  AND2_X1 U528 ( .A1(n661), .A2(KEYINPUT118), .ZN(n384) );
  NAND2_X1 U529 ( .A1(n389), .A2(n661), .ZN(n388) );
  NAND2_X2 U530 ( .A1(n394), .A2(n392), .ZN(n750) );
  NAND2_X1 U531 ( .A1(n396), .A2(n420), .ZN(n395) );
  XNOR2_X1 U532 ( .A(n471), .B(n397), .ZN(n438) );
  XNOR2_X2 U533 ( .A(n533), .B(n468), .ZN(n397) );
  XNOR2_X2 U534 ( .A(n398), .B(G143), .ZN(n533) );
  NAND2_X1 U535 ( .A1(n684), .A2(n759), .ZN(n399) );
  NOR2_X1 U536 ( .A1(n608), .A2(n603), .ZN(n586) );
  XNOR2_X2 U537 ( .A(n566), .B(n361), .ZN(n641) );
  NAND2_X1 U538 ( .A1(n401), .A2(n691), .ZN(n431) );
  NAND2_X1 U539 ( .A1(n401), .A2(n693), .ZN(n700) );
  XNOR2_X2 U540 ( .A(n521), .B(KEYINPUT39), .ZN(n401) );
  NAND2_X1 U541 ( .A1(n403), .A2(n580), .ZN(n402) );
  AND2_X1 U542 ( .A1(n657), .A2(n457), .ZN(n404) );
  XNOR2_X2 U543 ( .A(n406), .B(n405), .ZN(n640) );
  NOR2_X2 U544 ( .A1(n606), .A2(n593), .ZN(n406) );
  XNOR2_X2 U545 ( .A(n485), .B(n484), .ZN(n606) );
  INV_X1 U546 ( .A(n472), .ZN(n474) );
  INV_X1 U547 ( .A(n518), .ZN(n517) );
  NOR2_X2 U548 ( .A1(G902), .A2(n668), .ZN(n505) );
  AND2_X1 U549 ( .A1(n597), .A2(n641), .ZN(n604) );
  INV_X1 U550 ( .A(n597), .ZN(n410) );
  NAND2_X1 U551 ( .A1(n597), .A2(n414), .ZN(n413) );
  AND2_X1 U552 ( .A1(n641), .A2(n598), .ZN(n414) );
  XNOR2_X2 U553 ( .A(n415), .B(KEYINPUT32), .ZN(n759) );
  NAND2_X1 U554 ( .A1(n597), .A2(n596), .ZN(n415) );
  INV_X1 U555 ( .A(n554), .ZN(n578) );
  NOR2_X2 U556 ( .A1(n640), .A2(n566), .ZN(n614) );
  XNOR2_X2 U557 ( .A(n423), .B(n422), .ZN(n566) );
  XNOR2_X1 U558 ( .A(n495), .B(n504), .ZN(n713) );
  NAND2_X2 U559 ( .A1(n424), .A2(n628), .ZN(n521) );
  AND2_X1 U560 ( .A1(n424), .A2(n446), .ZN(n689) );
  XNOR2_X2 U561 ( .A(n510), .B(KEYINPUT73), .ZN(n424) );
  XNOR2_X1 U562 ( .A(n533), .B(n534), .ZN(n538) );
  NAND2_X1 U563 ( .A1(n558), .A2(n557), .ZN(n462) );
  XNOR2_X2 U564 ( .A(G125), .B(G146), .ZN(n426) );
  NAND2_X1 U565 ( .A1(n445), .A2(n447), .ZN(n428) );
  INV_X1 U566 ( .A(n568), .ZN(n686) );
  INV_X1 U567 ( .A(n560), .ZN(n451) );
  NAND2_X1 U568 ( .A1(n523), .A2(G210), .ZN(n456) );
  NOR2_X2 U569 ( .A1(n761), .A2(n762), .ZN(n552) );
  XNOR2_X1 U570 ( .A(n475), .B(n433), .ZN(n476) );
  XNOR2_X1 U571 ( .A(n602), .B(KEYINPUT72), .ZN(n470) );
  NOR2_X1 U572 ( .A1(n689), .A2(n360), .ZN(n445) );
  INV_X1 U573 ( .A(n640), .ZN(n434) );
  NAND2_X1 U574 ( .A1(n435), .A2(n470), .ZN(n469) );
  XNOR2_X2 U575 ( .A(n589), .B(KEYINPUT35), .ZN(n758) );
  NAND2_X1 U576 ( .A1(n444), .A2(n443), .ZN(n442) );
  XNOR2_X1 U577 ( .A(n458), .B(KEYINPUT69), .ZN(n443) );
  XNOR2_X1 U578 ( .A(n552), .B(KEYINPUT46), .ZN(n444) );
  XNOR2_X1 U579 ( .A(n556), .B(n448), .ZN(n447) );
  INV_X1 U580 ( .A(KEYINPUT79), .ZN(n448) );
  XNOR2_X1 U581 ( .A(n450), .B(n449), .ZN(n550) );
  NAND2_X1 U582 ( .A1(n647), .A2(n451), .ZN(n450) );
  XNOR2_X2 U583 ( .A(n505), .B(n452), .ZN(n559) );
  INV_X1 U584 ( .A(KEYINPUT118), .ZN(n457) );
  NAND2_X1 U585 ( .A1(n356), .A2(n572), .ZN(n458) );
  AND2_X4 U586 ( .A1(n464), .A2(n702), .ZN(n724) );
  NAND2_X1 U587 ( .A1(n703), .A2(n464), .ZN(n708) );
  NAND2_X2 U588 ( .A1(n667), .A2(n666), .ZN(n464) );
  XNOR2_X2 U589 ( .A(n469), .B(n620), .ZN(n741) );
  XNOR2_X1 U590 ( .A(n708), .B(n707), .ZN(n709) );
  NAND2_X1 U591 ( .A1(n750), .A2(n621), .ZN(n579) );
  NOR2_X2 U592 ( .A1(n721), .A2(n732), .ZN(n723) );
  NOR2_X2 U593 ( .A1(n671), .A2(n732), .ZN(n674) );
  XNOR2_X2 U594 ( .A(n501), .B(n500), .ZN(n511) );
  AND2_X1 U595 ( .A1(G224), .A2(n515), .ZN(n471) );
  XNOR2_X1 U596 ( .A(n584), .B(KEYINPUT103), .ZN(n585) );
  INV_X1 U597 ( .A(KEYINPUT99), .ZN(n542) );
  INV_X1 U598 ( .A(KEYINPUT102), .ZN(n598) );
  XNOR2_X1 U599 ( .A(n720), .B(n719), .ZN(n721) );
  XNOR2_X1 U600 ( .A(n672), .B(KEYINPUT63), .ZN(n673) );
  XNOR2_X1 U601 ( .A(n715), .B(n714), .ZN(n716) );
  XNOR2_X1 U602 ( .A(n474), .B(n473), .ZN(n475) );
  XOR2_X1 U603 ( .A(KEYINPUT10), .B(n513), .Z(n528) );
  XNOR2_X1 U604 ( .A(n476), .B(n528), .ZN(n480) );
  XOR2_X2 U605 ( .A(G953), .B(KEYINPUT64), .Z(n515) );
  NAND2_X1 U606 ( .A1(G234), .A2(n515), .ZN(n477) );
  NAND2_X1 U607 ( .A1(G221), .A2(n539), .ZN(n479) );
  XNOR2_X1 U608 ( .A(n480), .B(n479), .ZN(n728) );
  NOR2_X1 U609 ( .A1(n728), .A2(G902), .ZN(n485) );
  NAND2_X1 U610 ( .A1(G234), .A2(n664), .ZN(n481) );
  XNOR2_X1 U611 ( .A(KEYINPUT20), .B(n481), .ZN(n486) );
  NAND2_X1 U612 ( .A1(G217), .A2(n486), .ZN(n483) );
  NAND2_X1 U613 ( .A1(n486), .A2(G221), .ZN(n487) );
  INV_X1 U614 ( .A(n593), .ZN(n488) );
  XOR2_X1 U615 ( .A(G104), .B(n517), .Z(n493) );
  NAND2_X1 U616 ( .A1(G227), .A2(n515), .ZN(n491) );
  XNOR2_X1 U617 ( .A(n614), .B(KEYINPUT106), .ZN(n509) );
  NAND2_X1 U618 ( .A1(G234), .A2(G237), .ZN(n496) );
  XNOR2_X1 U619 ( .A(n496), .B(KEYINPUT14), .ZN(n626) );
  NOR2_X1 U620 ( .A1(n751), .A2(G900), .ZN(n497) );
  NAND2_X1 U621 ( .A1(G902), .A2(n497), .ZN(n498) );
  NAND2_X1 U622 ( .A1(G952), .A2(n580), .ZN(n581) );
  NAND2_X1 U623 ( .A1(n498), .A2(n581), .ZN(n499) );
  NAND2_X1 U624 ( .A1(n626), .A2(n499), .ZN(n547) );
  NAND2_X1 U625 ( .A1(G214), .A2(n519), .ZN(n627) );
  NAND2_X1 U626 ( .A1(n559), .A2(n627), .ZN(n506) );
  XNOR2_X1 U627 ( .A(KEYINPUT30), .B(n506), .ZN(n507) );
  NAND2_X1 U628 ( .A1(n509), .A2(n508), .ZN(n510) );
  XOR2_X1 U629 ( .A(G116), .B(G107), .Z(n543) );
  XOR2_X1 U630 ( .A(n522), .B(n543), .Z(n512) );
  XNOR2_X1 U631 ( .A(KEYINPUT17), .B(KEYINPUT91), .ZN(n514) );
  XNOR2_X1 U632 ( .A(n514), .B(n513), .ZN(n516) );
  NAND2_X1 U633 ( .A1(n519), .A2(G210), .ZN(n520) );
  NAND2_X1 U634 ( .A1(n523), .A2(G214), .ZN(n524) );
  XNOR2_X1 U635 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U636 ( .A(n527), .B(n526), .ZN(n530) );
  XNOR2_X1 U637 ( .A(n529), .B(n528), .ZN(n748) );
  XNOR2_X1 U638 ( .A(n530), .B(n748), .ZN(n718) );
  NOR2_X1 U639 ( .A1(G902), .A2(n718), .ZN(n532) );
  XNOR2_X1 U640 ( .A(KEYINPUT97), .B(KEYINPUT13), .ZN(n531) );
  XNOR2_X1 U641 ( .A(n536), .B(n535), .ZN(n537) );
  XOR2_X1 U642 ( .A(n538), .B(n537), .Z(n541) );
  NAND2_X1 U643 ( .A1(G217), .A2(n539), .ZN(n540) );
  XNOR2_X1 U644 ( .A(n543), .B(n542), .ZN(n544) );
  NOR2_X1 U645 ( .A1(n726), .A2(G902), .ZN(n545) );
  INV_X1 U646 ( .A(n558), .ZN(n553) );
  NAND2_X1 U647 ( .A1(n557), .A2(n553), .ZN(n630) );
  NAND2_X1 U648 ( .A1(n628), .A2(n627), .ZN(n632) );
  NOR2_X1 U649 ( .A1(n630), .A2(n632), .ZN(n546) );
  XNOR2_X1 U650 ( .A(n546), .B(KEYINPUT41), .ZN(n652) );
  NOR2_X1 U651 ( .A1(n547), .A2(n593), .ZN(n548) );
  NAND2_X1 U652 ( .A1(n466), .A2(n548), .ZN(n560) );
  INV_X1 U653 ( .A(n566), .ZN(n549) );
  NAND2_X1 U654 ( .A1(n550), .A2(n549), .ZN(n555) );
  NOR2_X1 U655 ( .A1(n652), .A2(n555), .ZN(n551) );
  NOR2_X1 U656 ( .A1(n557), .A2(n553), .ZN(n588) );
  NAND2_X1 U657 ( .A1(n568), .A2(KEYINPUT47), .ZN(n556) );
  NOR2_X1 U658 ( .A1(n558), .A2(n557), .ZN(n693) );
  NOR2_X1 U659 ( .A1(n561), .A2(n560), .ZN(n562) );
  NAND2_X1 U660 ( .A1(n590), .A2(n562), .ZN(n563) );
  XNOR2_X1 U661 ( .A(KEYINPUT104), .B(n563), .ZN(n574) );
  NOR2_X1 U662 ( .A1(n574), .A2(n564), .ZN(n565) );
  XNOR2_X1 U663 ( .A(n565), .B(KEYINPUT36), .ZN(n567) );
  NAND2_X1 U664 ( .A1(n567), .A2(n400), .ZN(n698) );
  XNOR2_X1 U665 ( .A(KEYINPUT80), .B(n633), .ZN(n617) );
  INV_X1 U666 ( .A(n617), .ZN(n570) );
  NOR2_X1 U667 ( .A1(KEYINPUT47), .A2(n568), .ZN(n569) );
  NAND2_X1 U668 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U669 ( .A(KEYINPUT105), .B(KEYINPUT43), .ZN(n576) );
  NAND2_X1 U670 ( .A1(n641), .A2(n627), .ZN(n573) );
  NOR2_X1 U671 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U672 ( .A(n576), .B(n575), .ZN(n577) );
  NAND2_X1 U673 ( .A1(n578), .A2(n577), .ZN(n701) );
  INV_X1 U674 ( .A(KEYINPUT2), .ZN(n621) );
  XNOR2_X1 U675 ( .A(n579), .B(KEYINPUT82), .ZN(n623) );
  XNOR2_X1 U676 ( .A(KEYINPUT92), .B(G898), .ZN(n738) );
  NOR2_X1 U677 ( .A1(n580), .A2(n738), .ZN(n735) );
  NAND2_X1 U678 ( .A1(n735), .A2(G902), .ZN(n582) );
  NAND2_X1 U679 ( .A1(n582), .A2(n581), .ZN(n583) );
  INV_X1 U680 ( .A(n590), .ZN(n603) );
  XNOR2_X1 U681 ( .A(KEYINPUT33), .B(KEYINPUT71), .ZN(n584) );
  XNOR2_X1 U682 ( .A(KEYINPUT34), .B(KEYINPUT74), .ZN(n587) );
  NOR2_X1 U683 ( .A1(n641), .A2(n590), .ZN(n591) );
  NAND2_X1 U684 ( .A1(n466), .A2(n591), .ZN(n592) );
  XNOR2_X1 U685 ( .A(n592), .B(KEYINPUT75), .ZN(n596) );
  OR2_X1 U686 ( .A1(n630), .A2(n593), .ZN(n594) );
  XNOR2_X2 U687 ( .A(n595), .B(KEYINPUT22), .ZN(n597) );
  INV_X1 U688 ( .A(n599), .ZN(n601) );
  NOR2_X1 U689 ( .A1(n758), .A2(KEYINPUT44), .ZN(n600) );
  NAND2_X1 U690 ( .A1(n601), .A2(n600), .ZN(n602) );
  NAND2_X1 U691 ( .A1(n604), .A2(n603), .ZN(n605) );
  NOR2_X1 U692 ( .A1(n466), .A2(n605), .ZN(n675) );
  INV_X1 U693 ( .A(n607), .ZN(n610) );
  NOR2_X1 U694 ( .A1(n609), .A2(n608), .ZN(n649) );
  NAND2_X1 U695 ( .A1(n610), .A2(n649), .ZN(n611) );
  XNOR2_X1 U696 ( .A(n611), .B(KEYINPUT31), .ZN(n694) );
  INV_X1 U697 ( .A(n612), .ZN(n613) );
  NAND2_X1 U698 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U699 ( .A1(n647), .A2(n615), .ZN(n681) );
  NOR2_X1 U700 ( .A1(n694), .A2(n681), .ZN(n616) );
  NOR2_X1 U701 ( .A1(n617), .A2(n616), .ZN(n618) );
  NOR2_X1 U702 ( .A1(n675), .A2(n618), .ZN(n619) );
  XOR2_X1 U703 ( .A(KEYINPUT45), .B(KEYINPUT84), .Z(n620) );
  NAND2_X1 U704 ( .A1(n741), .A2(n621), .ZN(n622) );
  NAND2_X1 U705 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U706 ( .A(n624), .B(KEYINPUT77), .ZN(n625) );
  NOR2_X2 U707 ( .A1(n741), .A2(n750), .ZN(n663) );
  NAND2_X1 U708 ( .A1(n663), .A2(KEYINPUT2), .ZN(n702) );
  NAND2_X1 U709 ( .A1(n625), .A2(n702), .ZN(n658) );
  OR2_X1 U710 ( .A1(n652), .A2(n637), .ZN(n656) );
  NAND2_X1 U711 ( .A1(G952), .A2(n626), .ZN(n655) );
  NOR2_X1 U712 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U713 ( .A1(n630), .A2(n629), .ZN(n631) );
  XOR2_X1 U714 ( .A(KEYINPUT115), .B(n631), .Z(n635) );
  NOR2_X1 U715 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U716 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U717 ( .A1(n488), .A2(n638), .ZN(n639) );
  XNOR2_X1 U718 ( .A(KEYINPUT49), .B(n639), .ZN(n645) );
  XOR2_X1 U719 ( .A(KEYINPUT50), .B(KEYINPUT113), .Z(n643) );
  NAND2_X1 U720 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U721 ( .A(n643), .B(n642), .ZN(n644) );
  NAND2_X1 U722 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U723 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U724 ( .A1(n649), .A2(n648), .ZN(n650) );
  XOR2_X1 U725 ( .A(KEYINPUT51), .B(n650), .Z(n651) );
  XNOR2_X1 U726 ( .A(KEYINPUT116), .B(n653), .ZN(n654) );
  INV_X1 U727 ( .A(KEYINPUT119), .ZN(n660) );
  INV_X1 U728 ( .A(KEYINPUT53), .ZN(n659) );
  XNOR2_X1 U729 ( .A(n660), .B(n659), .ZN(n661) );
  NAND2_X1 U730 ( .A1(n663), .A2(n662), .ZN(n667) );
  XNOR2_X1 U731 ( .A(KEYINPUT83), .B(n664), .ZN(n665) );
  NAND2_X1 U732 ( .A1(n665), .A2(KEYINPUT2), .ZN(n666) );
  NAND2_X1 U733 ( .A1(n724), .A2(G472), .ZN(n670) );
  XNOR2_X1 U734 ( .A(n668), .B(KEYINPUT62), .ZN(n669) );
  XNOR2_X1 U735 ( .A(n670), .B(n669), .ZN(n671) );
  XNOR2_X1 U736 ( .A(KEYINPUT89), .B(KEYINPUT90), .ZN(n672) );
  XNOR2_X1 U737 ( .A(n674), .B(n673), .ZN(G57) );
  XNOR2_X1 U738 ( .A(G101), .B(n675), .ZN(n676) );
  XNOR2_X1 U739 ( .A(n676), .B(KEYINPUT107), .ZN(G3) );
  NAND2_X1 U740 ( .A1(n681), .A2(n691), .ZN(n677) );
  XNOR2_X1 U741 ( .A(n677), .B(G104), .ZN(G6) );
  XOR2_X1 U742 ( .A(KEYINPUT27), .B(KEYINPUT109), .Z(n679) );
  XNOR2_X1 U743 ( .A(G107), .B(KEYINPUT26), .ZN(n678) );
  XNOR2_X1 U744 ( .A(n679), .B(n678), .ZN(n680) );
  XOR2_X1 U745 ( .A(KEYINPUT108), .B(n680), .Z(n683) );
  NAND2_X1 U746 ( .A1(n681), .A2(n693), .ZN(n682) );
  XNOR2_X1 U747 ( .A(n683), .B(n682), .ZN(G9) );
  XNOR2_X1 U748 ( .A(G110), .B(KEYINPUT110), .ZN(n685) );
  XNOR2_X1 U749 ( .A(n685), .B(n684), .ZN(G12) );
  XOR2_X1 U750 ( .A(G128), .B(KEYINPUT29), .Z(n688) );
  NAND2_X1 U751 ( .A1(n686), .A2(n693), .ZN(n687) );
  XNOR2_X1 U752 ( .A(n688), .B(n687), .ZN(G30) );
  XOR2_X1 U753 ( .A(n689), .B(G143), .Z(G45) );
  NAND2_X1 U754 ( .A1(n686), .A2(n691), .ZN(n690) );
  XNOR2_X1 U755 ( .A(n690), .B(G146), .ZN(G48) );
  NAND2_X1 U756 ( .A1(n694), .A2(n691), .ZN(n692) );
  XNOR2_X1 U757 ( .A(n692), .B(G113), .ZN(G15) );
  NAND2_X1 U758 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U759 ( .A(n695), .B(G116), .ZN(G18) );
  XOR2_X1 U760 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n697) );
  XNOR2_X1 U761 ( .A(G125), .B(KEYINPUT37), .ZN(n696) );
  XNOR2_X1 U762 ( .A(n697), .B(n696), .ZN(n699) );
  XOR2_X1 U763 ( .A(n699), .B(n698), .Z(G27) );
  XNOR2_X1 U764 ( .A(G134), .B(n700), .ZN(G36) );
  XNOR2_X1 U765 ( .A(G140), .B(n701), .ZN(G42) );
  AND2_X1 U766 ( .A1(n702), .A2(G210), .ZN(n703) );
  INV_X1 U767 ( .A(n704), .ZN(n706) );
  XOR2_X1 U768 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n705) );
  XNOR2_X1 U769 ( .A(KEYINPUT86), .B(KEYINPUT56), .ZN(n710) );
  XNOR2_X1 U770 ( .A(n711), .B(n710), .ZN(G51) );
  NAND2_X1 U771 ( .A1(n724), .A2(G469), .ZN(n715) );
  XOR2_X1 U772 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n712) );
  NOR2_X1 U773 ( .A1(n732), .A2(n716), .ZN(G54) );
  NAND2_X1 U774 ( .A1(n724), .A2(G475), .ZN(n720) );
  XOR2_X1 U775 ( .A(KEYINPUT120), .B(KEYINPUT59), .Z(n717) );
  XOR2_X1 U776 ( .A(KEYINPUT60), .B(KEYINPUT121), .Z(n722) );
  XNOR2_X1 U777 ( .A(n723), .B(n722), .ZN(G60) );
  NAND2_X1 U778 ( .A1(n724), .A2(G478), .ZN(n725) );
  XNOR2_X1 U779 ( .A(n726), .B(n725), .ZN(n727) );
  NOR2_X1 U780 ( .A1(n732), .A2(n727), .ZN(G63) );
  XNOR2_X1 U781 ( .A(n728), .B(KEYINPUT122), .ZN(n730) );
  NAND2_X1 U782 ( .A1(n724), .A2(G217), .ZN(n729) );
  XNOR2_X1 U783 ( .A(n730), .B(n729), .ZN(n731) );
  NOR2_X1 U784 ( .A1(n732), .A2(n731), .ZN(G66) );
  XNOR2_X1 U785 ( .A(KEYINPUT125), .B(KEYINPUT126), .ZN(n747) );
  XNOR2_X1 U786 ( .A(n733), .B(G110), .ZN(n734) );
  XNOR2_X1 U787 ( .A(n734), .B(KEYINPUT124), .ZN(n736) );
  NOR2_X1 U788 ( .A1(n736), .A2(n735), .ZN(n745) );
  NAND2_X1 U789 ( .A1(G953), .A2(G224), .ZN(n737) );
  XNOR2_X1 U790 ( .A(n737), .B(KEYINPUT61), .ZN(n739) );
  NAND2_X1 U791 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U792 ( .A(n740), .B(KEYINPUT123), .ZN(n743) );
  NOR2_X1 U793 ( .A1(G953), .A2(n741), .ZN(n742) );
  NOR2_X1 U794 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U795 ( .A(n745), .B(n744), .ZN(n746) );
  XNOR2_X1 U796 ( .A(n747), .B(n746), .ZN(G69) );
  XNOR2_X1 U797 ( .A(n749), .B(n748), .ZN(n753) );
  XNOR2_X1 U798 ( .A(n750), .B(n753), .ZN(n752) );
  NAND2_X1 U799 ( .A1(n752), .A2(n751), .ZN(n757) );
  XNOR2_X1 U800 ( .A(G227), .B(n753), .ZN(n754) );
  NAND2_X1 U801 ( .A1(n754), .A2(G900), .ZN(n755) );
  NAND2_X1 U802 ( .A1(n755), .A2(G953), .ZN(n756) );
  NAND2_X1 U803 ( .A1(n757), .A2(n756), .ZN(G72) );
  XOR2_X1 U804 ( .A(n758), .B(G122), .Z(G24) );
  XOR2_X1 U805 ( .A(G119), .B(n759), .Z(n760) );
  XNOR2_X1 U806 ( .A(KEYINPUT127), .B(n760), .ZN(G21) );
  XOR2_X1 U807 ( .A(n761), .B(G131), .Z(G33) );
  XOR2_X1 U808 ( .A(G137), .B(n762), .Z(G39) );
endmodule

