//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 1 1 1 1 1 0 0 1 1 1 0 0 1 0 1 0 0 1 0 1 0 1 1 0 0 0 1 1 0 0 1 0 1 0 1 0 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n784, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n972, new_n973;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT31), .B(G50gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT72), .ZN(new_n205));
  XOR2_X1   g004(.A(G197gat), .B(G204gat), .Z(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(KEYINPUT70), .B(G211gat), .ZN(new_n208));
  INV_X1    g007(.A(G218gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(KEYINPUT69), .B(KEYINPUT22), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n207), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(G211gat), .B(G218gat), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n213), .B(new_n207), .C1(new_n210), .C2(new_n211), .ZN(new_n216));
  AND3_X1   g015(.A1(new_n215), .A2(KEYINPUT71), .A3(new_n216), .ZN(new_n217));
  XOR2_X1   g016(.A(KEYINPUT70), .B(G211gat), .Z(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(G218gat), .ZN(new_n219));
  INV_X1    g018(.A(new_n211), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n206), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NOR3_X1   g020(.A1(new_n221), .A2(KEYINPUT71), .A3(new_n213), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n205), .B1(new_n217), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n222), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n215), .A2(KEYINPUT71), .A3(new_n216), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n224), .A2(KEYINPUT72), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(G148gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(G141gat), .ZN(new_n229));
  INV_X1    g028(.A(G141gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(G148gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(G155gat), .A2(G162gat), .ZN(new_n232));
  AOI22_X1  g031(.A1(new_n229), .A2(new_n231), .B1(KEYINPUT2), .B2(new_n232), .ZN(new_n233));
  NOR2_X1   g032(.A1(G155gat), .A2(G162gat), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(new_n232), .ZN(new_n236));
  AND2_X1   g035(.A1(new_n233), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT77), .ZN(new_n238));
  XNOR2_X1  g037(.A(G141gat), .B(G148gat), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT2), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n240), .B1(G155gat), .B2(G162gat), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n235), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n232), .A2(KEYINPUT76), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT76), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n244), .A2(G155gat), .A3(G162gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n238), .B1(new_n242), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n246), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n229), .A2(new_n231), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n232), .A2(KEYINPUT2), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n248), .A2(new_n251), .A3(KEYINPUT77), .A4(new_n235), .ZN(new_n252));
  AOI211_X1 g051(.A(KEYINPUT3), .B(new_n237), .C1(new_n247), .C2(new_n252), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n253), .A2(KEYINPUT29), .ZN(new_n254));
  OAI21_X1  g053(.A(KEYINPUT81), .B1(new_n227), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(G228gat), .ZN(new_n256));
  INV_X1    g055(.A(G233gat), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT3), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n224), .A2(new_n225), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n259), .B1(new_n260), .B2(KEYINPUT29), .ZN(new_n261));
  INV_X1    g060(.A(new_n237), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n234), .B1(new_n249), .B2(new_n250), .ZN(new_n263));
  AOI21_X1  g062(.A(KEYINPUT77), .B1(new_n263), .B2(new_n248), .ZN(new_n264));
  NOR4_X1   g063(.A1(new_n233), .A2(new_n246), .A3(new_n238), .A4(new_n234), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n262), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n261), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n254), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT81), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n268), .A2(new_n269), .A3(new_n223), .A4(new_n226), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n255), .A2(new_n258), .A3(new_n267), .A4(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(G22gat), .ZN(new_n272));
  INV_X1    g071(.A(new_n260), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n273), .A2(new_n254), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n237), .B1(new_n247), .B2(new_n252), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n215), .A2(new_n216), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT29), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n275), .B1(new_n278), .B2(new_n259), .ZN(new_n279));
  OAI22_X1  g078(.A1(new_n274), .A2(new_n279), .B1(new_n256), .B2(new_n257), .ZN(new_n280));
  AND3_X1   g079(.A1(new_n271), .A2(new_n272), .A3(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n272), .B1(new_n271), .B2(new_n280), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n204), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n271), .A2(new_n280), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(G22gat), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n271), .A2(new_n272), .A3(new_n280), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT82), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n204), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n285), .A2(new_n286), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n281), .A2(new_n287), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n283), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  OR2_X1    g090(.A1(new_n291), .A2(KEYINPUT83), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(KEYINPUT83), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n247), .A2(new_n252), .ZN(new_n295));
  INV_X1    g094(.A(G127gat), .ZN(new_n296));
  INV_X1    g095(.A(G134gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(G127gat), .A2(G134gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT67), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT68), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT1), .ZN(new_n303));
  AOI22_X1  g102(.A1(new_n300), .A2(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(KEYINPUT68), .A2(KEYINPUT1), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT66), .ZN(new_n306));
  INV_X1    g105(.A(G113gat), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n306), .B1(new_n307), .B2(G120gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(G120gat), .ZN(new_n309));
  INV_X1    g108(.A(G120gat), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n310), .A2(KEYINPUT66), .A3(G113gat), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n308), .A2(new_n309), .A3(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n298), .A2(KEYINPUT67), .A3(new_n299), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n304), .A2(new_n305), .A3(new_n312), .A4(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT65), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n310), .A2(G113gat), .ZN(new_n316));
  AOI21_X1  g115(.A(KEYINPUT1), .B1(new_n309), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n315), .B1(new_n317), .B2(new_n300), .ZN(new_n318));
  AND2_X1   g117(.A1(G127gat), .A2(G134gat), .ZN(new_n319));
  NOR2_X1   g118(.A1(G127gat), .A2(G134gat), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g120(.A(G113gat), .B(G120gat), .ZN(new_n322));
  OAI211_X1 g121(.A(new_n321), .B(KEYINPUT65), .C1(new_n322), .C2(KEYINPUT1), .ZN(new_n323));
  AND2_X1   g122(.A1(new_n318), .A2(new_n323), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n295), .A2(new_n314), .A3(new_n324), .A4(new_n262), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(KEYINPUT4), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n301), .B1(new_n319), .B2(new_n320), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n302), .A2(new_n303), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n312), .A2(new_n313), .A3(new_n327), .A4(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n305), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n318), .A2(new_n323), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT4), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n333), .A2(new_n275), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n326), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n266), .A2(KEYINPUT3), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n314), .A2(new_n318), .A3(new_n323), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n275), .A2(new_n259), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n336), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(G225gat), .A2(G233gat), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  NOR3_X1   g142(.A1(new_n341), .A2(KEYINPUT5), .A3(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n259), .B1(new_n295), .B2(new_n262), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n346), .A2(new_n253), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n343), .B1(new_n347), .B2(new_n338), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n335), .A2(KEYINPUT78), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT78), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n333), .A2(new_n275), .A3(new_n350), .A4(new_n334), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n349), .A2(new_n326), .A3(new_n351), .ZN(new_n352));
  AND2_X1   g151(.A1(new_n348), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT80), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n266), .A2(new_n338), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT79), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(new_n356), .A3(new_n325), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n266), .A2(KEYINPUT79), .A3(new_n338), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n357), .A2(new_n343), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(KEYINPUT5), .ZN(new_n360));
  NOR3_X1   g159(.A1(new_n353), .A2(new_n354), .A3(new_n360), .ZN(new_n361));
  AND2_X1   g160(.A1(new_n359), .A2(KEYINPUT5), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n348), .A2(new_n352), .ZN(new_n363));
  AOI21_X1  g162(.A(KEYINPUT80), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n345), .B1(new_n361), .B2(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(G1gat), .B(G29gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n366), .B(G85gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(KEYINPUT0), .B(G57gat), .ZN(new_n368));
  XOR2_X1   g167(.A(new_n367), .B(new_n368), .Z(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n365), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT6), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n354), .B1(new_n353), .B2(new_n360), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n362), .A2(KEYINPUT80), .A3(new_n363), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n344), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(KEYINPUT6), .B1(new_n377), .B2(new_n369), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(new_n371), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n374), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(G226gat), .A2(G233gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n381), .B(KEYINPUT73), .ZN(new_n382));
  INV_X1    g181(.A(G169gat), .ZN(new_n383));
  INV_X1    g182(.A(G176gat), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n383), .A2(new_n384), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(KEYINPUT26), .ZN(new_n388));
  NOR2_X1   g187(.A1(G169gat), .A2(G176gat), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT26), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n386), .A2(new_n388), .A3(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(G190gat), .ZN(new_n393));
  AND2_X1   g192(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n394));
  NOR2_X1   g193(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n393), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(KEYINPUT28), .ZN(new_n397));
  XNOR2_X1  g196(.A(KEYINPUT27), .B(G183gat), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT28), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n398), .A2(new_n399), .A3(new_n393), .ZN(new_n400));
  NAND2_X1  g199(.A1(G183gat), .A2(G190gat), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n392), .A2(new_n397), .A3(new_n400), .A4(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  OR2_X1    g202(.A1(G183gat), .A2(G190gat), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n404), .A2(KEYINPUT24), .A3(new_n401), .ZN(new_n405));
  OR2_X1    g204(.A1(new_n401), .A2(KEYINPUT24), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT23), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n387), .A2(new_n407), .ZN(new_n408));
  AND4_X1   g207(.A1(new_n386), .A2(new_n405), .A3(new_n406), .A4(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n389), .A2(KEYINPUT23), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT64), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n409), .B(new_n410), .C1(new_n411), .C2(KEYINPUT25), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n385), .B1(new_n407), .B2(new_n387), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n413), .A2(new_n411), .A3(new_n406), .A4(new_n405), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n413), .A2(new_n406), .A3(new_n405), .A4(new_n410), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT25), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n403), .B1(new_n412), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n382), .B1(new_n418), .B2(KEYINPUT29), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT74), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n412), .A2(new_n417), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(new_n402), .ZN(new_n423));
  INV_X1    g222(.A(new_n381), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  OAI211_X1 g224(.A(KEYINPUT74), .B(new_n382), .C1(new_n418), .C2(KEYINPUT29), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n421), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n227), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n424), .B1(new_n423), .B2(new_n277), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n418), .A2(new_n382), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AOI22_X1  g230(.A1(new_n427), .A2(new_n428), .B1(new_n431), .B2(new_n273), .ZN(new_n432));
  XNOR2_X1  g231(.A(G8gat), .B(G36gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(G64gat), .B(G92gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n433), .B(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n427), .A2(new_n428), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n431), .A2(new_n273), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n438), .A2(new_n439), .A3(new_n436), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n437), .B1(new_n441), .B2(KEYINPUT30), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT75), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT30), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n432), .A2(KEYINPUT75), .A3(new_n436), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n442), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n380), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n294), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g250(.A(G15gat), .B(G43gat), .ZN(new_n452));
  XNOR2_X1  g251(.A(G71gat), .B(G99gat), .ZN(new_n453));
  XOR2_X1   g252(.A(new_n452), .B(new_n453), .Z(new_n454));
  NAND2_X1  g253(.A1(new_n423), .A2(new_n338), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n418), .A2(new_n333), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n457), .A2(G227gat), .A3(G233gat), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n454), .B1(new_n459), .B2(KEYINPUT33), .ZN(new_n460));
  INV_X1    g259(.A(G227gat), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n455), .B(new_n456), .C1(new_n461), .C2(new_n257), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT34), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n463), .B1(new_n458), .B2(KEYINPUT32), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n458), .A2(KEYINPUT32), .A3(new_n463), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n466), .ZN(new_n468));
  INV_X1    g267(.A(new_n462), .ZN(new_n469));
  NOR3_X1   g268(.A1(new_n468), .A2(new_n464), .A3(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n460), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n469), .B1(new_n468), .B2(new_n464), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n465), .A2(new_n466), .A3(new_n462), .ZN(new_n473));
  INV_X1    g272(.A(new_n460), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  AND3_X1   g274(.A1(new_n471), .A2(KEYINPUT36), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT36), .B1(new_n471), .B2(new_n475), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT84), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n478), .B1(new_n365), .B2(new_n370), .ZN(new_n479));
  NOR3_X1   g278(.A1(new_n377), .A2(KEYINPUT84), .A3(new_n369), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n378), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT37), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n436), .B1(new_n432), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n260), .B1(new_n429), .B2(new_n430), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n484), .B1(new_n427), .B2(new_n428), .ZN(new_n485));
  AOI21_X1  g284(.A(KEYINPUT38), .B1(new_n485), .B2(KEYINPUT37), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n487), .A2(new_n444), .A3(new_n446), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT38), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n438), .A2(new_n439), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT37), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n489), .B1(new_n483), .B2(new_n491), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n481), .A2(new_n493), .A3(new_n374), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n341), .A2(new_n343), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n357), .A2(new_n358), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(new_n342), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n495), .A2(KEYINPUT39), .A3(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT40), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n342), .B1(new_n336), .B2(new_n340), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT39), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n370), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  AND3_X1   g301(.A1(new_n498), .A2(new_n499), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n499), .B1(new_n498), .B2(new_n502), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT84), .B1(new_n377), .B2(new_n369), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n365), .A2(new_n478), .A3(new_n370), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n291), .B1(new_n508), .B2(new_n448), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT85), .ZN(new_n510));
  AND3_X1   g309(.A1(new_n494), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n510), .B1(new_n494), .B2(new_n509), .ZN(new_n512));
  OAI221_X1 g311(.A(new_n451), .B1(new_n476), .B2(new_n477), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n471), .A2(new_n475), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n514), .A2(new_n291), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(KEYINPUT35), .B1(new_n450), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n481), .A2(new_n374), .ZN(new_n518));
  XOR2_X1   g317(.A(KEYINPUT86), .B(KEYINPUT35), .Z(new_n519));
  NAND4_X1  g318(.A1(new_n518), .A2(new_n515), .A3(new_n449), .A4(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n513), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(G29gat), .ZN(new_n523));
  INV_X1    g322(.A(G36gat), .ZN(new_n524));
  OR3_X1    g323(.A1(new_n523), .A2(new_n524), .A3(KEYINPUT88), .ZN(new_n525));
  OAI21_X1  g324(.A(KEYINPUT88), .B1(new_n523), .B2(new_n524), .ZN(new_n526));
  OAI21_X1  g325(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  NOR3_X1   g327(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n525), .B(new_n526), .C1(new_n528), .C2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(G50gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(G43gat), .ZN(new_n532));
  AOI21_X1  g331(.A(KEYINPUT15), .B1(new_n532), .B2(KEYINPUT89), .ZN(new_n533));
  OR2_X1    g332(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(G43gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(G50gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n532), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  OR2_X1    g337(.A1(new_n534), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT15), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n537), .B1(new_n530), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n534), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(KEYINPUT17), .ZN(new_n544));
  XNOR2_X1  g343(.A(G15gat), .B(G22gat), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT16), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n545), .B1(new_n546), .B2(G1gat), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n547), .B1(G1gat), .B2(new_n545), .ZN(new_n548));
  INV_X1    g347(.A(G8gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n548), .B(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(KEYINPUT90), .ZN(new_n552));
  OR2_X1    g351(.A1(new_n551), .A2(KEYINPUT90), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n544), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n543), .A2(new_n551), .ZN(new_n555));
  NAND2_X1  g354(.A1(G229gat), .A2(G233gat), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT91), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(KEYINPUT18), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n543), .B(new_n551), .ZN(new_n560));
  XOR2_X1   g359(.A(new_n556), .B(KEYINPUT13), .Z(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT18), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n557), .A2(KEYINPUT91), .A3(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n559), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  XOR2_X1   g364(.A(KEYINPUT87), .B(KEYINPUT11), .Z(new_n566));
  XNOR2_X1  g365(.A(G169gat), .B(G197gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G113gat), .B(G141gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(new_n570), .B(KEYINPUT12), .Z(new_n571));
  NAND2_X1  g370(.A1(new_n565), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n571), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n559), .A2(new_n573), .A3(new_n562), .A4(new_n564), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n572), .A2(KEYINPUT92), .A3(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT92), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n565), .A2(new_n576), .A3(new_n571), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(G85gat), .A2(G92gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(KEYINPUT7), .ZN(new_n581));
  INV_X1    g380(.A(G99gat), .ZN(new_n582));
  INV_X1    g381(.A(G106gat), .ZN(new_n583));
  OAI21_X1  g382(.A(KEYINPUT8), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  OAI211_X1 g383(.A(new_n581), .B(new_n584), .C1(G85gat), .C2(G92gat), .ZN(new_n585));
  XOR2_X1   g384(.A(G99gat), .B(G106gat), .Z(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(KEYINPUT95), .ZN(new_n588));
  AND2_X1   g387(.A1(new_n544), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT96), .ZN(new_n590));
  INV_X1    g389(.A(new_n543), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT41), .ZN(new_n592));
  NAND2_X1  g391(.A1(G232gat), .A2(G233gat), .ZN(new_n593));
  OAI22_X1  g392(.A1(new_n591), .A2(new_n587), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  OR3_X1    g393(.A1(new_n589), .A2(new_n590), .A3(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n590), .B1(new_n589), .B2(new_n594), .ZN(new_n596));
  XNOR2_X1  g395(.A(G190gat), .B(G218gat), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  OR2_X1    g397(.A1(new_n596), .A2(new_n597), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G134gat), .B(G162gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n593), .A2(new_n592), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n603), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n598), .A2(new_n599), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G127gat), .B(G155gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(G211gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(G71gat), .B(G78gat), .ZN(new_n612));
  XOR2_X1   g411(.A(new_n612), .B(KEYINPUT93), .Z(new_n613));
  XNOR2_X1  g412(.A(G57gat), .B(G64gat), .ZN(new_n614));
  AOI21_X1  g413(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n615), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT94), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n617), .B1(new_n614), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n614), .A2(new_n618), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(new_n612), .ZN(new_n621));
  OAI22_X1  g420(.A1(new_n613), .A2(new_n616), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT21), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n550), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(G183gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n622), .A2(new_n623), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  AND2_X1   g426(.A1(G231gat), .A2(G233gat), .ZN(new_n628));
  AND2_X1   g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n627), .A2(new_n628), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n611), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NOR3_X1   g431(.A1(new_n629), .A2(new_n630), .A3(new_n611), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n609), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n633), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n635), .A2(new_n608), .A3(new_n631), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n607), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G120gat), .B(G148gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(G176gat), .B(G204gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(G230gat), .A2(G233gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(KEYINPUT99), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n587), .B1(new_n622), .B2(KEYINPUT97), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n622), .A2(KEYINPUT97), .ZN(new_n646));
  XOR2_X1   g445(.A(new_n645), .B(new_n646), .Z(new_n647));
  INV_X1    g446(.A(KEYINPUT10), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT98), .ZN(new_n649));
  NOR3_X1   g448(.A1(new_n587), .A2(new_n622), .A3(new_n648), .ZN(new_n650));
  AOI22_X1  g449(.A1(new_n647), .A2(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  OR2_X1    g450(.A1(new_n650), .A2(new_n649), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n643), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT100), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI211_X1 g454(.A(KEYINPUT100), .B(new_n643), .C1(new_n651), .C2(new_n652), .ZN(new_n656));
  OAI221_X1 g455(.A(new_n641), .B1(new_n644), .B2(new_n647), .C1(new_n655), .C2(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n647), .A2(new_n644), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n640), .B1(new_n653), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n637), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n522), .A2(new_n579), .A3(new_n661), .ZN(new_n662));
  AND2_X1   g461(.A1(new_n662), .A2(KEYINPUT101), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n662), .A2(KEYINPUT101), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n380), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g468(.A1(new_n665), .A2(new_n449), .ZN(new_n670));
  NAND2_X1  g469(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n546), .A2(new_n549), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT42), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n670), .A2(KEYINPUT42), .A3(new_n671), .A4(new_n672), .ZN(new_n676));
  OAI211_X1 g475(.A(new_n675), .B(new_n676), .C1(new_n549), .C2(new_n670), .ZN(G1325gat));
  INV_X1    g476(.A(new_n514), .ZN(new_n678));
  AOI21_X1  g477(.A(G15gat), .B1(new_n666), .B2(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(KEYINPUT102), .B1(new_n476), .B2(new_n477), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT36), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n514), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT102), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n471), .A2(KEYINPUT36), .A3(new_n475), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n680), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  OR2_X1    g486(.A1(new_n687), .A2(KEYINPUT103), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(KEYINPUT103), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(G15gat), .ZN(new_n692));
  XOR2_X1   g491(.A(new_n692), .B(KEYINPUT104), .Z(new_n693));
  AOI21_X1  g492(.A(new_n679), .B1(new_n666), .B2(new_n693), .ZN(G1326gat));
  NAND3_X1  g493(.A1(new_n666), .A2(new_n272), .A3(new_n294), .ZN(new_n695));
  INV_X1    g494(.A(new_n294), .ZN(new_n696));
  OAI21_X1  g495(.A(G22gat), .B1(new_n665), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(KEYINPUT105), .B(KEYINPUT43), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1327gat));
  AOI21_X1  g499(.A(new_n607), .B1(new_n513), .B2(new_n521), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n634), .A2(new_n636), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n703), .A2(new_n578), .A3(new_n660), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n705), .A2(new_n523), .A3(new_n667), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(KEYINPUT45), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708));
  OAI211_X1 g507(.A(new_n451), .B(new_n686), .C1(new_n511), .C2(new_n512), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT106), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n372), .B1(new_n365), .B2(new_n370), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n712), .B1(new_n506), .B2(new_n507), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n483), .A2(new_n491), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(KEYINPUT38), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n444), .A2(new_n446), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n715), .A2(new_n716), .A3(new_n487), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n713), .A2(new_n717), .A3(new_n373), .ZN(new_n718));
  INV_X1    g517(.A(new_n291), .ZN(new_n719));
  INV_X1    g518(.A(new_n505), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n720), .B1(new_n479), .B2(new_n480), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n719), .B1(new_n721), .B2(new_n449), .ZN(new_n722));
  OAI21_X1  g521(.A(KEYINPUT85), .B1(new_n718), .B2(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n494), .A2(new_n509), .A3(new_n510), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n725), .A2(KEYINPUT106), .A3(new_n451), .A4(new_n686), .ZN(new_n726));
  AOI22_X1  g525(.A1(new_n711), .A2(new_n726), .B1(new_n517), .B2(new_n520), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n708), .B1(new_n727), .B2(new_n607), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n701), .A2(KEYINPUT44), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n728), .A2(new_n729), .A3(new_n704), .ZN(new_n730));
  OAI21_X1  g529(.A(G29gat), .B1(new_n730), .B2(new_n380), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n707), .A2(new_n731), .ZN(G1328gat));
  OR2_X1    g531(.A1(new_n730), .A2(new_n449), .ZN(new_n733));
  OR2_X1    g532(.A1(new_n733), .A2(KEYINPUT107), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(KEYINPUT107), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n734), .A2(G36gat), .A3(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n705), .A2(new_n524), .A3(new_n448), .ZN(new_n737));
  XOR2_X1   g536(.A(new_n737), .B(KEYINPUT46), .Z(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(new_n738), .ZN(G1329gat));
  OAI21_X1  g538(.A(G43gat), .B1(new_n730), .B2(new_n686), .ZN(new_n740));
  AND3_X1   g539(.A1(new_n705), .A2(new_n535), .A3(new_n678), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n740), .A2(KEYINPUT47), .A3(new_n742), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n728), .A2(new_n691), .A3(new_n729), .A4(new_n704), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT108), .ZN(new_n745));
  AND3_X1   g544(.A1(new_n744), .A2(new_n745), .A3(G43gat), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n745), .B1(new_n744), .B2(G43gat), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n746), .A2(new_n747), .A3(new_n741), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n743), .B1(new_n748), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g548(.A(KEYINPUT48), .ZN(new_n750));
  OAI21_X1  g549(.A(G50gat), .B1(new_n730), .B2(new_n719), .ZN(new_n751));
  AND3_X1   g550(.A1(new_n705), .A2(new_n531), .A3(new_n294), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(KEYINPUT109), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n750), .B1(new_n751), .B2(new_n753), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n752), .B1(KEYINPUT109), .B2(KEYINPUT48), .ZN(new_n755));
  OAI211_X1 g554(.A(new_n750), .B(G50gat), .C1(new_n730), .C2(new_n696), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n754), .B1(new_n755), .B2(new_n756), .ZN(G1331gat));
  INV_X1    g556(.A(new_n660), .ZN(new_n758));
  NOR4_X1   g557(.A1(new_n727), .A2(new_n579), .A3(new_n637), .A4(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(new_n667), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g560(.A1(new_n711), .A2(new_n726), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n521), .ZN(new_n763));
  INV_X1    g562(.A(new_n637), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n579), .A2(new_n758), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT110), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n767), .A2(new_n449), .ZN(new_n768));
  NOR2_X1   g567(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n769));
  AND2_X1   g568(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n768), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n771), .B1(new_n768), .B2(new_n769), .ZN(G1333gat));
  INV_X1    g571(.A(KEYINPUT50), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n759), .A2(KEYINPUT110), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT110), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n766), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n691), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(G71gat), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n766), .A2(G71gat), .A3(new_n514), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n773), .B1(new_n778), .B2(new_n780), .ZN(new_n781));
  AOI211_X1 g580(.A(KEYINPUT50), .B(new_n779), .C1(new_n777), .C2(G71gat), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n781), .A2(new_n782), .ZN(G1334gat));
  NOR2_X1   g582(.A1(new_n767), .A2(new_n696), .ZN(new_n784));
  XOR2_X1   g583(.A(new_n784), .B(G78gat), .Z(G1335gat));
  INV_X1    g584(.A(new_n607), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n579), .A2(new_n703), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n763), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(KEYINPUT51), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n607), .B1(new_n762), .B2(new_n521), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT51), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n790), .A2(new_n791), .A3(new_n787), .ZN(new_n792));
  AND3_X1   g591(.A1(new_n789), .A2(new_n660), .A3(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(G85gat), .B1(new_n793), .B2(new_n667), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n579), .A2(new_n703), .A3(new_n758), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n729), .B(new_n795), .C1(new_n790), .C2(KEYINPUT44), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(KEYINPUT111), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT111), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n728), .A2(new_n798), .A3(new_n729), .A4(new_n795), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n380), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n794), .B1(G85gat), .B2(new_n800), .ZN(G1336gat));
  INV_X1    g600(.A(G92gat), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n797), .A2(new_n799), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n802), .B1(new_n803), .B2(new_n448), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n449), .A2(G92gat), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n789), .A2(new_n660), .A3(new_n792), .A4(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(KEYINPUT52), .B1(new_n804), .B2(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(G92gat), .B1(new_n796), .B2(new_n449), .ZN(new_n809));
  XNOR2_X1  g608(.A(KEYINPUT112), .B(KEYINPUT52), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n806), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(KEYINPUT113), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT113), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n806), .A2(new_n809), .A3(new_n813), .A4(new_n810), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n808), .A2(new_n815), .ZN(G1337gat));
  XNOR2_X1  g615(.A(KEYINPUT115), .B(G99gat), .ZN(new_n817));
  AOI21_X1  g616(.A(KEYINPUT114), .B1(new_n803), .B2(new_n691), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT114), .ZN(new_n819));
  AOI211_X1 g618(.A(new_n819), .B(new_n690), .C1(new_n797), .C2(new_n799), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n817), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n817), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n793), .A2(new_n678), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(new_n823), .ZN(G1338gat));
  AOI21_X1  g623(.A(new_n583), .B1(new_n803), .B2(new_n294), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n789), .A2(new_n583), .A3(new_n660), .A4(new_n792), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n826), .A2(new_n719), .ZN(new_n827));
  OAI21_X1  g626(.A(KEYINPUT53), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n827), .A2(KEYINPUT53), .ZN(new_n829));
  OAI21_X1  g628(.A(G106gat), .B1(new_n796), .B2(new_n719), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n828), .A2(new_n831), .ZN(G1339gat));
  NOR3_X1   g631(.A1(new_n579), .A2(new_n637), .A3(new_n660), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n556), .B1(new_n554), .B2(new_n555), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n560), .A2(new_n561), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n570), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OR2_X1    g635(.A1(new_n836), .A2(KEYINPUT116), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(KEYINPUT116), .ZN(new_n838));
  AND3_X1   g637(.A1(new_n574), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n660), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n651), .A2(new_n643), .A3(new_n652), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n841), .B(KEYINPUT54), .C1(new_n655), .C2(new_n656), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT55), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n641), .B1(new_n653), .B2(new_n844), .ZN(new_n845));
  AND3_X1   g644(.A1(new_n842), .A2(new_n843), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n843), .B1(new_n842), .B2(new_n845), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n657), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI211_X1 g647(.A(new_n607), .B(new_n840), .C1(new_n848), .C2(new_n578), .ZN(new_n849));
  OAI211_X1 g648(.A(new_n657), .B(new_n839), .C1(new_n846), .C2(new_n847), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n703), .B1(new_n850), .B2(new_n786), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n833), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n852), .A2(new_n516), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n380), .A2(new_n448), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n307), .B1(new_n855), .B2(new_n578), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n852), .A2(new_n294), .A3(new_n514), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n854), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n579), .A2(G113gat), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n856), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  XOR2_X1   g659(.A(new_n860), .B(KEYINPUT117), .Z(G1340gat));
  OAI21_X1  g660(.A(G120gat), .B1(new_n858), .B2(new_n758), .ZN(new_n862));
  XOR2_X1   g661(.A(new_n862), .B(KEYINPUT118), .Z(new_n863));
  NAND2_X1  g662(.A1(new_n660), .A2(new_n310), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n863), .B1(new_n855), .B2(new_n864), .ZN(G1341gat));
  NOR3_X1   g664(.A1(new_n858), .A2(new_n296), .A3(new_n702), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT119), .ZN(new_n867));
  OR2_X1    g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n296), .B1(new_n855), .B2(new_n702), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n866), .A2(new_n867), .ZN(new_n870));
  AND3_X1   g669(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(G1342gat));
  NAND2_X1  g670(.A1(new_n786), .A2(new_n449), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n872), .B(KEYINPUT120), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n853), .A2(new_n297), .A3(new_n667), .A4(new_n873), .ZN(new_n874));
  XOR2_X1   g673(.A(new_n874), .B(KEYINPUT56), .Z(new_n875));
  OAI21_X1  g674(.A(G134gat), .B1(new_n858), .B2(new_n607), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(G1343gat));
  NAND2_X1  g676(.A1(new_n849), .A2(new_n851), .ZN(new_n878));
  INV_X1    g677(.A(new_n833), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(new_n291), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n881), .A2(new_n691), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n882), .A2(new_n230), .A3(new_n579), .A4(new_n854), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT58), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT57), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n880), .A2(new_n886), .A3(new_n291), .ZN(new_n887));
  OAI21_X1  g686(.A(KEYINPUT57), .B1(new_n852), .B2(new_n696), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n686), .A2(new_n854), .ZN(new_n889));
  INV_X1    g688(.A(new_n889), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n887), .A2(new_n888), .A3(new_n579), .A4(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT121), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n891), .B(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n885), .B1(new_n893), .B2(G141gat), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n891), .A2(G141gat), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n884), .B1(new_n895), .B2(new_n883), .ZN(new_n896));
  OAI21_X1  g695(.A(KEYINPUT122), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n887), .A2(new_n890), .A3(new_n888), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n892), .A3(new_n579), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n891), .A2(KEYINPUT121), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n899), .A2(G141gat), .A3(new_n900), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n901), .A2(new_n884), .A3(new_n883), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT122), .ZN(new_n903));
  INV_X1    g702(.A(new_n896), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n897), .A2(new_n905), .ZN(G1344gat));
  INV_X1    g705(.A(KEYINPUT59), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n881), .A2(KEYINPUT57), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n880), .A2(new_n886), .A3(new_n294), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n910), .A2(new_n660), .A3(new_n890), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n907), .B1(new_n911), .B2(G148gat), .ZN(new_n912));
  AOI211_X1 g711(.A(KEYINPUT59), .B(new_n228), .C1(new_n898), .C2(new_n660), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n882), .A2(new_n854), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n660), .A2(new_n228), .ZN(new_n915));
  OAI22_X1  g714(.A1(new_n912), .A2(new_n913), .B1(new_n914), .B2(new_n915), .ZN(G1345gat));
  NAND3_X1  g715(.A1(new_n882), .A2(new_n703), .A3(new_n854), .ZN(new_n917));
  INV_X1    g716(.A(G155gat), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n702), .A2(new_n918), .ZN(new_n919));
  AOI22_X1  g718(.A1(new_n917), .A2(new_n918), .B1(new_n898), .B2(new_n919), .ZN(G1346gat));
  INV_X1    g719(.A(G162gat), .ZN(new_n921));
  NAND4_X1  g720(.A1(new_n882), .A2(new_n921), .A3(new_n667), .A4(new_n873), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n898), .A2(new_n786), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n922), .B1(new_n923), .B2(new_n921), .ZN(G1347gat));
  NOR2_X1   g723(.A1(new_n667), .A2(new_n449), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n853), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n926), .B(KEYINPUT123), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n927), .A2(new_n383), .A3(new_n579), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n857), .A2(new_n925), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(G169gat), .B1(new_n930), .B2(new_n578), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n928), .A2(new_n931), .ZN(G1348gat));
  AOI21_X1  g731(.A(G176gat), .B1(new_n927), .B2(new_n660), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n758), .A2(new_n384), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n933), .B1(new_n929), .B2(new_n934), .ZN(G1349gat));
  INV_X1    g734(.A(new_n398), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n926), .A2(new_n936), .A3(new_n702), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n929), .A2(new_n703), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n937), .B1(new_n938), .B2(G183gat), .ZN(new_n939));
  AND4_X1   g738(.A1(KEYINPUT124), .A2(new_n939), .A3(KEYINPUT125), .A4(KEYINPUT60), .ZN(new_n940));
  AOI21_X1  g739(.A(KEYINPUT60), .B1(new_n939), .B2(KEYINPUT125), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n939), .A2(KEYINPUT124), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(G1350gat));
  NAND3_X1  g742(.A1(new_n927), .A2(new_n393), .A3(new_n786), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n393), .B1(new_n929), .B2(new_n786), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT61), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n945), .A2(new_n946), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n944), .B1(new_n947), .B2(new_n948), .ZN(G1351gat));
  AND2_X1   g748(.A1(new_n690), .A2(new_n925), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n950), .A2(new_n291), .A3(new_n880), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(G197gat), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n952), .A2(new_n953), .A3(new_n579), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n910), .A2(new_n950), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n955), .A2(new_n579), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n954), .B1(new_n956), .B2(new_n953), .ZN(G1352gat));
  NOR3_X1   g756(.A1(new_n951), .A2(G204gat), .A3(new_n758), .ZN(new_n958));
  XNOR2_X1  g757(.A(new_n958), .B(KEYINPUT62), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n910), .A2(new_n660), .A3(new_n950), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(G204gat), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n959), .A2(new_n961), .ZN(G1353gat));
  NAND3_X1  g761(.A1(new_n952), .A2(new_n208), .A3(new_n703), .ZN(new_n963));
  NAND4_X1  g762(.A1(new_n908), .A2(new_n703), .A3(new_n909), .A4(new_n950), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(KEYINPUT126), .ZN(new_n965));
  AOI21_X1  g764(.A(KEYINPUT63), .B1(new_n965), .B2(G211gat), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT126), .ZN(new_n967));
  OR2_X1    g766(.A1(new_n964), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n964), .A2(new_n967), .ZN(new_n969));
  AND4_X1   g768(.A1(KEYINPUT63), .A2(new_n968), .A3(G211gat), .A4(new_n969), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n963), .B1(new_n966), .B2(new_n970), .ZN(G1354gat));
  NAND3_X1  g770(.A1(new_n952), .A2(new_n209), .A3(new_n786), .ZN(new_n972));
  AND2_X1   g771(.A1(new_n955), .A2(new_n786), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n972), .B1(new_n973), .B2(new_n209), .ZN(G1355gat));
endmodule


