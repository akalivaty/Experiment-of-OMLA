

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589;

  INV_X1 U324 ( .A(n392), .ZN(n375) );
  XNOR2_X1 U325 ( .A(n406), .B(n380), .ZN(n381) );
  XNOR2_X1 U326 ( .A(n413), .B(n412), .ZN(n414) );
  INV_X1 U327 ( .A(n411), .ZN(n412) );
  XNOR2_X1 U328 ( .A(n490), .B(n489), .ZN(n530) );
  XNOR2_X1 U329 ( .A(n376), .B(n375), .ZN(n383) );
  XOR2_X1 U330 ( .A(KEYINPUT45), .B(n422), .Z(n292) );
  XOR2_X1 U331 ( .A(G85GAT), .B(KEYINPUT73), .Z(n293) );
  INV_X1 U332 ( .A(KEYINPUT54), .ZN(n455) );
  XNOR2_X1 U333 ( .A(n455), .B(KEYINPUT118), .ZN(n456) );
  XNOR2_X1 U334 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U335 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U336 ( .A(n410), .B(n332), .ZN(n333) );
  XNOR2_X1 U337 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U338 ( .A(n488), .B(KEYINPUT105), .ZN(n489) );
  XNOR2_X1 U339 ( .A(n334), .B(n333), .ZN(n338) );
  XNOR2_X1 U340 ( .A(n383), .B(n382), .ZN(n385) );
  NOR2_X1 U341 ( .A1(n518), .A2(n448), .ZN(n449) );
  INV_X1 U342 ( .A(G127GAT), .ZN(n450) );
  INV_X1 U343 ( .A(G43GAT), .ZN(n493) );
  XOR2_X1 U344 ( .A(n342), .B(n384), .Z(n534) );
  XNOR2_X1 U345 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U346 ( .A(n450), .B(KEYINPUT50), .ZN(n451) );
  XNOR2_X1 U347 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U348 ( .A(n470), .B(n469), .ZN(G1351GAT) );
  XNOR2_X1 U349 ( .A(n496), .B(n495), .ZN(G1330GAT) );
  XOR2_X1 U350 ( .A(G78GAT), .B(G211GAT), .Z(n295) );
  XNOR2_X1 U351 ( .A(G22GAT), .B(G155GAT), .ZN(n294) );
  XNOR2_X1 U352 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U353 ( .A(G64GAT), .B(G71GAT), .Z(n297) );
  XNOR2_X1 U354 ( .A(G183GAT), .B(G127GAT), .ZN(n296) );
  XNOR2_X1 U355 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U356 ( .A(n299), .B(n298), .Z(n304) );
  XOR2_X1 U357 ( .A(KEYINPUT14), .B(KEYINPUT82), .Z(n301) );
  NAND2_X1 U358 ( .A1(G231GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U359 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U360 ( .A(KEYINPUT12), .B(n302), .ZN(n303) );
  XNOR2_X1 U361 ( .A(n304), .B(n303), .ZN(n308) );
  XOR2_X1 U362 ( .A(KEYINPUT84), .B(KEYINPUT15), .Z(n306) );
  XNOR2_X1 U363 ( .A(G8GAT), .B(KEYINPUT83), .ZN(n305) );
  XNOR2_X1 U364 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U365 ( .A(n308), .B(n307), .Z(n313) );
  XNOR2_X1 U366 ( .A(G15GAT), .B(G1GAT), .ZN(n309) );
  XNOR2_X1 U367 ( .A(n309), .B(KEYINPUT65), .ZN(n397) );
  XOR2_X1 U368 ( .A(KEYINPUT68), .B(KEYINPUT69), .Z(n311) );
  XNOR2_X1 U369 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n310) );
  XNOR2_X1 U370 ( .A(n311), .B(n310), .ZN(n411) );
  XNOR2_X1 U371 ( .A(n397), .B(n411), .ZN(n312) );
  XOR2_X1 U372 ( .A(n313), .B(n312), .Z(n581) );
  INV_X1 U373 ( .A(n581), .ZN(n567) );
  XOR2_X1 U374 ( .A(KEYINPUT23), .B(G106GAT), .Z(n315) );
  XNOR2_X1 U375 ( .A(G50GAT), .B(G218GAT), .ZN(n314) );
  XNOR2_X1 U376 ( .A(n315), .B(n314), .ZN(n330) );
  XOR2_X1 U377 ( .A(KEYINPUT24), .B(KEYINPUT90), .Z(n317) );
  NAND2_X1 U378 ( .A1(G228GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U379 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U380 ( .A(n318), .B(KEYINPUT22), .Z(n324) );
  XOR2_X1 U381 ( .A(G155GAT), .B(KEYINPUT3), .Z(n320) );
  XNOR2_X1 U382 ( .A(KEYINPUT91), .B(KEYINPUT2), .ZN(n319) );
  XNOR2_X1 U383 ( .A(n320), .B(n319), .ZN(n361) );
  XOR2_X1 U384 ( .A(G204GAT), .B(G211GAT), .Z(n322) );
  XNOR2_X1 U385 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n321) );
  XNOR2_X1 U386 ( .A(n322), .B(n321), .ZN(n331) );
  XNOR2_X1 U387 ( .A(n361), .B(n331), .ZN(n323) );
  XNOR2_X1 U388 ( .A(n324), .B(n323), .ZN(n326) );
  XNOR2_X1 U389 ( .A(G78GAT), .B(KEYINPUT72), .ZN(n325) );
  XNOR2_X1 U390 ( .A(n325), .B(G148GAT), .ZN(n407) );
  XOR2_X1 U391 ( .A(n326), .B(n407), .Z(n328) );
  XOR2_X1 U392 ( .A(G141GAT), .B(G22GAT), .Z(n398) );
  XOR2_X1 U393 ( .A(KEYINPUT74), .B(G162GAT), .Z(n379) );
  XNOR2_X1 U394 ( .A(n398), .B(n379), .ZN(n327) );
  XNOR2_X1 U395 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U396 ( .A(n330), .B(n329), .ZN(n476) );
  XNOR2_X1 U397 ( .A(KEYINPUT28), .B(n476), .ZN(n541) );
  INV_X1 U398 ( .A(n541), .ZN(n518) );
  XOR2_X1 U399 ( .A(KEYINPUT95), .B(n331), .Z(n334) );
  XOR2_X1 U400 ( .A(G176GAT), .B(G64GAT), .Z(n410) );
  NAND2_X1 U401 ( .A1(G226GAT), .A2(G233GAT), .ZN(n332) );
  XOR2_X1 U402 ( .A(G169GAT), .B(G8GAT), .Z(n395) );
  XOR2_X1 U403 ( .A(G183GAT), .B(KEYINPUT18), .Z(n336) );
  XNOR2_X1 U404 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n335) );
  XNOR2_X1 U405 ( .A(n336), .B(n335), .ZN(n443) );
  XOR2_X1 U406 ( .A(n395), .B(n443), .Z(n337) );
  XNOR2_X1 U407 ( .A(n338), .B(n337), .ZN(n342) );
  XOR2_X1 U408 ( .A(KEYINPUT80), .B(G92GAT), .Z(n340) );
  XNOR2_X1 U409 ( .A(G190GAT), .B(G218GAT), .ZN(n339) );
  XNOR2_X1 U410 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U411 ( .A(G36GAT), .B(n341), .ZN(n384) );
  XOR2_X1 U412 ( .A(n534), .B(KEYINPUT27), .Z(n343) );
  XNOR2_X1 U413 ( .A(n343), .B(KEYINPUT96), .ZN(n479) );
  XOR2_X1 U414 ( .A(G85GAT), .B(G148GAT), .Z(n345) );
  XNOR2_X1 U415 ( .A(G29GAT), .B(G162GAT), .ZN(n344) );
  XNOR2_X1 U416 ( .A(n345), .B(n344), .ZN(n349) );
  XOR2_X1 U417 ( .A(KEYINPUT94), .B(G120GAT), .Z(n347) );
  XNOR2_X1 U418 ( .A(G141GAT), .B(G1GAT), .ZN(n346) );
  XNOR2_X1 U419 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U420 ( .A(n349), .B(n348), .Z(n354) );
  XOR2_X1 U421 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n351) );
  NAND2_X1 U422 ( .A1(G225GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U423 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U424 ( .A(KEYINPUT93), .B(n352), .ZN(n353) );
  XNOR2_X1 U425 ( .A(n354), .B(n353), .ZN(n358) );
  XOR2_X1 U426 ( .A(G57GAT), .B(KEYINPUT92), .Z(n356) );
  XNOR2_X1 U427 ( .A(KEYINPUT1), .B(KEYINPUT6), .ZN(n355) );
  XNOR2_X1 U428 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U429 ( .A(n358), .B(n357), .Z(n363) );
  XOR2_X1 U430 ( .A(G127GAT), .B(KEYINPUT0), .Z(n360) );
  XNOR2_X1 U431 ( .A(G113GAT), .B(G134GAT), .ZN(n359) );
  XNOR2_X1 U432 ( .A(n360), .B(n359), .ZN(n442) );
  XNOR2_X1 U433 ( .A(n442), .B(n361), .ZN(n362) );
  XOR2_X1 U434 ( .A(n363), .B(n362), .Z(n532) );
  INV_X1 U435 ( .A(KEYINPUT10), .ZN(n367) );
  XOR2_X1 U436 ( .A(KEYINPUT78), .B(KEYINPUT11), .Z(n365) );
  XNOR2_X1 U437 ( .A(KEYINPUT76), .B(KEYINPUT77), .ZN(n364) );
  XNOR2_X1 U438 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U439 ( .A(n367), .B(n366), .ZN(n369) );
  NAND2_X1 U440 ( .A1(G232GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U441 ( .A(n369), .B(n368), .ZN(n371) );
  INV_X1 U442 ( .A(KEYINPUT75), .ZN(n370) );
  XNOR2_X1 U443 ( .A(n371), .B(n370), .ZN(n376) );
  XOR2_X1 U444 ( .A(KEYINPUT8), .B(G50GAT), .Z(n373) );
  XNOR2_X1 U445 ( .A(G43GAT), .B(G29GAT), .ZN(n372) );
  XNOR2_X1 U446 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U447 ( .A(KEYINPUT7), .B(n374), .Z(n392) );
  XNOR2_X1 U448 ( .A(G99GAT), .B(G106GAT), .ZN(n377) );
  XNOR2_X1 U449 ( .A(n293), .B(n377), .ZN(n406) );
  XOR2_X1 U450 ( .A(KEYINPUT9), .B(KEYINPUT79), .Z(n378) );
  XNOR2_X1 U451 ( .A(n381), .B(G134GAT), .ZN(n382) );
  XNOR2_X1 U452 ( .A(n385), .B(n384), .ZN(n560) );
  XOR2_X1 U453 ( .A(KEYINPUT29), .B(KEYINPUT64), .Z(n387) );
  NAND2_X1 U454 ( .A1(G229GAT), .A2(G233GAT), .ZN(n386) );
  XNOR2_X1 U455 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U456 ( .A(n388), .B(KEYINPUT30), .Z(n394) );
  XOR2_X1 U457 ( .A(KEYINPUT66), .B(G113GAT), .Z(n390) );
  XNOR2_X1 U458 ( .A(G36GAT), .B(G197GAT), .ZN(n389) );
  XNOR2_X1 U459 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U460 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U461 ( .A(n394), .B(n393), .ZN(n396) );
  XOR2_X1 U462 ( .A(n396), .B(n395), .Z(n400) );
  XNOR2_X1 U463 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U464 ( .A(n400), .B(n399), .ZN(n571) );
  XOR2_X1 U465 ( .A(KEYINPUT32), .B(KEYINPUT71), .Z(n402) );
  XNOR2_X1 U466 ( .A(G204GAT), .B(G92GAT), .ZN(n401) );
  XNOR2_X1 U467 ( .A(n402), .B(n401), .ZN(n417) );
  XOR2_X1 U468 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n404) );
  NAND2_X1 U469 ( .A1(G230GAT), .A2(G233GAT), .ZN(n403) );
  XNOR2_X1 U470 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U471 ( .A(n405), .B(KEYINPUT70), .Z(n409) );
  XNOR2_X1 U472 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U473 ( .A(n409), .B(n408), .ZN(n415) );
  XOR2_X1 U474 ( .A(G120GAT), .B(G71GAT), .Z(n433) );
  XNOR2_X1 U475 ( .A(n433), .B(n410), .ZN(n413) );
  XOR2_X1 U476 ( .A(n417), .B(n416), .Z(n577) );
  XOR2_X1 U477 ( .A(KEYINPUT41), .B(n577), .Z(n554) );
  NAND2_X1 U478 ( .A1(n571), .A2(n554), .ZN(n418) );
  XNOR2_X1 U479 ( .A(KEYINPUT46), .B(n418), .ZN(n419) );
  NAND2_X1 U480 ( .A1(n419), .A2(n567), .ZN(n420) );
  NOR2_X1 U481 ( .A1(n560), .A2(n420), .ZN(n421) );
  XNOR2_X1 U482 ( .A(n421), .B(KEYINPUT47), .ZN(n425) );
  XNOR2_X1 U483 ( .A(KEYINPUT81), .B(n560), .ZN(n466) );
  XNOR2_X1 U484 ( .A(KEYINPUT36), .B(n466), .ZN(n587) );
  NOR2_X1 U485 ( .A1(n587), .A2(n567), .ZN(n422) );
  NOR2_X1 U486 ( .A1(n292), .A2(n577), .ZN(n423) );
  XNOR2_X1 U487 ( .A(n571), .B(KEYINPUT67), .ZN(n563) );
  NAND2_X1 U488 ( .A1(n423), .A2(n563), .ZN(n424) );
  NAND2_X1 U489 ( .A1(n425), .A2(n424), .ZN(n427) );
  XOR2_X1 U490 ( .A(KEYINPUT112), .B(KEYINPUT48), .Z(n426) );
  XNOR2_X1 U491 ( .A(n427), .B(n426), .ZN(n454) );
  NOR2_X1 U492 ( .A1(n532), .A2(n454), .ZN(n428) );
  NAND2_X1 U493 ( .A1(n479), .A2(n428), .ZN(n429) );
  XNOR2_X1 U494 ( .A(KEYINPUT113), .B(n429), .ZN(n551) );
  XOR2_X1 U495 ( .A(G99GAT), .B(G190GAT), .Z(n431) );
  XNOR2_X1 U496 ( .A(G43GAT), .B(G15GAT), .ZN(n430) );
  XNOR2_X1 U497 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U498 ( .A(n433), .B(n432), .Z(n435) );
  NAND2_X1 U499 ( .A1(G227GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U500 ( .A(n435), .B(n434), .ZN(n447) );
  XOR2_X1 U501 ( .A(KEYINPUT89), .B(G176GAT), .Z(n437) );
  XNOR2_X1 U502 ( .A(G169GAT), .B(KEYINPUT20), .ZN(n436) );
  XNOR2_X1 U503 ( .A(n437), .B(n436), .ZN(n441) );
  XOR2_X1 U504 ( .A(KEYINPUT87), .B(KEYINPUT85), .Z(n439) );
  XNOR2_X1 U505 ( .A(KEYINPUT86), .B(KEYINPUT88), .ZN(n438) );
  XNOR2_X1 U506 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U507 ( .A(n441), .B(n440), .Z(n445) );
  XNOR2_X1 U508 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U509 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U510 ( .A(n447), .B(n446), .Z(n536) );
  INV_X1 U511 ( .A(n536), .ZN(n492) );
  NAND2_X1 U512 ( .A1(n551), .A2(n492), .ZN(n448) );
  XOR2_X1 U513 ( .A(KEYINPUT114), .B(n449), .Z(n548) );
  NOR2_X1 U514 ( .A1(n567), .A2(n548), .ZN(n452) );
  XNOR2_X1 U515 ( .A(n452), .B(n451), .ZN(G1342GAT) );
  INV_X1 U516 ( .A(n532), .ZN(n512) );
  XOR2_X1 U517 ( .A(n534), .B(KEYINPUT117), .Z(n453) );
  NOR2_X1 U518 ( .A1(n454), .A2(n453), .ZN(n457) );
  NOR2_X1 U519 ( .A1(n512), .A2(n458), .ZN(n570) );
  NAND2_X1 U520 ( .A1(n570), .A2(n476), .ZN(n460) );
  XOR2_X1 U521 ( .A(KEYINPUT55), .B(KEYINPUT119), .Z(n459) );
  XNOR2_X1 U522 ( .A(n460), .B(n459), .ZN(n461) );
  NAND2_X1 U523 ( .A1(n492), .A2(n461), .ZN(n462) );
  XNOR2_X1 U524 ( .A(n462), .B(KEYINPUT120), .ZN(n566) );
  INV_X1 U525 ( .A(n554), .ZN(n545) );
  NOR2_X1 U526 ( .A1(n566), .A2(n545), .ZN(n465) );
  XNOR2_X1 U527 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n463) );
  XNOR2_X1 U528 ( .A(n463), .B(G176GAT), .ZN(n464) );
  XNOR2_X1 U529 ( .A(n465), .B(n464), .ZN(G1349GAT) );
  NOR2_X1 U530 ( .A1(n566), .A2(n466), .ZN(n470) );
  XNOR2_X1 U531 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n468) );
  INV_X1 U532 ( .A(G190GAT), .ZN(n467) );
  NOR2_X1 U533 ( .A1(n492), .A2(n518), .ZN(n471) );
  NAND2_X1 U534 ( .A1(n479), .A2(n471), .ZN(n472) );
  NOR2_X1 U535 ( .A1(n532), .A2(n472), .ZN(n473) );
  XNOR2_X1 U536 ( .A(n473), .B(KEYINPUT97), .ZN(n484) );
  INV_X1 U537 ( .A(n534), .ZN(n515) );
  NAND2_X1 U538 ( .A1(n515), .A2(n492), .ZN(n474) );
  NAND2_X1 U539 ( .A1(n476), .A2(n474), .ZN(n475) );
  XOR2_X1 U540 ( .A(KEYINPUT25), .B(n475), .Z(n481) );
  NOR2_X1 U541 ( .A1(n492), .A2(n476), .ZN(n478) );
  XNOR2_X1 U542 ( .A(KEYINPUT98), .B(KEYINPUT26), .ZN(n477) );
  XNOR2_X1 U543 ( .A(n478), .B(n477), .ZN(n569) );
  NAND2_X1 U544 ( .A1(n479), .A2(n569), .ZN(n480) );
  NAND2_X1 U545 ( .A1(n481), .A2(n480), .ZN(n482) );
  NAND2_X1 U546 ( .A1(n532), .A2(n482), .ZN(n483) );
  NAND2_X1 U547 ( .A1(n484), .A2(n483), .ZN(n485) );
  XOR2_X1 U548 ( .A(KEYINPUT99), .B(n485), .Z(n499) );
  NAND2_X1 U549 ( .A1(n499), .A2(n567), .ZN(n486) );
  XNOR2_X1 U550 ( .A(n486), .B(KEYINPUT104), .ZN(n487) );
  NOR2_X1 U551 ( .A1(n587), .A2(n487), .ZN(n490) );
  XNOR2_X1 U552 ( .A(KEYINPUT106), .B(KEYINPUT37), .ZN(n488) );
  NOR2_X1 U553 ( .A1(n577), .A2(n563), .ZN(n500) );
  NAND2_X1 U554 ( .A1(n530), .A2(n500), .ZN(n491) );
  XOR2_X1 U555 ( .A(KEYINPUT38), .B(n491), .Z(n519) );
  NAND2_X1 U556 ( .A1(n519), .A2(n492), .ZN(n496) );
  XOR2_X1 U557 ( .A(KEYINPUT108), .B(KEYINPUT40), .Z(n494) );
  NAND2_X1 U558 ( .A1(n466), .A2(n581), .ZN(n497) );
  XOR2_X1 U559 ( .A(KEYINPUT16), .B(n497), .Z(n498) );
  AND2_X1 U560 ( .A1(n499), .A2(n498), .ZN(n521) );
  NAND2_X1 U561 ( .A1(n500), .A2(n521), .ZN(n509) );
  NOR2_X1 U562 ( .A1(n532), .A2(n509), .ZN(n502) );
  XNOR2_X1 U563 ( .A(KEYINPUT100), .B(KEYINPUT34), .ZN(n501) );
  XNOR2_X1 U564 ( .A(n502), .B(n501), .ZN(n503) );
  XOR2_X1 U565 ( .A(G1GAT), .B(n503), .Z(G1324GAT) );
  NOR2_X1 U566 ( .A1(n534), .A2(n509), .ZN(n504) );
  XOR2_X1 U567 ( .A(G8GAT), .B(n504), .Z(G1325GAT) );
  NOR2_X1 U568 ( .A1(n509), .A2(n536), .ZN(n508) );
  XOR2_X1 U569 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n506) );
  XNOR2_X1 U570 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n505) );
  XNOR2_X1 U571 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U572 ( .A(n508), .B(n507), .ZN(G1326GAT) );
  NOR2_X1 U573 ( .A1(n541), .A2(n509), .ZN(n511) );
  XNOR2_X1 U574 ( .A(G22GAT), .B(KEYINPUT103), .ZN(n510) );
  XNOR2_X1 U575 ( .A(n511), .B(n510), .ZN(G1327GAT) );
  NAND2_X1 U576 ( .A1(n512), .A2(n519), .ZN(n514) );
  XOR2_X1 U577 ( .A(G29GAT), .B(KEYINPUT39), .Z(n513) );
  XNOR2_X1 U578 ( .A(n514), .B(n513), .ZN(G1328GAT) );
  XOR2_X1 U579 ( .A(G36GAT), .B(KEYINPUT107), .Z(n517) );
  NAND2_X1 U580 ( .A1(n515), .A2(n519), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n517), .B(n516), .ZN(G1329GAT) );
  NAND2_X1 U582 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U583 ( .A(n520), .B(G50GAT), .ZN(G1331GAT) );
  NOR2_X1 U584 ( .A1(n571), .A2(n545), .ZN(n531) );
  NAND2_X1 U585 ( .A1(n531), .A2(n521), .ZN(n526) );
  NOR2_X1 U586 ( .A1(n532), .A2(n526), .ZN(n522) );
  XOR2_X1 U587 ( .A(G57GAT), .B(n522), .Z(n523) );
  XNOR2_X1 U588 ( .A(KEYINPUT42), .B(n523), .ZN(G1332GAT) );
  NOR2_X1 U589 ( .A1(n534), .A2(n526), .ZN(n524) );
  XOR2_X1 U590 ( .A(G64GAT), .B(n524), .Z(G1333GAT) );
  NOR2_X1 U591 ( .A1(n536), .A2(n526), .ZN(n525) );
  XOR2_X1 U592 ( .A(G71GAT), .B(n525), .Z(G1334GAT) );
  NOR2_X1 U593 ( .A1(n541), .A2(n526), .ZN(n528) );
  XNOR2_X1 U594 ( .A(KEYINPUT43), .B(KEYINPUT109), .ZN(n527) );
  XNOR2_X1 U595 ( .A(n528), .B(n527), .ZN(n529) );
  XOR2_X1 U596 ( .A(G78GAT), .B(n529), .Z(G1335GAT) );
  NAND2_X1 U597 ( .A1(n531), .A2(n530), .ZN(n540) );
  NOR2_X1 U598 ( .A1(n532), .A2(n540), .ZN(n533) );
  XOR2_X1 U599 ( .A(G85GAT), .B(n533), .Z(G1336GAT) );
  NOR2_X1 U600 ( .A1(n534), .A2(n540), .ZN(n535) );
  XOR2_X1 U601 ( .A(G92GAT), .B(n535), .Z(G1337GAT) );
  NOR2_X1 U602 ( .A1(n536), .A2(n540), .ZN(n538) );
  XNOR2_X1 U603 ( .A(KEYINPUT110), .B(KEYINPUT111), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U605 ( .A(G99GAT), .B(n539), .ZN(G1338GAT) );
  NOR2_X1 U606 ( .A1(n541), .A2(n540), .ZN(n542) );
  XOR2_X1 U607 ( .A(G106GAT), .B(n542), .Z(n543) );
  XNOR2_X1 U608 ( .A(KEYINPUT44), .B(n543), .ZN(G1339GAT) );
  NOR2_X1 U609 ( .A1(n548), .A2(n563), .ZN(n544) );
  XOR2_X1 U610 ( .A(G113GAT), .B(n544), .Z(G1340GAT) );
  NOR2_X1 U611 ( .A1(n548), .A2(n545), .ZN(n547) );
  XNOR2_X1 U612 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(G1341GAT) );
  NOR2_X1 U614 ( .A1(n548), .A2(n466), .ZN(n550) );
  XNOR2_X1 U615 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(G1343GAT) );
  XOR2_X1 U617 ( .A(G141GAT), .B(KEYINPUT115), .Z(n553) );
  AND2_X1 U618 ( .A1(n569), .A2(n551), .ZN(n561) );
  NAND2_X1 U619 ( .A1(n561), .A2(n571), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(G1344GAT) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(KEYINPUT116), .ZN(n558) );
  XOR2_X1 U622 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n556) );
  NAND2_X1 U623 ( .A1(n561), .A2(n554), .ZN(n555) );
  XNOR2_X1 U624 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(G1345GAT) );
  NAND2_X1 U626 ( .A1(n581), .A2(n561), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n559), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U628 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n562), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U630 ( .A1(n566), .A2(n563), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n564), .B(G169GAT), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n565), .B(KEYINPUT121), .ZN(G1348GAT) );
  NOR2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U634 ( .A(G183GAT), .B(n568), .Z(G1350GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT124), .B(KEYINPUT60), .Z(n573) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n586) );
  INV_X1 U637 ( .A(n586), .ZN(n582) );
  NAND2_X1 U638 ( .A1(n582), .A2(n571), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(n574) );
  XOR2_X1 U640 ( .A(n574), .B(KEYINPUT59), .Z(n576) );
  XNOR2_X1 U641 ( .A(G197GAT), .B(KEYINPUT123), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(G1352GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n579) );
  NAND2_X1 U644 ( .A1(n582), .A2(n577), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(n580) );
  XOR2_X1 U646 ( .A(G204GAT), .B(n580), .Z(G1353GAT) );
  XOR2_X1 U647 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n584) );
  NAND2_X1 U648 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U650 ( .A(G211GAT), .B(n585), .ZN(G1354GAT) );
  NOR2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U652 ( .A(KEYINPUT62), .B(n588), .Z(n589) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(n589), .ZN(G1355GAT) );
endmodule

