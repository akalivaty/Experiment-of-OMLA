//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 0 1 1 1 0 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 1 1 0 1 0 1 0 0 0 0 0 0 1 1 0 0 1 0 1 1 1 1 1 1 0 0 1 0 1 0 1 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:33 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1310, new_n1311, new_n1312, new_n1313, new_n1314,
    new_n1315, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1381, new_n1382, new_n1383,
    new_n1384, new_n1385, new_n1386, new_n1387, new_n1388, new_n1389;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT64), .Z(new_n210));
  AOI22_X1  g0010(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n214));
  NAND4_X1  g0014(.A1(new_n211), .A2(new_n212), .A3(new_n213), .A4(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n210), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT1), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n210), .A2(G13), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT0), .Z(new_n220));
  XNOR2_X1  g0020(.A(KEYINPUT65), .B(G20), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(new_n201), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(G50), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  AOI211_X1 g0026(.A(new_n217), .B(new_n220), .C1(new_n223), .C2(new_n226), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n231), .B(new_n234), .Z(G358));
  XOR2_X1   g0035(.A(G87), .B(G97), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT66), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  NAND2_X1  g0043(.A1(G33), .A2(G41), .ZN(new_n244));
  NAND3_X1  g0044(.A1(new_n244), .A2(G1), .A3(G13), .ZN(new_n245));
  INV_X1    g0045(.A(new_n245), .ZN(new_n246));
  OR2_X1    g0046(.A1(KEYINPUT3), .A2(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(KEYINPUT3), .A2(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  OAI21_X1  g0049(.A(new_n246), .B1(new_n249), .B2(G77), .ZN(new_n250));
  OR2_X1    g0050(.A1(G222), .A2(G1698), .ZN(new_n251));
  XNOR2_X1  g0051(.A(KEYINPUT68), .B(G223), .ZN(new_n252));
  INV_X1    g0052(.A(G1698), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n251), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n250), .B1(new_n249), .B2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G41), .ZN(new_n256));
  INV_X1    g0056(.A(G45), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G1), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT67), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT67), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G1), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n258), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n263), .A2(G226), .A3(new_n245), .ZN(new_n264));
  INV_X1    g0064(.A(G274), .ZN(new_n265));
  AND2_X1   g0065(.A1(G1), .A2(G13), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n265), .B1(new_n266), .B2(new_n244), .ZN(new_n267));
  AOI21_X1  g0067(.A(G1), .B1(new_n256), .B2(new_n257), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n264), .A2(new_n269), .ZN(new_n270));
  OR2_X1    g0070(.A1(new_n255), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G169), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(new_n222), .ZN(new_n275));
  OR2_X1    g0075(.A1(KEYINPUT8), .A2(G58), .ZN(new_n276));
  AND2_X1   g0076(.A1(KEYINPUT69), .A2(G58), .ZN(new_n277));
  NOR2_X1   g0077(.A1(KEYINPUT69), .A2(G58), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT8), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n276), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n221), .A2(G33), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n203), .A2(G20), .ZN(new_n284));
  OAI21_X1  g0084(.A(KEYINPUT70), .B1(G20), .B2(G33), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NOR3_X1   g0086(.A1(KEYINPUT70), .A2(G20), .A3(G33), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G150), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n284), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n275), .B1(new_n283), .B2(new_n290), .ZN(new_n291));
  XNOR2_X1  g0091(.A(KEYINPUT67), .B(G1), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n275), .B1(new_n292), .B2(G20), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G50), .ZN(new_n294));
  AND4_X1   g0094(.A1(G13), .A2(new_n260), .A3(new_n262), .A4(G20), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(new_n202), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n291), .A2(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n255), .A2(new_n270), .ZN(new_n299));
  INV_X1    g0099(.A(G179), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AND3_X1   g0101(.A1(new_n273), .A2(new_n298), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n298), .A2(KEYINPUT9), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT9), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n291), .A2(new_n304), .A3(new_n297), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n271), .A2(G200), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n299), .A2(G190), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n307), .A2(KEYINPUT72), .A3(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(KEYINPUT10), .B1(new_n306), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n303), .A2(new_n305), .ZN(new_n311));
  AND2_X1   g0111(.A1(new_n308), .A2(KEYINPUT72), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT10), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n311), .A2(new_n312), .A3(new_n313), .A4(new_n307), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n302), .B1(new_n310), .B2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT13), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n263), .A2(G238), .A3(new_n245), .ZN(new_n317));
  INV_X1    g0117(.A(G33), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n318), .A2(new_n205), .ZN(new_n319));
  NOR2_X1   g0119(.A1(G226), .A2(G1698), .ZN(new_n320));
  INV_X1    g0120(.A(G232), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n320), .B1(new_n321), .B2(G1698), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n319), .B1(new_n322), .B2(new_n249), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n269), .B(new_n317), .C1(new_n323), .C2(new_n245), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT73), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n316), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  AND3_X1   g0126(.A1(new_n268), .A2(new_n245), .A3(G274), .ZN(new_n327));
  INV_X1    g0127(.A(new_n319), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n321), .A2(G1698), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n329), .B1(G226), .B2(G1698), .ZN(new_n330));
  AND2_X1   g0130(.A1(KEYINPUT3), .A2(G33), .ZN(new_n331));
  NOR2_X1   g0131(.A1(KEYINPUT3), .A2(G33), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n328), .B1(new_n330), .B2(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n327), .B1(new_n334), .B2(new_n246), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n335), .A2(KEYINPUT73), .A3(new_n317), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n326), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n334), .A2(new_n246), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n338), .A2(new_n316), .A3(new_n269), .A4(new_n317), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n337), .A2(G179), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n324), .A2(KEYINPUT13), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(new_n339), .ZN(new_n342));
  AOI21_X1  g0142(.A(KEYINPUT14), .B1(new_n342), .B2(G169), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT14), .ZN(new_n344));
  AOI211_X1 g0144(.A(new_n344), .B(new_n272), .C1(new_n341), .C2(new_n339), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n340), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n221), .A2(G33), .A3(G77), .ZN(new_n347));
  OAI21_X1  g0147(.A(G50), .B1(new_n286), .B2(new_n287), .ZN(new_n348));
  INV_X1    g0148(.A(G68), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(G20), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n347), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n275), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT11), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n351), .A2(KEYINPUT11), .A3(new_n275), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n292), .A2(G13), .A3(G20), .ZN(new_n356));
  OAI21_X1  g0156(.A(KEYINPUT12), .B1(new_n356), .B2(G68), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT12), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n295), .A2(new_n358), .A3(new_n349), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n357), .A2(new_n359), .B1(G68), .B2(new_n293), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n354), .A2(new_n355), .A3(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n337), .A2(G190), .A3(new_n339), .ZN(new_n362));
  INV_X1    g0162(.A(G200), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n363), .B1(new_n341), .B2(new_n339), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n364), .A2(new_n361), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n346), .A2(new_n361), .B1(new_n362), .B2(new_n365), .ZN(new_n366));
  NOR2_X1   g0166(.A1(G232), .A2(G1698), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n253), .A2(G238), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n249), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n369), .B(new_n246), .C1(G107), .C2(new_n249), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n263), .A2(G244), .A3(new_n245), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n370), .A2(new_n269), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n272), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n373), .B1(G179), .B2(new_n372), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n293), .A2(G77), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(G77), .B2(new_n356), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT71), .ZN(new_n377));
  XNOR2_X1  g0177(.A(KEYINPUT15), .B(G87), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n377), .B1(new_n282), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n378), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n380), .A2(KEYINPUT71), .A3(G33), .A4(new_n221), .ZN(new_n381));
  OR3_X1    g0181(.A1(KEYINPUT70), .A2(G20), .A3(G33), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n285), .ZN(new_n383));
  XOR2_X1   g0183(.A(KEYINPUT8), .B(G58), .Z(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(G20), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(KEYINPUT65), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT65), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(G20), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(G77), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n379), .A2(new_n381), .A3(new_n385), .A4(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n376), .B1(new_n392), .B2(new_n275), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n374), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(G190), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n372), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n396), .B1(G200), .B2(new_n372), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n394), .B1(new_n393), .B2(new_n397), .ZN(new_n398));
  AND3_X1   g0198(.A1(new_n315), .A2(new_n366), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n321), .B1(new_n266), .B2(new_n244), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n263), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT75), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n401), .A2(new_n269), .A3(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n402), .B1(new_n401), .B2(new_n269), .ZN(new_n405));
  INV_X1    g0205(.A(G223), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n253), .ZN(new_n407));
  INV_X1    g0207(.A(G226), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(G1698), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n407), .B(new_n409), .C1(new_n331), .C2(new_n332), .ZN(new_n410));
  NAND2_X1  g0210(.A1(G33), .A2(G87), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n245), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NOR4_X1   g0212(.A1(new_n404), .A2(new_n405), .A3(G179), .A4(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n401), .A2(new_n269), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n412), .B1(new_n414), .B2(KEYINPUT75), .ZN(new_n415));
  AOI21_X1  g0215(.A(G169), .B1(new_n415), .B2(new_n403), .ZN(new_n416));
  OAI21_X1  g0216(.A(KEYINPUT76), .B1(new_n413), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n281), .A2(new_n356), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(new_n281), .B2(new_n293), .ZN(new_n419));
  OAI21_X1  g0219(.A(G68), .B1(new_n277), .B2(new_n278), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n224), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n421), .A2(G20), .B1(new_n383), .B2(G159), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT7), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n333), .A2(new_n221), .A3(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n247), .A2(new_n386), .A3(new_n248), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT7), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n424), .A2(new_n426), .A3(G68), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n422), .A2(new_n427), .A3(KEYINPUT16), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n275), .ZN(new_n429));
  XNOR2_X1  g0229(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n333), .A2(new_n423), .A3(new_n386), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n249), .A2(new_n390), .ZN(new_n433));
  OAI211_X1 g0233(.A(G68), .B(new_n432), .C1(new_n433), .C2(new_n423), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n431), .B1(new_n434), .B2(new_n422), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n419), .B1(new_n429), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n415), .A2(new_n300), .A3(new_n403), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT76), .ZN(new_n438));
  NOR3_X1   g0238(.A1(new_n404), .A2(new_n405), .A3(new_n412), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n437), .B(new_n438), .C1(new_n439), .C2(G169), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n417), .A2(new_n436), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(KEYINPUT18), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT18), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n417), .A2(new_n443), .A3(new_n440), .A4(new_n436), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n415), .A2(new_n395), .A3(new_n403), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n445), .B1(new_n439), .B2(G200), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n434), .A2(new_n422), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n430), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n448), .A2(new_n275), .A3(new_n428), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n446), .A2(new_n449), .A3(new_n419), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT17), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n446), .A2(new_n449), .A3(KEYINPUT17), .A4(new_n419), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n442), .A2(new_n444), .A3(new_n452), .A4(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n399), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n387), .A2(new_n389), .A3(G33), .A4(G97), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT19), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n249), .A2(new_n221), .A3(G68), .ZN(new_n460));
  NAND3_X1  g0260(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n387), .A2(new_n389), .A3(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(G97), .A2(G107), .ZN(new_n463));
  INV_X1    g0263(.A(G87), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n459), .A2(new_n460), .A3(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT81), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n459), .A2(new_n460), .A3(new_n466), .A4(KEYINPUT81), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n469), .A2(new_n275), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n295), .A2(new_n378), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT78), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n260), .A2(new_n262), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n473), .B1(new_n474), .B2(new_n318), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n292), .A2(KEYINPUT78), .A3(G33), .ZN(new_n476));
  INV_X1    g0276(.A(new_n275), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n475), .A2(new_n356), .A3(new_n476), .A4(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(G87), .ZN(new_n480));
  AND3_X1   g0280(.A1(new_n471), .A2(new_n472), .A3(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n260), .A2(new_n262), .A3(G45), .ZN(new_n482));
  INV_X1    g0282(.A(G250), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n483), .B1(new_n266), .B2(new_n244), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(KEYINPUT80), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT80), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n482), .A2(new_n484), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(G33), .A2(G116), .ZN(new_n490));
  INV_X1    g0290(.A(G244), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(G1698), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n492), .B1(G238), .B2(G1698), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n490), .B1(new_n493), .B2(new_n333), .ZN(new_n494));
  AND3_X1   g0294(.A1(new_n260), .A2(new_n262), .A3(G45), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n494), .A2(new_n246), .B1(new_n267), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n489), .A2(new_n496), .A3(new_n395), .ZN(new_n497));
  INV_X1    g0297(.A(new_n488), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n487), .B1(new_n482), .B2(new_n484), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n495), .A2(new_n267), .ZN(new_n501));
  INV_X1    g0301(.A(new_n490), .ZN(new_n502));
  NOR2_X1   g0302(.A1(G238), .A2(G1698), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n503), .B1(new_n491), .B2(G1698), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n502), .B1(new_n504), .B2(new_n249), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n501), .B1(new_n505), .B2(new_n245), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n500), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n497), .B1(new_n507), .B2(G200), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n481), .A2(new_n508), .ZN(new_n509));
  NOR3_X1   g0309(.A1(new_n500), .A2(new_n506), .A3(G179), .ZN(new_n510));
  AOI21_X1  g0310(.A(G169), .B1(new_n489), .B2(new_n496), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n479), .A2(new_n380), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n471), .A2(new_n513), .A3(new_n472), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n509), .A2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(G77), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n288), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G97), .A2(G107), .ZN(new_n519));
  AND2_X1   g0319(.A1(KEYINPUT6), .A2(G107), .ZN(new_n520));
  NOR2_X1   g0320(.A1(KEYINPUT77), .A2(KEYINPUT6), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n207), .B(new_n519), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n519), .ZN(new_n523));
  OAI22_X1  g0323(.A1(new_n523), .A2(new_n463), .B1(KEYINPUT77), .B2(KEYINPUT6), .ZN(new_n524));
  AND2_X1   g0324(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n518), .B1(new_n525), .B2(new_n390), .ZN(new_n526));
  OAI211_X1 g0326(.A(G107), .B(new_n432), .C1(new_n433), .C2(new_n423), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n477), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n295), .A2(new_n205), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n529), .B1(new_n478), .B2(new_n205), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n491), .A2(G1698), .ZN(new_n532));
  AOI21_X1  g0332(.A(KEYINPUT4), .B1(new_n249), .B2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(G250), .A2(G1698), .ZN(new_n535));
  NAND2_X1  g0335(.A1(KEYINPUT4), .A2(G244), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n535), .B1(new_n536), .B2(G1698), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n249), .A2(new_n537), .B1(G33), .B2(G283), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n245), .B1(new_n534), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n256), .A2(KEYINPUT5), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT5), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(G41), .ZN(new_n542));
  AND2_X1   g0342(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n495), .A2(new_n267), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n540), .A2(new_n542), .ZN(new_n545));
  OAI211_X1 g0345(.A(G257), .B(new_n245), .C1(new_n482), .C2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n539), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n548), .A2(KEYINPUT79), .A3(G190), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT79), .ZN(new_n550));
  AND2_X1   g0350(.A1(new_n544), .A2(new_n546), .ZN(new_n551));
  NAND2_X1  g0351(.A1(G33), .A2(G283), .ZN(new_n552));
  INV_X1    g0352(.A(new_n537), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n552), .B1(new_n553), .B2(new_n333), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n246), .B1(new_n554), .B2(new_n533), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n550), .B1(new_n556), .B2(new_n395), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(G200), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n531), .A2(new_n549), .A3(new_n557), .A4(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n551), .A2(new_n555), .A3(new_n300), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n272), .B1(new_n539), .B2(new_n547), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n560), .B(new_n561), .C1(new_n528), .C2(new_n530), .ZN(new_n562));
  AND2_X1   g0362(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT25), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(new_n356), .B2(G107), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n295), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n479), .A2(G107), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  OAI211_X1 g0368(.A(G264), .B(new_n245), .C1(new_n482), .C2(new_n545), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n483), .A2(new_n253), .ZN(new_n570));
  INV_X1    g0370(.A(G257), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(G1698), .ZN(new_n572));
  AND2_X1   g0372(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n573), .A2(new_n249), .B1(G33), .B2(G294), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n569), .B(new_n544), .C1(new_n574), .C2(new_n245), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n363), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(G190), .B2(new_n575), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT82), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT23), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n390), .A2(new_n578), .A3(new_n579), .A4(new_n206), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n206), .ZN(new_n581));
  OAI21_X1  g0381(.A(KEYINPUT82), .B1(new_n221), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n249), .A2(new_n221), .A3(KEYINPUT22), .A4(G87), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n249), .A2(new_n221), .A3(G87), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT22), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n206), .A2(G20), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(KEYINPUT23), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n590), .B1(G20), .B2(new_n490), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g0393(.A(KEYINPUT24), .B1(new_n585), .B2(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n591), .B1(new_n586), .B2(new_n587), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT24), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n595), .A2(new_n583), .A3(new_n596), .A4(new_n584), .ZN(new_n597));
  AND2_X1   g0397(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n568), .B(new_n577), .C1(new_n598), .C2(new_n477), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n246), .B1(new_n495), .B2(new_n543), .ZN(new_n600));
  NAND2_X1  g0400(.A1(G33), .A2(G294), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n570), .A2(new_n572), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n601), .B1(new_n602), .B2(new_n333), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n600), .A2(G264), .B1(new_n603), .B2(new_n246), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n604), .A2(new_n300), .A3(new_n544), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n575), .A2(new_n272), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n477), .B1(new_n594), .B2(new_n597), .ZN(new_n607));
  INV_X1    g0407(.A(new_n568), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n605), .B(new_n606), .C1(new_n607), .C2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(G303), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n247), .A2(new_n610), .A3(new_n248), .ZN(new_n611));
  MUX2_X1   g0411(.A(G257), .B(G264), .S(G1698), .Z(new_n612));
  OAI211_X1 g0412(.A(new_n246), .B(new_n611), .C1(new_n612), .C2(new_n333), .ZN(new_n613));
  OAI211_X1 g0413(.A(G270), .B(new_n245), .C1(new_n482), .C2(new_n545), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n613), .A2(new_n544), .A3(new_n614), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n615), .A2(G169), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n318), .A2(G97), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n221), .A2(new_n552), .A3(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(G116), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n274), .A2(new_n222), .B1(G20), .B2(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n618), .A2(KEYINPUT20), .A3(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(KEYINPUT20), .B1(new_n618), .B2(new_n620), .ZN(new_n623));
  OAI22_X1  g0423(.A1(new_n622), .A2(new_n623), .B1(G116), .B2(new_n356), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n478), .A2(new_n619), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n616), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT21), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n295), .A2(new_n619), .ZN(new_n628));
  OAI221_X1 g0428(.A(new_n628), .B1(new_n478), .B2(new_n619), .C1(new_n623), .C2(new_n622), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n615), .A2(KEYINPUT21), .A3(G169), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n544), .A2(new_n613), .A3(new_n614), .A4(G179), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n626), .A2(new_n627), .B1(new_n629), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n615), .A2(G200), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n634), .B1(new_n395), .B2(new_n615), .ZN(new_n635));
  OR2_X1    g0435(.A1(new_n635), .A2(new_n629), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n599), .A2(new_n609), .A3(new_n633), .A4(new_n636), .ZN(new_n637));
  NOR4_X1   g0437(.A1(new_n456), .A2(new_n516), .A3(new_n564), .A4(new_n637), .ZN(G372));
  NAND2_X1  g0438(.A1(new_n310), .A2(new_n314), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n452), .A2(new_n453), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n346), .A2(new_n361), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n362), .A2(new_n365), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n394), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n640), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n442), .A2(new_n444), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n639), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n302), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(KEYINPUT83), .B1(new_n507), .B2(G169), .ZN(new_n650));
  INV_X1    g0450(.A(new_n510), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT83), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n511), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n650), .A2(new_n514), .A3(new_n651), .A4(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n562), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(new_n509), .A3(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT26), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AOI22_X1  g0458(.A1(new_n481), .A2(new_n508), .B1(new_n512), .B2(new_n514), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n659), .A2(KEYINPUT26), .A3(new_n655), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n609), .A2(new_n633), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n563), .A2(new_n509), .A3(new_n662), .A4(new_n599), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n661), .A2(new_n663), .A3(new_n654), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n649), .B1(new_n456), .B2(new_n665), .ZN(G369));
  INV_X1    g0466(.A(KEYINPUT85), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT84), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n221), .A2(G13), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n668), .B1(new_n669), .B2(new_n474), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT27), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n221), .A2(new_n292), .A3(KEYINPUT84), .A4(G13), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(G213), .ZN(new_n674));
  INV_X1    g0474(.A(G343), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n671), .B1(new_n670), .B2(new_n672), .ZN(new_n676));
  NOR3_X1   g0476(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n629), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n633), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n633), .A2(new_n636), .A3(new_n678), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n667), .B1(new_n681), .B2(G330), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n681), .A2(new_n667), .A3(G330), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n599), .A2(new_n609), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n677), .B1(new_n607), .B2(new_n608), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n609), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n677), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n685), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n677), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n629), .A2(new_n632), .ZN(new_n695));
  AOI21_X1  g0495(.A(KEYINPUT21), .B1(new_n629), .B2(new_n616), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n694), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  OAI22_X1  g0497(.A1(new_n686), .A2(new_n697), .B1(new_n609), .B2(new_n677), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n693), .A2(new_n699), .ZN(G399));
  INV_X1    g0500(.A(new_n218), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(G41), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n465), .A2(G116), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NOR3_X1   g0504(.A1(new_n702), .A2(new_n259), .A3(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n705), .B1(new_n226), .B2(new_n702), .ZN(new_n706));
  XOR2_X1   g0506(.A(new_n706), .B(KEYINPUT28), .Z(new_n707));
  NAND4_X1  g0507(.A1(new_n659), .A2(new_n562), .A3(new_n559), .A4(new_n694), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT30), .ZN(new_n709));
  AND4_X1   g0509(.A1(G179), .A2(new_n613), .A3(new_n544), .A4(new_n614), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n710), .A2(new_n489), .A3(new_n604), .A4(new_n496), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n709), .B1(new_n711), .B2(new_n556), .ZN(new_n712));
  OAI211_X1 g0512(.A(new_n300), .B(new_n615), .C1(new_n500), .C2(new_n506), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n575), .B1(new_n539), .B2(new_n547), .ZN(new_n714));
  OR2_X1    g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n489), .A2(new_n496), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n569), .B1(new_n574), .B2(new_n245), .ZN(new_n717));
  NOR3_X1   g0517(.A1(new_n716), .A2(new_n717), .A3(new_n631), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n551), .A2(new_n555), .A3(KEYINPUT30), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n712), .A2(new_n715), .A3(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(KEYINPUT31), .B1(new_n722), .B2(new_n677), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT86), .ZN(new_n724));
  OAI22_X1  g0524(.A1(new_n637), .A2(new_n708), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(KEYINPUT30), .B1(new_n718), .B2(new_n548), .ZN(new_n726));
  OAI22_X1  g0526(.A1(new_n711), .A2(new_n719), .B1(new_n713), .B2(new_n714), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n677), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT31), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n722), .A2(KEYINPUT31), .A3(new_n677), .ZN(new_n731));
  AOI21_X1  g0531(.A(KEYINPUT86), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(G330), .B1(new_n725), .B2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  XNOR2_X1  g0534(.A(KEYINPUT88), .B(KEYINPUT29), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT87), .ZN(new_n737));
  AND3_X1   g0537(.A1(new_n664), .A2(new_n737), .A3(new_n694), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n737), .B1(new_n664), .B2(new_n694), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n736), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n654), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n599), .A2(new_n559), .A3(new_n509), .A4(new_n562), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n741), .B1(new_n743), .B2(new_n662), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n657), .B1(new_n516), .B2(new_n562), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n654), .A2(new_n509), .A3(new_n655), .A4(KEYINPUT26), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n677), .B1(new_n744), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(KEYINPUT29), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n734), .B1(new_n740), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n707), .B1(new_n750), .B2(G1), .ZN(G364));
  INV_X1    g0551(.A(KEYINPUT89), .ZN(new_n752));
  INV_X1    g0552(.A(new_n684), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n752), .B1(new_n753), .B2(new_n682), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n683), .A2(KEYINPUT89), .A3(new_n684), .ZN(new_n755));
  INV_X1    g0555(.A(new_n669), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n259), .B1(new_n756), .B2(G45), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n702), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(G330), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n679), .A2(new_n761), .A3(new_n680), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n754), .A2(new_n755), .A3(new_n760), .A4(new_n762), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n763), .B(KEYINPUT90), .ZN(new_n764));
  NOR4_X1   g0564(.A1(new_n386), .A2(new_n395), .A3(new_n363), .A4(G179), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n249), .B1(new_n765), .B2(G303), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n221), .A2(new_n300), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n767), .A2(G190), .A3(G200), .ZN(new_n768));
  INV_X1    g0568(.A(G326), .ZN(new_n769));
  NOR4_X1   g0569(.A1(new_n221), .A2(new_n300), .A3(G190), .A4(G200), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(G311), .ZN(new_n772));
  OAI221_X1 g0572(.A(new_n766), .B1(new_n768), .B2(new_n769), .C1(new_n771), .C2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n395), .A2(G200), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n221), .B1(new_n300), .B2(new_n774), .ZN(new_n775));
  OR2_X1    g0575(.A1(new_n775), .A2(KEYINPUT95), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(KEYINPUT95), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n773), .B1(G294), .B2(new_n779), .ZN(new_n780));
  NOR3_X1   g0580(.A1(new_n363), .A2(G179), .A3(G190), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n390), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR3_X1   g0583(.A1(G179), .A2(G190), .A3(G200), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n390), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI22_X1  g0586(.A1(G283), .A2(new_n783), .B1(new_n786), .B2(G329), .ZN(new_n787));
  XOR2_X1   g0587(.A(new_n787), .B(KEYINPUT96), .Z(new_n788));
  NAND3_X1  g0588(.A1(new_n767), .A2(new_n395), .A3(G200), .ZN(new_n789));
  XOR2_X1   g0589(.A(KEYINPUT33), .B(G317), .Z(new_n790));
  NAND2_X1  g0590(.A1(new_n767), .A2(new_n774), .ZN(new_n791));
  INV_X1    g0591(.A(G322), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n789), .A2(new_n790), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n793), .B(KEYINPUT97), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n780), .A2(new_n788), .A3(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(G159), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n785), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g0597(.A(KEYINPUT94), .B(KEYINPUT32), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n783), .A2(G107), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n333), .B1(new_n765), .B2(G87), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n202), .A2(new_n768), .B1(new_n789), .B2(new_n349), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n797), .A2(new_n798), .B1(new_n791), .B2(new_n279), .ZN(new_n804));
  NOR3_X1   g0604(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n779), .A2(G97), .ZN(new_n806));
  AND2_X1   g0606(.A1(new_n770), .A2(KEYINPUT93), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n770), .A2(KEYINPUT93), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n805), .B(new_n806), .C1(new_n517), .C2(new_n809), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n266), .B1(new_n386), .B2(G169), .ZN(new_n811));
  OR2_X1    g0611(.A1(new_n811), .A2(KEYINPUT92), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(KEYINPUT92), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n795), .A2(new_n810), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n812), .A2(new_n813), .ZN(new_n815));
  NOR2_X1   g0615(.A1(G13), .A2(G33), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n817), .A2(G20), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n701), .A2(new_n249), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n226), .A2(new_n257), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n820), .B(new_n821), .C1(new_n257), .C2(new_n242), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n218), .A2(new_n249), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT91), .ZN(new_n824));
  INV_X1    g0624(.A(G355), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n822), .B1(G116), .B2(new_n218), .C1(new_n824), .C2(new_n825), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n760), .B(new_n814), .C1(new_n819), .C2(new_n826), .ZN(new_n827));
  XOR2_X1   g0627(.A(new_n827), .B(KEYINPUT98), .Z(new_n828));
  INV_X1    g0628(.A(new_n818), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n828), .B1(new_n681), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n764), .A2(new_n830), .ZN(G396));
  NOR2_X1   g0631(.A1(new_n782), .A2(new_n464), .ZN(new_n832));
  INV_X1    g0632(.A(new_n765), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n333), .B1(new_n785), .B2(new_n772), .C1(new_n833), .C2(new_n206), .ZN(new_n834));
  INV_X1    g0634(.A(new_n791), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n832), .B(new_n834), .C1(G294), .C2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n809), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(G116), .ZN(new_n838));
  INV_X1    g0638(.A(new_n789), .ZN(new_n839));
  INV_X1    g0639(.A(new_n768), .ZN(new_n840));
  AOI22_X1  g0640(.A1(G283), .A2(new_n839), .B1(new_n840), .B2(G303), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n836), .A2(new_n838), .A3(new_n806), .A4(new_n841), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n840), .A2(G137), .B1(new_n835), .B2(G143), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n843), .B1(new_n289), .B2(new_n789), .C1(new_n809), .C2(new_n796), .ZN(new_n844));
  XOR2_X1   g0644(.A(new_n844), .B(KEYINPUT34), .Z(new_n845));
  OAI21_X1  g0645(.A(new_n249), .B1(new_n833), .B2(new_n202), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n846), .B1(G132), .B2(new_n786), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n782), .A2(new_n349), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n847), .B(new_n849), .C1(new_n279), .C2(new_n778), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n842), .B1(new_n845), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(new_n815), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n815), .A2(new_n816), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n852), .B(new_n759), .C1(G77), .C2(new_n854), .ZN(new_n855));
  OR2_X1    g0655(.A1(new_n374), .A2(new_n393), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n397), .A2(new_n393), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n856), .B(new_n857), .C1(new_n393), .C2(new_n694), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n394), .A2(KEYINPUT99), .A3(new_n677), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(KEYINPUT99), .B1(new_n394), .B2(new_n677), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n858), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n816), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n855), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT99), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n867), .B1(new_n856), .B2(new_n694), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(new_n859), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n677), .B1(new_n869), .B2(new_n858), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n664), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n738), .A2(new_n739), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n871), .B1(new_n872), .B2(new_n862), .ZN(new_n873));
  OR2_X1    g0673(.A1(new_n873), .A2(new_n733), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n759), .B1(new_n873), .B2(new_n733), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n866), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(G384));
  NAND2_X1  g0677(.A1(new_n394), .A2(new_n694), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n878), .B(KEYINPUT100), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n879), .B1(new_n664), .B2(new_n870), .ZN(new_n880));
  INV_X1    g0680(.A(new_n361), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n694), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n339), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n316), .B1(new_n335), .B2(new_n317), .ZN(new_n885));
  OAI21_X1  g0685(.A(G169), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n344), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n342), .A2(KEYINPUT14), .A3(G169), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n884), .B1(new_n326), .B2(new_n336), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n887), .A2(new_n888), .B1(G179), .B2(new_n889), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n642), .B(new_n883), .C1(new_n890), .C2(new_n881), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT101), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n366), .A2(KEYINPUT101), .A3(new_n883), .ZN(new_n894));
  AND2_X1   g0694(.A1(new_n362), .A2(new_n365), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n882), .B1(new_n895), .B2(new_n346), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(KEYINPUT102), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT102), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n898), .B(new_n882), .C1(new_n895), .C2(new_n346), .ZN(new_n899));
  AOI22_X1  g0699(.A1(new_n893), .A2(new_n894), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n880), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n431), .B1(new_n422), .B2(new_n427), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n419), .B1(new_n429), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n674), .A2(new_n676), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n454), .A2(new_n906), .ZN(new_n907));
  AND3_X1   g0707(.A1(new_n417), .A2(new_n440), .A3(new_n903), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n450), .A2(new_n905), .ZN(new_n909));
  OAI21_X1  g0709(.A(KEYINPUT37), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n436), .A2(new_n904), .ZN(new_n911));
  XOR2_X1   g0711(.A(KEYINPUT103), .B(KEYINPUT37), .Z(new_n912));
  NAND4_X1  g0712(.A1(new_n441), .A2(new_n450), .A3(new_n911), .A4(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n907), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT38), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI22_X1  g0717(.A1(new_n454), .A2(new_n906), .B1(new_n910), .B2(new_n913), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(KEYINPUT38), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n901), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n904), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n645), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n641), .A2(new_n677), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n441), .A2(new_n450), .A3(new_n911), .ZN(new_n927));
  INV_X1    g0727(.A(new_n912), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT104), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n929), .A2(new_n930), .A3(new_n913), .ZN(new_n931));
  INV_X1    g0731(.A(new_n911), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n454), .A2(new_n932), .ZN(new_n933));
  OR2_X1    g0733(.A1(new_n913), .A2(new_n930), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n931), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n916), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT39), .B1(new_n918), .B2(KEYINPUT38), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AND3_X1   g0738(.A1(new_n907), .A2(KEYINPUT38), .A3(new_n914), .ZN(new_n939));
  AOI21_X1  g0739(.A(KEYINPUT38), .B1(new_n907), .B2(new_n914), .ZN(new_n940));
  OAI21_X1  g0740(.A(KEYINPUT39), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n926), .B1(new_n938), .B2(new_n941), .ZN(new_n942));
  NOR3_X1   g0742(.A1(new_n924), .A2(new_n942), .A3(KEYINPUT105), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT105), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n938), .A2(new_n941), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n925), .ZN(new_n946));
  AOI22_X1  g0746(.A1(new_n901), .A2(new_n920), .B1(new_n645), .B2(new_n922), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n944), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n943), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n664), .A2(new_n694), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(KEYINPUT87), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n664), .A2(new_n737), .A3(new_n694), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n735), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n456), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n749), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n649), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n949), .B(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n936), .A2(new_n919), .ZN(new_n958));
  OAI211_X1 g0758(.A(new_n730), .B(new_n731), .C1(new_n708), .C2(new_n637), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n862), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n891), .A2(new_n892), .ZN(new_n962));
  AOI21_X1  g0762(.A(KEYINPUT101), .B1(new_n366), .B2(new_n883), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n890), .A2(new_n642), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n898), .B1(new_n964), .B2(new_n882), .ZN(new_n965));
  INV_X1    g0765(.A(new_n899), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n962), .A2(new_n963), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT106), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n961), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(KEYINPUT106), .B1(new_n900), .B2(new_n960), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n958), .A2(new_n969), .A3(new_n970), .A4(KEYINPUT40), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n961), .B(new_n967), .C1(new_n939), .C2(new_n940), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT40), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n954), .A2(new_n959), .ZN(new_n976));
  AND2_X1   g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n975), .A2(new_n976), .ZN(new_n978));
  NOR3_X1   g0778(.A1(new_n977), .A2(new_n978), .A3(new_n761), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  AOI22_X1  g0780(.A1(new_n957), .A2(new_n980), .B1(new_n474), .B2(new_n669), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n980), .B2(new_n957), .ZN(new_n982));
  INV_X1    g0782(.A(new_n525), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT35), .ZN(new_n984));
  OAI211_X1 g0784(.A(G116), .B(new_n223), .C1(new_n983), .C2(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(new_n984), .B2(new_n983), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT36), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n226), .A2(G77), .A3(new_n420), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n202), .A2(G68), .ZN(new_n989));
  AOI211_X1 g0789(.A(G13), .B(new_n292), .C1(new_n988), .C2(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n982), .A2(new_n991), .ZN(G367));
  AOI211_X1 g0792(.A(new_n818), .B(new_n815), .C1(new_n701), .C2(new_n380), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n820), .A2(new_n234), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n760), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(G317), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n333), .B1(new_n785), .B2(new_n996), .C1(new_n205), .C2(new_n782), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n765), .A2(G116), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n998), .B(KEYINPUT46), .Z(new_n999));
  AOI211_X1 g0799(.A(new_n997), .B(new_n999), .C1(G303), .C2(new_n835), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(G294), .A2(new_n839), .B1(new_n840), .B2(G311), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n837), .A2(G283), .B1(G107), .B2(new_n779), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n837), .A2(G50), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(KEYINPUT69), .B(G58), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n333), .B1(new_n765), .B2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n390), .A2(G77), .A3(new_n781), .ZN(new_n1007));
  INV_X1    g0807(.A(G137), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n1006), .B(new_n1007), .C1(new_n1008), .C2(new_n785), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(G150), .B2(new_n835), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(G143), .A2(new_n840), .B1(new_n839), .B2(G159), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n779), .A2(G68), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1004), .A2(new_n1010), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1003), .A2(KEYINPUT47), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n815), .ZN(new_n1015));
  AOI21_X1  g0815(.A(KEYINPUT47), .B1(new_n1003), .B2(new_n1013), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n471), .A2(new_n472), .A3(new_n480), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n677), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT107), .ZN(new_n1019));
  NOR3_X1   g0819(.A1(new_n654), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1019), .B1(new_n654), .B2(new_n1018), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n654), .A2(new_n509), .A3(new_n1018), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1020), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n995), .B1(new_n1015), .B2(new_n1016), .C1(new_n829), .C2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT112), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n740), .A2(new_n749), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(new_n733), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n677), .B1(new_n528), .B2(new_n530), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n559), .A2(new_n562), .A3(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n655), .A2(new_n677), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(KEYINPUT110), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT110), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1030), .A2(new_n1034), .A3(new_n1031), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1033), .A2(new_n698), .A3(new_n1035), .ZN(new_n1036));
  XOR2_X1   g0836(.A(KEYINPUT111), .B(KEYINPUT44), .Z(new_n1037));
  XNOR2_X1  g0837(.A(new_n1036), .B(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT45), .ZN(new_n1039));
  AND3_X1   g0839(.A1(new_n1030), .A2(new_n1034), .A3(new_n1031), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1034), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1039), .B1(new_n1042), .B2(new_n698), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1044), .A2(KEYINPUT45), .A3(new_n699), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  AND3_X1   g0846(.A1(new_n1038), .A2(new_n693), .A3(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n693), .B1(new_n1038), .B2(new_n1046), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n697), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n687), .A2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n692), .B2(new_n1050), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n754), .A2(new_n755), .A3(new_n1052), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n685), .B(new_n1051), .C1(new_n692), .C2(new_n1050), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1028), .B1(new_n1049), .B2(new_n1056), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n702), .B(KEYINPUT41), .Z(new_n1058));
  OAI21_X1  g0858(.A(new_n757), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(KEYINPUT42), .B1(new_n1042), .B2(new_n1051), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT42), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1044), .A2(new_n1061), .A3(new_n687), .A4(new_n1050), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n655), .B1(new_n1044), .B2(new_n690), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1060), .B(new_n1062), .C1(new_n1063), .C2(new_n677), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1024), .A2(KEYINPUT43), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1020), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1023), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1067), .B1(new_n1068), .B2(new_n1021), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT108), .ZN(new_n1070));
  AOI21_X1  g0870(.A(KEYINPUT43), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT109), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1024), .A2(KEYINPUT108), .ZN(new_n1073));
  AND3_X1   g0873(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1072), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1066), .A2(new_n1076), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1064), .B(new_n1065), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n693), .A2(new_n1042), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1077), .A2(new_n1080), .A3(new_n1078), .ZN(new_n1083));
  AND2_X1   g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1026), .B1(new_n1059), .B2(new_n1084), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n683), .A2(new_n684), .B1(new_n689), .B2(new_n691), .ZN(new_n1086));
  AND2_X1   g0886(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1037), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1036), .B(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1086), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1038), .A2(new_n693), .A3(new_n1046), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n750), .B1(new_n1092), .B2(new_n1055), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1058), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n758), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1096));
  NOR3_X1   g0896(.A1(new_n1095), .A2(new_n1096), .A3(KEYINPUT112), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1025), .B1(new_n1085), .B2(new_n1097), .ZN(G387));
  NAND2_X1  g0898(.A1(new_n1028), .A2(new_n1055), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1056), .A2(new_n750), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1099), .A2(new_n702), .A3(new_n1100), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n809), .A2(new_n610), .B1(new_n996), .B2(new_n791), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT114), .ZN(new_n1103));
  OR2_X1    g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(G311), .A2(new_n839), .B1(new_n840), .B2(G322), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT48), .ZN(new_n1108));
  OR2_X1    g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n779), .A2(G283), .B1(G294), .B2(new_n765), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1109), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  XOR2_X1   g0912(.A(new_n1112), .B(KEYINPUT49), .Z(new_n1113));
  OAI221_X1 g0913(.A(new_n333), .B1(new_n785), .B2(new_n769), .C1(new_n619), .C2(new_n782), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n796), .A2(new_n768), .B1(new_n789), .B2(new_n281), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n765), .A2(G77), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n249), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(G97), .B2(new_n783), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n835), .A2(G50), .B1(G68), .B2(new_n770), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1119), .B(new_n1120), .C1(new_n289), .C2(new_n785), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n1116), .B(new_n1121), .C1(new_n380), .C2(new_n779), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n815), .B1(new_n1115), .B2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n692), .A2(new_n829), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n257), .B1(new_n349), .B2(new_n517), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(new_n704), .B2(KEYINPUT113), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1126), .B1(KEYINPUT113), .B2(new_n704), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n384), .A2(new_n202), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(new_n1128), .B(KEYINPUT50), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n820), .B1(new_n1127), .B2(new_n1129), .C1(new_n231), .C2(new_n257), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n1130), .B1(G107), .B2(new_n218), .C1(new_n703), .C2(new_n824), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n760), .B(new_n1124), .C1(new_n819), .C2(new_n1131), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n1123), .A2(new_n1132), .B1(new_n1056), .B2(new_n758), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1101), .A2(new_n1133), .ZN(G393));
  NAND2_X1  g0934(.A1(new_n1049), .A2(new_n758), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1044), .A2(new_n829), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n1136), .B(KEYINPUT115), .ZN(new_n1137));
  NOR3_X1   g0937(.A1(new_n239), .A2(new_n701), .A3(new_n249), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n819), .B1(new_n205), .B2(new_n218), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n759), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n800), .ZN(new_n1141));
  INV_X1    g0941(.A(G283), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n333), .B1(new_n833), .B2(new_n1142), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1144), .B1(new_n792), .B2(new_n785), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1145), .B1(G294), .B2(new_n770), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n1146), .B1(new_n619), .B2(new_n778), .C1(new_n610), .C2(new_n789), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n768), .A2(new_n996), .B1(new_n791), .B2(new_n772), .ZN(new_n1148));
  XOR2_X1   g0948(.A(new_n1148), .B(KEYINPUT52), .Z(new_n1149));
  NAND2_X1  g0949(.A1(new_n837), .A2(new_n384), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n779), .A2(G77), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n839), .A2(G50), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n249), .B1(new_n833), .B2(new_n349), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n832), .B(new_n1153), .C1(G143), .C2(new_n786), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1150), .A2(new_n1151), .A3(new_n1152), .A4(new_n1154), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n768), .A2(new_n289), .B1(new_n791), .B2(new_n796), .ZN(new_n1156));
  XOR2_X1   g0956(.A(KEYINPUT116), .B(KEYINPUT51), .Z(new_n1157));
  XNOR2_X1  g0957(.A(new_n1156), .B(new_n1157), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n1147), .A2(new_n1149), .B1(new_n1155), .B2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1140), .B1(new_n1159), .B2(new_n815), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1137), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1135), .A2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1100), .A2(new_n1092), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n702), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1100), .A2(new_n1092), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1162), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(G390));
  INV_X1    g0968(.A(new_n879), .ZN(new_n1169));
  AND2_X1   g0969(.A1(new_n745), .A2(new_n746), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n662), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n654), .B1(new_n1171), .B2(new_n742), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n694), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1169), .B1(new_n1173), .B2(new_n863), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(new_n967), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n925), .B1(new_n936), .B2(new_n919), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n926), .B1(new_n880), .B2(new_n900), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1178), .A2(new_n938), .A3(new_n941), .ZN(new_n1179));
  OAI211_X1 g0979(.A(G330), .B(new_n862), .C1(new_n725), .C2(new_n732), .ZN(new_n1180));
  OR2_X1    g0980(.A1(new_n1180), .A2(new_n900), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1177), .A2(new_n1179), .A3(new_n1181), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n920), .A2(KEYINPUT39), .B1(new_n936), .B2(new_n937), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n1183), .A2(new_n1178), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1184));
  AND3_X1   g0984(.A1(new_n959), .A2(G330), .A3(new_n862), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT117), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1185), .A2(new_n967), .A3(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n959), .A2(G330), .A3(new_n862), .ZN(new_n1188));
  OAI21_X1  g0988(.A(KEYINPUT117), .B1(new_n900), .B2(new_n1188), .ZN(new_n1189));
  AND2_X1   g0989(.A1(new_n1187), .A2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1182), .B1(new_n1184), .B2(new_n1190), .ZN(new_n1191));
  OR2_X1    g0991(.A1(new_n1191), .A2(new_n757), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n760), .B1(new_n281), .B2(new_n853), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(KEYINPUT54), .B(G143), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n837), .A2(new_n1195), .B1(G159), .B2(new_n779), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n249), .B1(new_n782), .B2(new_n202), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(G125), .B2(new_n786), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n765), .A2(G150), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(new_n1199), .B(KEYINPUT53), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(G132), .B2(new_n835), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(G128), .A2(new_n840), .B1(new_n839), .B2(G137), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1196), .A2(new_n1198), .A3(new_n1201), .A4(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n837), .A2(G97), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n786), .A2(G294), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n249), .B1(new_n765), .B2(G87), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n849), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(G116), .B2(new_n835), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(G107), .A2(new_n839), .B1(new_n840), .B2(G283), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1204), .A2(new_n1151), .A3(new_n1208), .A4(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1203), .A2(new_n1210), .ZN(new_n1211));
  AND2_X1   g1011(.A1(new_n1211), .A2(KEYINPUT119), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n815), .B1(new_n1211), .B2(KEYINPUT119), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1193), .B1(new_n1212), .B2(new_n1213), .C1(new_n945), .C2(new_n817), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1180), .A2(new_n900), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1187), .A2(new_n1189), .A3(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n880), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n879), .B1(new_n748), .B2(new_n862), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1181), .B(new_n1219), .C1(new_n967), .C2(new_n1185), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1218), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n959), .ZN(new_n1222));
  NOR3_X1   g1022(.A1(new_n456), .A2(new_n761), .A3(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n456), .B1(KEYINPUT29), .B2(new_n748), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n648), .B(new_n1223), .C1(new_n740), .C2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1221), .A2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT118), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1221), .A2(new_n1225), .A3(KEYINPUT118), .ZN(new_n1229));
  AND3_X1   g1029(.A1(new_n1228), .A2(new_n1191), .A3(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n702), .B1(new_n1191), .B2(new_n1226), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1192), .B(new_n1214), .C1(new_n1230), .C2(new_n1231), .ZN(G378));
  AOI21_X1  g1032(.A(new_n761), .B1(new_n972), .B2(new_n973), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n904), .A2(new_n298), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(new_n315), .B(new_n1235), .ZN(new_n1236));
  XNOR2_X1  g1036(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1237));
  XNOR2_X1  g1037(.A(new_n1236), .B(new_n1237), .ZN(new_n1238));
  AND3_X1   g1038(.A1(new_n1233), .A2(new_n971), .A3(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1238), .B1(new_n1233), .B2(new_n971), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n943), .A2(new_n948), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1233), .A2(new_n971), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1238), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  OAI21_X1  g1044(.A(KEYINPUT105), .B1(new_n924), .B2(new_n942), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n946), .A2(new_n944), .A3(new_n947), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1233), .A2(new_n971), .A3(new_n1238), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1244), .A2(new_n1245), .A3(new_n1246), .A4(new_n1247), .ZN(new_n1248));
  AND2_X1   g1048(.A1(new_n1241), .A2(new_n1248), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1225), .B1(new_n1191), .B2(new_n1226), .ZN(new_n1250));
  AOI21_X1  g1050(.A(KEYINPUT57), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1250), .A2(KEYINPUT57), .A3(new_n1248), .A4(new_n1241), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(new_n702), .ZN(new_n1253));
  OR2_X1    g1053(.A1(new_n1251), .A2(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1241), .A2(new_n1248), .A3(new_n758), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n759), .B1(G50), .B2(new_n854), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n249), .A2(G41), .ZN(new_n1257));
  AOI211_X1 g1057(.A(G50), .B(new_n1257), .C1(new_n318), .C2(new_n256), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n783), .A2(new_n1005), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n786), .A2(G283), .ZN(new_n1260));
  AND4_X1   g1060(.A1(new_n1117), .A2(new_n1259), .A3(new_n1260), .A4(new_n1257), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n835), .A2(G107), .B1(new_n380), .B2(new_n770), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(G97), .A2(new_n839), .B1(new_n840), .B2(G116), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1012), .A2(new_n1261), .A3(new_n1262), .A4(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT58), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1258), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  OAI22_X1  g1066(.A1(new_n771), .A2(new_n1008), .B1(new_n833), .B2(new_n1194), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1267), .B1(G128), .B2(new_n835), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(G125), .A2(new_n840), .B1(new_n839), .B2(G132), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1268), .B(new_n1269), .C1(new_n289), .C2(new_n778), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(KEYINPUT59), .ZN(new_n1271));
  OAI211_X1 g1071(.A(new_n318), .B(new_n256), .C1(new_n782), .C2(new_n796), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1272), .B1(G124), .B2(new_n786), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1271), .A2(new_n1273), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1270), .A2(KEYINPUT59), .ZN(new_n1275));
  OAI221_X1 g1075(.A(new_n1266), .B1(new_n1265), .B2(new_n1264), .C1(new_n1274), .C2(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1256), .B1(new_n1276), .B2(new_n815), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1277), .B1(new_n1238), .B2(new_n817), .ZN(new_n1278));
  AND2_X1   g1078(.A1(new_n1255), .A2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1254), .A2(new_n1279), .ZN(G375));
  INV_X1    g1080(.A(new_n1223), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n649), .B(new_n1281), .C1(new_n953), .C2(new_n955), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1282), .A2(new_n1218), .A3(new_n1220), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1228), .A2(new_n1094), .A3(new_n1229), .A4(new_n1283), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1259), .B(new_n249), .C1(new_n796), .C2(new_n833), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1285), .B1(G128), .B2(new_n786), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n779), .A2(G50), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(new_n835), .A2(G137), .B1(G150), .B2(new_n770), .ZN(new_n1288));
  AOI22_X1  g1088(.A1(G132), .A2(new_n840), .B1(new_n839), .B2(new_n1195), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1286), .A2(new_n1287), .A3(new_n1288), .A4(new_n1289), .ZN(new_n1290));
  OAI22_X1  g1090(.A1(new_n778), .A2(new_n378), .B1(new_n1142), .B2(new_n791), .ZN(new_n1291));
  XNOR2_X1  g1091(.A(new_n1291), .B(KEYINPUT120), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n786), .A2(G303), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n249), .B1(new_n765), .B2(G97), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1293), .A2(new_n1007), .A3(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1295), .B1(G294), .B2(new_n840), .ZN(new_n1296));
  OAI221_X1 g1096(.A(new_n1296), .B1(new_n206), .B2(new_n809), .C1(new_n619), .C2(new_n789), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1290), .B1(new_n1292), .B2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT121), .ZN(new_n1299));
  AND2_X1   g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n815), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1301));
  OAI221_X1 g1101(.A(new_n759), .B1(G68), .B2(new_n854), .C1(new_n1300), .C2(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1302), .B1(new_n816), .B2(new_n900), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1303), .B1(new_n1221), .B2(new_n758), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1284), .A2(new_n1304), .ZN(G381));
  NAND2_X1  g1105(.A1(new_n1192), .A2(new_n1214), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1231), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1228), .A2(new_n1191), .A3(new_n1229), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1306), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1254), .A2(new_n1309), .A3(new_n1279), .ZN(new_n1310));
  OAI211_X1 g1110(.A(new_n1025), .B(new_n1167), .C1(new_n1085), .C2(new_n1097), .ZN(new_n1311));
  INV_X1    g1111(.A(G396), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1312), .A2(new_n1101), .A3(new_n1133), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(new_n876), .ZN(new_n1315));
  OR4_X1    g1115(.A1(G381), .A2(new_n1310), .A3(new_n1311), .A4(new_n1315), .ZN(G407));
  OAI211_X1 g1116(.A(G407), .B(G213), .C1(G343), .C2(new_n1310), .ZN(G409));
  INV_X1    g1117(.A(KEYINPUT122), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1255), .A2(new_n1318), .A3(new_n1278), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1250), .A2(new_n1094), .A3(new_n1248), .A4(new_n1241), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1318), .B1(new_n1255), .B2(new_n1278), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1309), .B1(new_n1321), .B2(new_n1322), .ZN(new_n1323));
  OAI211_X1 g1123(.A(G378), .B(new_n1279), .C1(new_n1251), .C2(new_n1253), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(G213), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1326), .A2(G343), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT60), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1283), .A2(new_n1329), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1282), .A2(new_n1218), .A3(KEYINPUT60), .A4(new_n1220), .ZN(new_n1331));
  NAND4_X1  g1131(.A1(new_n1330), .A2(new_n702), .A3(new_n1226), .A4(new_n1331), .ZN(new_n1332));
  AND3_X1   g1132(.A1(new_n1332), .A2(G384), .A3(new_n1304), .ZN(new_n1333));
  AOI21_X1  g1133(.A(G384), .B1(new_n1332), .B2(new_n1304), .ZN(new_n1334));
  NOR2_X1   g1134(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1325), .A2(new_n1328), .A3(new_n1335), .ZN(new_n1336));
  NOR2_X1   g1136(.A1(new_n1336), .A2(KEYINPUT62), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT61), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1327), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1327), .A2(G2897), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1340), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1332), .A2(new_n1304), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1342), .A2(new_n876), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1332), .A2(G384), .A3(new_n1304), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1340), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1343), .A2(new_n1344), .A3(new_n1345), .ZN(new_n1346));
  AND2_X1   g1146(.A1(new_n1341), .A2(new_n1346), .ZN(new_n1347));
  OAI21_X1  g1147(.A(new_n1338), .B1(new_n1339), .B2(new_n1347), .ZN(new_n1348));
  INV_X1    g1148(.A(KEYINPUT62), .ZN(new_n1349));
  AOI21_X1  g1149(.A(new_n1349), .B1(new_n1339), .B2(new_n1335), .ZN(new_n1350));
  NOR3_X1   g1150(.A1(new_n1337), .A2(new_n1348), .A3(new_n1350), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(G387), .A2(G390), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(G393), .A2(G396), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1353), .A2(new_n1313), .ZN(new_n1354));
  INV_X1    g1154(.A(KEYINPUT125), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1354), .A2(new_n1355), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1353), .A2(KEYINPUT125), .A3(new_n1313), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1356), .A2(new_n1357), .ZN(new_n1358));
  NAND3_X1  g1158(.A1(new_n1352), .A2(new_n1358), .A3(new_n1311), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1359), .A2(KEYINPUT126), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1352), .A2(new_n1311), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1361), .A2(new_n1354), .ZN(new_n1362));
  INV_X1    g1162(.A(KEYINPUT126), .ZN(new_n1363));
  NAND4_X1  g1163(.A1(new_n1352), .A2(new_n1358), .A3(new_n1363), .A4(new_n1311), .ZN(new_n1364));
  NAND3_X1  g1164(.A1(new_n1360), .A2(new_n1362), .A3(new_n1364), .ZN(new_n1365));
  XOR2_X1   g1165(.A(KEYINPUT123), .B(KEYINPUT63), .Z(new_n1366));
  NAND2_X1  g1166(.A1(new_n1336), .A2(new_n1366), .ZN(new_n1367));
  INV_X1    g1167(.A(KEYINPUT124), .ZN(new_n1368));
  AND3_X1   g1168(.A1(new_n1341), .A2(new_n1346), .A3(new_n1368), .ZN(new_n1369));
  AOI21_X1  g1169(.A(new_n1368), .B1(new_n1341), .B2(new_n1346), .ZN(new_n1370));
  NOR2_X1   g1170(.A1(new_n1369), .A2(new_n1370), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1325), .A2(new_n1328), .ZN(new_n1372));
  NAND2_X1  g1172(.A1(new_n1371), .A2(new_n1372), .ZN(new_n1373));
  NAND4_X1  g1173(.A1(new_n1367), .A2(new_n1373), .A3(new_n1365), .A4(new_n1338), .ZN(new_n1374));
  NAND4_X1  g1174(.A1(new_n1325), .A2(KEYINPUT63), .A3(new_n1328), .A4(new_n1335), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(new_n1375), .A2(KEYINPUT127), .ZN(new_n1376));
  INV_X1    g1176(.A(KEYINPUT127), .ZN(new_n1377));
  NAND4_X1  g1177(.A1(new_n1339), .A2(new_n1377), .A3(KEYINPUT63), .A4(new_n1335), .ZN(new_n1378));
  NAND2_X1  g1178(.A1(new_n1376), .A2(new_n1378), .ZN(new_n1379));
  OAI22_X1  g1179(.A1(new_n1351), .A2(new_n1365), .B1(new_n1374), .B2(new_n1379), .ZN(G405));
  AOI21_X1  g1180(.A(G378), .B1(new_n1254), .B2(new_n1279), .ZN(new_n1381));
  INV_X1    g1181(.A(new_n1324), .ZN(new_n1382));
  OAI21_X1  g1182(.A(new_n1335), .B1(new_n1381), .B2(new_n1382), .ZN(new_n1383));
  INV_X1    g1183(.A(new_n1383), .ZN(new_n1384));
  NOR3_X1   g1184(.A1(new_n1381), .A2(new_n1382), .A3(new_n1335), .ZN(new_n1385));
  NOR3_X1   g1185(.A1(new_n1384), .A2(new_n1365), .A3(new_n1385), .ZN(new_n1386));
  OR3_X1    g1186(.A1(new_n1381), .A2(new_n1382), .A3(new_n1335), .ZN(new_n1387));
  AND2_X1   g1187(.A1(new_n1362), .A2(new_n1364), .ZN(new_n1388));
  AOI22_X1  g1188(.A1(new_n1387), .A2(new_n1383), .B1(new_n1388), .B2(new_n1360), .ZN(new_n1389));
  NOR2_X1   g1189(.A1(new_n1386), .A2(new_n1389), .ZN(G402));
endmodule


