//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 1 0 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 0 0 0 0 1 1 1 1 1 0 1 1 0 0 0 0 0 1 1 1 1 0 0 1 1 1 1 1 1 1 1 0 1 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:18 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n793, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n994, new_n995, new_n996,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076;
  INV_X1    g000(.A(G140), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G125), .ZN(new_n188));
  INV_X1    g002(.A(G125), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G140), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n188), .A2(new_n190), .A3(KEYINPUT16), .ZN(new_n191));
  OR3_X1    g005(.A1(new_n189), .A2(KEYINPUT16), .A3(G140), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(new_n192), .A3(G146), .ZN(new_n193));
  XOR2_X1   g007(.A(new_n193), .B(KEYINPUT74), .Z(new_n194));
  INV_X1    g008(.A(G146), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n188), .A2(new_n190), .A3(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G128), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G119), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT23), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  OR2_X1    g014(.A1(new_n197), .A2(G119), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n197), .A2(KEYINPUT23), .A3(G119), .ZN(new_n202));
  AND3_X1   g016(.A1(new_n200), .A2(new_n201), .A3(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G110), .ZN(new_n204));
  AND2_X1   g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n201), .A2(new_n198), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT24), .B(G110), .ZN(new_n207));
  AND2_X1   g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  OAI211_X1 g022(.A(new_n194), .B(new_n196), .C1(new_n205), .C2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n193), .A2(KEYINPUT73), .ZN(new_n210));
  AOI21_X1  g024(.A(G146), .B1(new_n191), .B2(new_n192), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AOI211_X1 g026(.A(KEYINPUT73), .B(G146), .C1(new_n191), .C2(new_n192), .ZN(new_n213));
  OAI22_X1  g027(.A1(new_n203), .A2(new_n204), .B1(new_n206), .B2(new_n207), .ZN(new_n214));
  OR3_X1    g028(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n209), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(KEYINPUT22), .B(G137), .ZN(new_n217));
  INV_X1    g031(.A(G221), .ZN(new_n218));
  INV_X1    g032(.A(G234), .ZN(new_n219));
  NOR3_X1   g033(.A1(new_n218), .A2(new_n219), .A3(G953), .ZN(new_n220));
  XOR2_X1   g034(.A(new_n217), .B(new_n220), .Z(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n216), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G902), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n209), .A2(new_n215), .A3(new_n221), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT25), .ZN(new_n227));
  OAI21_X1  g041(.A(G217), .B1(new_n219), .B2(G902), .ZN(new_n228));
  XNOR2_X1  g042(.A(new_n228), .B(KEYINPUT72), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT25), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n223), .A2(new_n231), .A3(new_n224), .A4(new_n225), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n227), .A2(new_n230), .A3(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n230), .A2(G902), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n223), .A2(new_n225), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(G472), .A2(G902), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT66), .ZN(new_n240));
  XNOR2_X1  g054(.A(G134), .B(G137), .ZN(new_n241));
  INV_X1    g055(.A(G131), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n240), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT11), .ZN(new_n244));
  INV_X1    g058(.A(G134), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n244), .B1(new_n245), .B2(G137), .ZN(new_n246));
  INV_X1    g060(.A(G137), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n247), .A2(KEYINPUT11), .A3(G134), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n245), .A2(G137), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n246), .A2(new_n248), .A3(new_n242), .A4(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n245), .A2(G137), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n247), .A2(G134), .ZN(new_n252));
  OAI211_X1 g066(.A(KEYINPUT66), .B(G131), .C1(new_n251), .C2(new_n252), .ZN(new_n253));
  AND3_X1   g067(.A1(new_n243), .A2(new_n250), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n195), .A2(G143), .ZN(new_n255));
  INV_X1    g069(.A(G143), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G146), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n255), .A2(KEYINPUT1), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n258), .A2(new_n259), .A3(G128), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n255), .B(new_n257), .C1(KEYINPUT1), .C2(new_n197), .ZN(new_n261));
  AND3_X1   g075(.A1(new_n260), .A2(KEYINPUT67), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(KEYINPUT67), .B1(new_n260), .B2(new_n261), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n254), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(KEYINPUT0), .A2(G128), .ZN(new_n265));
  OAI21_X1  g079(.A(KEYINPUT65), .B1(new_n258), .B2(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(G143), .B(G146), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT65), .ZN(new_n268));
  AND2_X1   g082(.A1(KEYINPUT0), .A2(G128), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  NOR2_X1   g084(.A1(KEYINPUT0), .A2(G128), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  AOI22_X1  g086(.A1(new_n266), .A2(new_n270), .B1(new_n258), .B2(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n246), .A2(new_n249), .A3(new_n248), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(G131), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(new_n250), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  XNOR2_X1  g091(.A(G116), .B(G119), .ZN(new_n278));
  XNOR2_X1  g092(.A(KEYINPUT2), .B(G113), .ZN(new_n279));
  XNOR2_X1  g093(.A(new_n278), .B(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n264), .A2(new_n277), .A3(new_n280), .ZN(new_n281));
  AND2_X1   g095(.A1(new_n275), .A2(new_n250), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n258), .A2(new_n272), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n268), .B1(new_n267), .B2(new_n269), .ZN(new_n284));
  AND4_X1   g098(.A1(new_n268), .A2(new_n255), .A3(new_n257), .A4(new_n269), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n283), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n243), .A2(new_n250), .A3(new_n253), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n260), .A2(new_n261), .ZN(new_n288));
  OAI22_X1  g102(.A1(new_n282), .A2(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n280), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n281), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT28), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(KEYINPUT68), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT68), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n292), .A2(new_n295), .A3(KEYINPUT28), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT67), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n288), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n260), .A2(KEYINPUT67), .A3(new_n261), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n287), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n282), .A2(new_n286), .ZN(new_n301));
  OAI21_X1  g115(.A(KEYINPUT69), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT69), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n264), .A2(new_n277), .A3(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n302), .A2(new_n280), .A3(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT28), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n294), .A2(new_n296), .A3(new_n307), .ZN(new_n308));
  NOR2_X1   g122(.A1(G237), .A2(G953), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G210), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n310), .B(KEYINPUT27), .ZN(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT26), .B(G101), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n311), .B(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n308), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n264), .A2(new_n277), .A3(KEYINPUT30), .ZN(new_n316));
  XOR2_X1   g130(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n317));
  NAND2_X1  g131(.A1(new_n289), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n316), .A2(new_n318), .A3(new_n290), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n319), .A2(new_n313), .A3(new_n281), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(KEYINPUT31), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT31), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n319), .A2(new_n322), .A3(new_n313), .A4(new_n281), .ZN(new_n323));
  AND2_X1   g137(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n239), .B1(new_n315), .B2(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(KEYINPUT70), .B1(new_n325), .B2(KEYINPUT32), .ZN(new_n326));
  AOI22_X1  g140(.A1(new_n293), .A2(KEYINPUT68), .B1(new_n305), .B2(new_n306), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n313), .B1(new_n327), .B2(new_n296), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n321), .A2(new_n323), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n238), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT70), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT32), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n326), .A2(new_n333), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n239), .A2(new_n332), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n335), .B1(new_n328), .B2(new_n329), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT71), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n294), .A2(new_n313), .A3(new_n296), .A4(new_n307), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n313), .B1(new_n319), .B2(new_n281), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n340), .A2(KEYINPUT29), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n290), .B1(new_n300), .B2(new_n301), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n306), .B1(new_n343), .B2(new_n281), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n344), .B1(new_n306), .B2(new_n305), .ZN(new_n345));
  AND2_X1   g159(.A1(new_n313), .A2(KEYINPUT29), .ZN(new_n346));
  AOI21_X1  g160(.A(G902), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n342), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(G472), .ZN(new_n349));
  OAI211_X1 g163(.A(KEYINPUT71), .B(new_n335), .C1(new_n328), .C2(new_n329), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n338), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n237), .B1(new_n334), .B2(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(G214), .B1(G237), .B2(G902), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n353), .B(KEYINPUT81), .ZN(new_n354));
  INV_X1    g168(.A(G107), .ZN(new_n355));
  OAI21_X1  g169(.A(KEYINPUT76), .B1(new_n355), .B2(G104), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT76), .ZN(new_n357));
  INV_X1    g171(.A(G104), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(new_n358), .A3(G107), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n355), .A2(G104), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n356), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  AND2_X1   g175(.A1(new_n361), .A2(G101), .ZN(new_n362));
  INV_X1    g176(.A(G101), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n363), .B1(new_n355), .B2(G104), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n355), .A2(KEYINPUT75), .A3(G104), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT3), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n355), .A2(KEYINPUT75), .A3(KEYINPUT3), .A4(G104), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n364), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(KEYINPUT77), .B1(new_n362), .B2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n278), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n371), .A2(new_n279), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n278), .A2(KEYINPUT5), .ZN(new_n373));
  INV_X1    g187(.A(G116), .ZN(new_n374));
  NOR3_X1   g188(.A1(new_n374), .A2(KEYINPUT5), .A3(G119), .ZN(new_n375));
  INV_X1    g189(.A(G113), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n372), .B1(new_n373), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n364), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n358), .A2(G107), .ZN(new_n380));
  AOI21_X1  g194(.A(KEYINPUT3), .B1(new_n380), .B2(KEYINPUT75), .ZN(new_n381));
  INV_X1    g195(.A(new_n368), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n379), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT77), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n361), .A2(G101), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n370), .A2(new_n378), .A3(new_n386), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n355), .A2(G104), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n388), .B1(new_n367), .B2(new_n368), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n383), .B(KEYINPUT4), .C1(new_n363), .C2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT4), .ZN(new_n391));
  AND2_X1   g205(.A1(new_n367), .A2(new_n368), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n391), .B(G101), .C1(new_n392), .C2(new_n388), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n390), .A2(new_n290), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n387), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(KEYINPUT82), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT6), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT82), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n387), .A2(new_n394), .A3(new_n398), .ZN(new_n399));
  XNOR2_X1  g213(.A(G110), .B(G122), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n396), .A2(new_n397), .A3(new_n399), .A4(new_n401), .ZN(new_n402));
  AND3_X1   g216(.A1(new_n387), .A2(new_n394), .A3(new_n398), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n398), .B1(new_n387), .B2(new_n394), .ZN(new_n404));
  NOR3_X1   g218(.A1(new_n403), .A2(new_n404), .A3(new_n400), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n387), .A2(new_n394), .A3(new_n400), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(KEYINPUT6), .ZN(new_n407));
  OAI211_X1 g221(.A(KEYINPUT83), .B(new_n402), .C1(new_n405), .C2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n396), .A2(new_n399), .A3(new_n401), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT83), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n409), .A2(new_n410), .A3(KEYINPUT6), .A4(new_n406), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n288), .A2(new_n189), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n413), .B1(new_n273), .B2(new_n189), .ZN(new_n414));
  INV_X1    g228(.A(G224), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n415), .A2(G953), .ZN(new_n416));
  XOR2_X1   g230(.A(new_n414), .B(new_n416), .Z(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n412), .A2(new_n418), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n395), .A2(new_n401), .ZN(new_n420));
  OAI21_X1  g234(.A(KEYINPUT7), .B1(new_n415), .B2(G953), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n414), .A2(KEYINPUT84), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n414), .A2(new_n421), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT84), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n420), .B1(new_n422), .B2(new_n425), .ZN(new_n426));
  OR3_X1    g240(.A1(new_n414), .A2(KEYINPUT85), .A3(new_n421), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n383), .A2(new_n385), .ZN(new_n428));
  OR2_X1    g242(.A1(new_n378), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n378), .A2(new_n428), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n400), .B(KEYINPUT8), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n429), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(KEYINPUT85), .B1(new_n414), .B2(new_n421), .ZN(new_n433));
  AND3_X1   g247(.A1(new_n427), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(G902), .B1(new_n426), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(G210), .B1(G237), .B2(G902), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n419), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n436), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n417), .B1(new_n408), .B2(new_n411), .ZN(new_n439));
  INV_X1    g253(.A(new_n435), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n354), .B1(new_n437), .B2(new_n441), .ZN(new_n442));
  XNOR2_X1  g256(.A(G113), .B(G122), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n443), .B(new_n358), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT89), .ZN(new_n445));
  INV_X1    g259(.A(G237), .ZN(new_n446));
  INV_X1    g260(.A(G953), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(new_n447), .A3(G214), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n256), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n309), .A2(G143), .A3(G214), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(KEYINPUT18), .A2(G131), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(KEYINPUT86), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT86), .ZN(new_n455));
  AOI211_X1 g269(.A(new_n455), .B(new_n452), .C1(new_n449), .C2(new_n450), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n195), .B1(new_n188), .B2(new_n190), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n457), .B1(KEYINPUT87), .B2(new_n196), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n188), .A2(new_n190), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n459), .A2(KEYINPUT87), .A3(G146), .ZN(new_n460));
  OAI22_X1  g274(.A1(new_n454), .A2(new_n456), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n449), .A2(new_n450), .A3(new_n452), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT88), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n449), .A2(KEYINPUT88), .A3(new_n450), .A4(new_n452), .ZN(new_n465));
  AND2_X1   g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n445), .B1(new_n461), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n448), .A2(new_n256), .ZN(new_n468));
  AOI21_X1  g282(.A(G143), .B1(new_n309), .B2(G214), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n455), .B1(new_n470), .B2(new_n452), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n451), .A2(KEYINPUT86), .A3(new_n453), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n464), .A2(new_n465), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n196), .A2(KEYINPUT87), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n459), .A2(G146), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n475), .B(new_n476), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n473), .A2(KEYINPUT89), .A3(new_n474), .A4(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n467), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n470), .A2(new_n242), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n451), .A2(G131), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT19), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n459), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(KEYINPUT19), .B1(new_n188), .B2(new_n190), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n195), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT90), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AND2_X1   g302(.A1(new_n486), .A2(new_n487), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n194), .B(new_n482), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n444), .B1(new_n479), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT17), .ZN(new_n492));
  AND3_X1   g306(.A1(new_n480), .A2(new_n492), .A3(new_n481), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n451), .A2(KEYINPUT17), .A3(G131), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n191), .A2(new_n192), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n195), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n497), .A2(KEYINPUT73), .A3(new_n193), .ZN(new_n498));
  INV_X1    g312(.A(new_n213), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n495), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n493), .B1(new_n500), .B2(KEYINPUT91), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n494), .B1(new_n212), .B2(new_n213), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT91), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AOI22_X1  g318(.A1(new_n501), .A2(new_n504), .B1(new_n467), .B2(new_n478), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n491), .B1(new_n444), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(G475), .A2(G902), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(KEYINPUT20), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n491), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n501), .A2(new_n504), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n511), .A2(new_n444), .A3(new_n479), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT20), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n513), .A2(new_n514), .A3(new_n507), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n509), .A2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT94), .ZN(new_n517));
  OAI21_X1  g331(.A(KEYINPUT92), .B1(new_n197), .B2(G143), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT92), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n519), .A2(new_n256), .A3(G128), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  AND2_X1   g335(.A1(KEYINPUT93), .A2(KEYINPUT13), .ZN(new_n522));
  NOR2_X1   g336(.A1(KEYINPUT93), .A2(KEYINPUT13), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n517), .B1(new_n521), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n256), .A2(G128), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n526), .B1(new_n521), .B2(new_n524), .ZN(new_n527));
  XNOR2_X1  g341(.A(KEYINPUT93), .B(KEYINPUT13), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n528), .A2(KEYINPUT94), .A3(new_n518), .A4(new_n520), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n525), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(G134), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT95), .ZN(new_n532));
  AOI211_X1 g346(.A(new_n532), .B(new_n526), .C1(new_n518), .C2(new_n520), .ZN(new_n533));
  INV_X1    g347(.A(new_n526), .ZN(new_n534));
  AOI21_X1  g348(.A(KEYINPUT95), .B1(new_n521), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n245), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  XNOR2_X1  g350(.A(G116), .B(G122), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n537), .B(G107), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n531), .A2(new_n536), .A3(new_n539), .ZN(new_n540));
  OR2_X1    g354(.A1(new_n374), .A2(G122), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n355), .B1(new_n541), .B2(KEYINPUT14), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n542), .B(new_n537), .ZN(new_n543));
  NOR3_X1   g357(.A1(new_n533), .A2(new_n535), .A3(new_n245), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n519), .B1(G128), .B2(new_n256), .ZN(new_n545));
  NOR3_X1   g359(.A1(new_n197), .A2(KEYINPUT92), .A3(G143), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n534), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n532), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n521), .A2(KEYINPUT95), .A3(new_n534), .ZN(new_n549));
  AOI21_X1  g363(.A(G134), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n543), .B1(new_n544), .B2(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(KEYINPUT9), .B(G234), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n553), .A2(G217), .A3(new_n447), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n540), .A2(new_n551), .A3(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n555), .B1(new_n540), .B2(new_n551), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n224), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(G478), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n561), .A2(KEYINPUT15), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n559), .A2(new_n562), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  AND3_X1   g381(.A1(new_n511), .A2(new_n444), .A3(new_n479), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n444), .B1(new_n511), .B2(new_n479), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n224), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(G475), .ZN(new_n571));
  AND2_X1   g385(.A1(new_n447), .A2(G952), .ZN(new_n572));
  NAND2_X1  g386(.A1(G234), .A2(G237), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n573), .A2(G902), .A3(G953), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(KEYINPUT21), .B(G898), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n575), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n516), .A2(new_n567), .A3(new_n571), .A4(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n218), .B1(new_n553), .B2(new_n224), .ZN(new_n583));
  INV_X1    g397(.A(G469), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n584), .A2(new_n224), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n428), .A2(new_n288), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n383), .A2(new_n261), .A3(new_n260), .A4(new_n385), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n586), .A2(KEYINPUT79), .A3(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT79), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n428), .A2(new_n589), .A3(new_n288), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(KEYINPUT80), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT80), .ZN(new_n593));
  OR2_X1    g407(.A1(new_n593), .A2(KEYINPUT78), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n588), .B(new_n590), .C1(KEYINPUT12), .C2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n592), .A2(new_n276), .A3(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT10), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n587), .A2(new_n597), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n370), .A2(new_n386), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n597), .B1(new_n298), .B2(new_n299), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n390), .A2(new_n273), .A3(new_n393), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n601), .A2(new_n282), .A3(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(G110), .B(G140), .ZN(new_n604));
  INV_X1    g418(.A(G227), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n605), .A2(G953), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n604), .B(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  OR2_X1    g422(.A1(new_n282), .A2(KEYINPUT78), .ZN(new_n609));
  OAI21_X1  g423(.A(KEYINPUT12), .B1(new_n591), .B2(new_n609), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n596), .A2(new_n603), .A3(new_n608), .A4(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n282), .B1(new_n601), .B2(new_n602), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n298), .A2(new_n299), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n613), .A2(KEYINPUT10), .A3(new_n370), .A4(new_n386), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n587), .A2(new_n597), .ZN(new_n615));
  AND4_X1   g429(.A1(new_n282), .A2(new_n614), .A3(new_n602), .A4(new_n615), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n607), .B1(new_n612), .B2(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(G902), .B1(new_n611), .B2(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n585), .B1(new_n618), .B2(new_n584), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n596), .A2(new_n603), .A3(new_n610), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n607), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n614), .A2(new_n602), .A3(new_n615), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n276), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n603), .A2(new_n623), .A3(new_n608), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n621), .A2(G469), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n583), .B1(new_n619), .B2(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n442), .A2(new_n582), .A3(new_n626), .ZN(new_n627));
  OR2_X1    g441(.A1(new_n352), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(G101), .ZN(G3));
  NAND2_X1  g443(.A1(new_n437), .A2(new_n441), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n630), .A2(new_n353), .A3(new_n580), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT99), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n560), .A2(G478), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT33), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n634), .B1(new_n557), .B2(new_n558), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n550), .A2(new_n538), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n548), .A2(new_n549), .A3(G134), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n536), .A2(new_n638), .ZN(new_n639));
  AOI22_X1  g453(.A1(new_n637), .A2(new_n531), .B1(new_n639), .B2(new_n543), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n554), .B1(new_n640), .B2(KEYINPUT96), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n540), .A2(new_n551), .A3(KEYINPUT96), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  OAI21_X1  g457(.A(KEYINPUT33), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n640), .A2(KEYINPUT97), .A3(new_n555), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT97), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n556), .A2(new_n646), .ZN(new_n647));
  AND2_X1   g461(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  OAI21_X1  g462(.A(KEYINPUT98), .B1(new_n644), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n540), .A2(new_n551), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT96), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n555), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n634), .B1(new_n652), .B2(new_n642), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT98), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n645), .A2(new_n647), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n636), .B1(new_n649), .B2(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n561), .A2(G902), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n633), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  AOI22_X1  g473(.A1(new_n509), .A2(new_n515), .B1(G475), .B2(new_n570), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n632), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n650), .A2(new_n651), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n662), .A2(new_n554), .A3(new_n642), .ZN(new_n663));
  AND4_X1   g477(.A1(new_n654), .A2(new_n655), .A3(KEYINPUT33), .A4(new_n663), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n654), .B1(new_n653), .B2(new_n655), .ZN(new_n665));
  OAI211_X1 g479(.A(new_n635), .B(new_n658), .C1(new_n664), .C2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n633), .ZN(new_n667));
  AOI22_X1  g481(.A1(new_n666), .A2(new_n667), .B1(new_n516), .B2(new_n571), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(KEYINPUT99), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n631), .B1(new_n661), .B2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n626), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n224), .B1(new_n328), .B2(new_n329), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n325), .B1(G472), .B2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n671), .A2(new_n674), .A3(new_n236), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n670), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT34), .B(G104), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G6));
  INV_X1    g492(.A(new_n353), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n679), .B1(new_n437), .B2(new_n441), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n579), .B(KEYINPUT101), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT100), .ZN(new_n682));
  OAI22_X1  g496(.A1(new_n502), .A2(new_n503), .B1(KEYINPUT17), .B2(new_n482), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n500), .A2(KEYINPUT91), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n479), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n444), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g501(.A(G902), .B1(new_n687), .B2(new_n512), .ZN(new_n688));
  INV_X1    g502(.A(G475), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n682), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n570), .A2(KEYINPUT100), .A3(G475), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AND2_X1   g506(.A1(new_n692), .A2(new_n516), .ZN(new_n693));
  AND4_X1   g507(.A1(new_n566), .A2(new_n680), .A3(new_n681), .A4(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n675), .ZN(new_n695));
  XOR2_X1   g509(.A(KEYINPUT35), .B(G107), .Z(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G9));
  INV_X1    g511(.A(KEYINPUT102), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n222), .A2(KEYINPUT36), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n216), .B(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n234), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n233), .A2(new_n698), .A3(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n698), .B1(new_n233), .B2(new_n701), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n673), .ZN(new_n706));
  OR2_X1    g520(.A1(new_n627), .A2(new_n706), .ZN(new_n707));
  XOR2_X1   g521(.A(KEYINPUT37), .B(G110), .Z(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G12));
  INV_X1    g523(.A(new_n704), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n702), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n325), .A2(KEYINPUT70), .A3(KEYINPUT32), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n331), .B1(new_n330), .B2(new_n332), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  AND3_X1   g528(.A1(new_n338), .A2(new_n349), .A3(new_n350), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n711), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT104), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n436), .B1(new_n419), .B2(new_n435), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n439), .A2(new_n440), .A3(new_n438), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n353), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n447), .A2(G900), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n573), .A2(G902), .ZN(new_n723));
  OR3_X1    g537(.A1(new_n722), .A2(KEYINPUT103), .A3(new_n723), .ZN(new_n724));
  OAI21_X1  g538(.A(KEYINPUT103), .B1(new_n722), .B2(new_n723), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n724), .A2(new_n574), .A3(new_n725), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n692), .A2(new_n516), .A3(new_n566), .A4(new_n726), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n717), .B1(new_n720), .B2(new_n727), .ZN(new_n728));
  AND4_X1   g542(.A1(new_n516), .A2(new_n692), .A3(new_n566), .A4(new_n726), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n729), .A2(KEYINPUT104), .A3(new_n680), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n716), .A2(new_n728), .A3(new_n730), .A4(new_n626), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(KEYINPUT105), .ZN(new_n732));
  OAI211_X1 g546(.A(new_n626), .B(new_n705), .C1(new_n334), .C2(new_n351), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT105), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n734), .A2(new_n735), .A3(new_n728), .A4(new_n730), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n732), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(KEYINPUT106), .B(G128), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n737), .B(new_n738), .ZN(G30));
  NAND2_X1  g553(.A1(new_n315), .A2(new_n324), .ZN(new_n740));
  AOI21_X1  g554(.A(KEYINPUT71), .B1(new_n740), .B2(new_n335), .ZN(new_n741));
  INV_X1    g555(.A(new_n350), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(G472), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n319), .A2(new_n281), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(new_n313), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n343), .A2(new_n314), .A3(new_n281), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n748), .A2(KEYINPUT107), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n748), .A2(KEYINPUT107), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n749), .A2(new_n750), .A3(G902), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n743), .B1(new_n744), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n752), .A2(new_n334), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n233), .A2(new_n701), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n660), .A2(new_n567), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  NOR4_X1   g570(.A1(new_n753), .A2(new_n679), .A3(new_n754), .A4(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n726), .B(KEYINPUT39), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n671), .A2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  OR2_X1    g575(.A1(new_n761), .A2(KEYINPUT40), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(KEYINPUT40), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n630), .B(KEYINPUT38), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n757), .A2(new_n762), .A3(new_n763), .A4(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G143), .ZN(G45));
  INV_X1    g580(.A(KEYINPUT109), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n743), .A2(new_n326), .A3(new_n333), .A4(new_n349), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n768), .A2(new_n626), .A3(new_n680), .A4(new_n705), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n516), .A2(new_n571), .ZN(new_n770));
  INV_X1    g584(.A(new_n666), .ZN(new_n771));
  OAI211_X1 g585(.A(new_n770), .B(new_n726), .C1(new_n771), .C2(new_n633), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(KEYINPUT108), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT108), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n668), .A2(new_n774), .A3(new_n726), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n767), .B1(new_n769), .B2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(new_n726), .ZN(new_n778));
  NOR4_X1   g592(.A1(new_n659), .A2(KEYINPUT108), .A3(new_n660), .A4(new_n778), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n774), .B1(new_n668), .B2(new_n726), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n734), .A2(new_n781), .A3(KEYINPUT109), .A4(new_n680), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n777), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G146), .ZN(G48));
  NOR2_X1   g598(.A1(new_n618), .A2(new_n584), .ZN(new_n785));
  AOI211_X1 g599(.A(G469), .B(G902), .C1(new_n611), .C2(new_n617), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n785), .A2(new_n786), .A3(new_n583), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n237), .B(new_n787), .C1(new_n334), .C2(new_n351), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n670), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(KEYINPUT41), .B(G113), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n790), .B(new_n791), .ZN(G15));
  NAND2_X1  g606(.A1(new_n789), .A2(new_n694), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G116), .ZN(G18));
  INV_X1    g608(.A(new_n787), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n720), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n716), .A2(new_n582), .A3(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G119), .ZN(G21));
  NAND2_X1  g612(.A1(new_n680), .A2(new_n755), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n321), .B(new_n323), .C1(new_n345), .C2(new_n313), .ZN(new_n800));
  AOI22_X1  g614(.A1(new_n672), .A2(G472), .B1(new_n238), .B2(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n787), .A2(new_n801), .A3(new_n237), .A4(new_n681), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n799), .A2(new_n802), .ZN(new_n803));
  XOR2_X1   g617(.A(new_n803), .B(G122), .Z(G24));
  NAND2_X1  g618(.A1(new_n672), .A2(G472), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n800), .A2(new_n238), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n805), .A2(new_n754), .A3(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  AND4_X1   g622(.A1(new_n773), .A2(new_n796), .A3(new_n775), .A4(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(new_n189), .ZN(G27));
  NAND3_X1  g624(.A1(new_n437), .A2(new_n441), .A3(new_n353), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n618), .A2(new_n584), .ZN(new_n812));
  INV_X1    g626(.A(new_n585), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n624), .A2(KEYINPUT110), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT110), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n603), .A2(new_n623), .A3(new_n815), .A4(new_n608), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n621), .A2(G469), .A3(new_n814), .A4(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n812), .A2(new_n813), .A3(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n583), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n352), .A2(new_n811), .A3(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT42), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n821), .A2(new_n822), .A3(new_n781), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n349), .A2(new_n336), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n330), .A2(new_n332), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n236), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n811), .A2(new_n820), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OAI21_X1  g642(.A(KEYINPUT42), .B1(new_n776), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n823), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(new_n242), .ZN(G33));
  NAND2_X1  g645(.A1(new_n821), .A2(new_n729), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(G134), .ZN(G36));
  OAI21_X1  g647(.A(KEYINPUT111), .B1(new_n659), .B2(new_n770), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT43), .ZN(new_n835));
  OR2_X1    g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n834), .A2(new_n835), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n673), .B1(new_n233), .B2(new_n701), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  OR2_X1    g654(.A1(new_n840), .A2(KEYINPUT44), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(KEYINPUT44), .ZN(new_n842));
  AOI21_X1  g656(.A(KEYINPUT45), .B1(new_n621), .B2(new_n624), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n843), .A2(new_n584), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n621), .A2(KEYINPUT45), .A3(new_n814), .A4(new_n816), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(new_n813), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT46), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n786), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n849), .B1(new_n848), .B2(new_n847), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(new_n819), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n851), .A2(new_n759), .A3(new_n811), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n841), .A2(new_n842), .A3(new_n852), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(G137), .ZN(G39));
  INV_X1    g668(.A(KEYINPUT47), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n850), .A2(KEYINPUT47), .A3(new_n819), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n768), .A2(new_n237), .A3(new_n811), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n858), .A2(new_n781), .A3(new_n859), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n860), .B(G140), .ZN(G42));
  INV_X1    g675(.A(KEYINPUT123), .ZN(new_n862));
  NOR2_X1   g676(.A1(G952), .A2(G953), .ZN(new_n863));
  INV_X1    g677(.A(new_n811), .ZN(new_n864));
  OR2_X1    g678(.A1(new_n820), .A2(new_n807), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n865), .A2(new_n779), .A3(new_n780), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n693), .A2(new_n567), .A3(new_n726), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n733), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n864), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n869), .A2(new_n829), .A3(new_n823), .A4(new_n832), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n627), .B1(new_n352), .B2(new_n706), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n442), .A2(new_n681), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n668), .A2(new_n626), .A3(new_n673), .A4(new_n237), .ZN(new_n873));
  OAI22_X1  g687(.A1(new_n872), .A2(new_n873), .B1(new_n799), .B2(new_n802), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n789), .B1(new_n670), .B2(new_n694), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n506), .A2(KEYINPUT20), .A3(new_n508), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n514), .B1(new_n513), .B2(new_n507), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n571), .B(new_n566), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(KEYINPUT113), .ZN(new_n880));
  OAI21_X1  g694(.A(KEYINPUT114), .B1(new_n880), .B2(new_n872), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT113), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n879), .B(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT114), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n883), .A2(new_n884), .A3(new_n442), .A4(new_n681), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n881), .A2(new_n885), .A3(new_n675), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n875), .A2(new_n797), .A3(new_n876), .A4(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT53), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n870), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n809), .B1(new_n732), .B2(new_n736), .ZN(new_n890));
  OR3_X1    g704(.A1(new_n820), .A2(new_n754), .A3(new_n778), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n753), .A2(new_n891), .A3(new_n799), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n892), .B1(new_n777), .B2(new_n782), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n890), .A2(new_n893), .A3(KEYINPUT52), .ZN(new_n894));
  AOI21_X1  g708(.A(KEYINPUT52), .B1(new_n890), .B2(new_n893), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n889), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT116), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n889), .B(KEYINPUT116), .C1(new_n894), .C2(new_n895), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n870), .A2(new_n887), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT52), .ZN(new_n902));
  AOI211_X1 g716(.A(new_n902), .B(new_n892), .C1(new_n777), .C2(new_n782), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n890), .A2(KEYINPUT115), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT115), .ZN(new_n905));
  AOI211_X1 g719(.A(new_n905), .B(new_n809), .C1(new_n732), .C2(new_n736), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n903), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n890), .A2(new_n893), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(new_n902), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n901), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  OAI211_X1 g724(.A(new_n898), .B(new_n899), .C1(new_n910), .C2(KEYINPUT53), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n907), .A2(new_n909), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n900), .B1(new_n894), .B2(new_n895), .ZN(new_n913));
  AOI22_X1  g727(.A1(new_n912), .A2(new_n889), .B1(new_n913), .B2(new_n888), .ZN(new_n914));
  XOR2_X1   g728(.A(KEYINPUT117), .B(KEYINPUT54), .Z(new_n915));
  AOI22_X1  g729(.A1(new_n911), .A2(KEYINPUT54), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n795), .A2(new_n811), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n753), .A2(new_n237), .A3(new_n575), .A4(new_n917), .ZN(new_n918));
  NOR4_X1   g732(.A1(new_n918), .A2(new_n770), .A3(new_n771), .A4(new_n633), .ZN(new_n919));
  OR3_X1    g733(.A1(new_n785), .A2(new_n786), .A3(KEYINPUT118), .ZN(new_n920));
  OAI21_X1  g734(.A(KEYINPUT118), .B1(new_n785), .B2(new_n786), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n920), .A2(new_n583), .A3(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n856), .A2(new_n857), .A3(new_n922), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n801), .A2(new_n237), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n836), .A2(new_n575), .A3(new_n924), .A4(new_n837), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n925), .A2(new_n811), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n919), .B1(new_n923), .B2(new_n926), .ZN(new_n927));
  OR3_X1    g741(.A1(new_n764), .A2(new_n353), .A3(new_n795), .ZN(new_n928));
  NOR2_X1   g742(.A1(KEYINPUT119), .A2(KEYINPUT50), .ZN(new_n929));
  OR3_X1    g743(.A1(new_n928), .A2(new_n925), .A3(new_n929), .ZN(new_n930));
  AND2_X1   g744(.A1(KEYINPUT119), .A2(KEYINPUT50), .ZN(new_n931));
  OAI22_X1  g745(.A1(new_n928), .A2(new_n925), .B1(new_n931), .B2(new_n929), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n836), .A2(new_n575), .A3(new_n837), .A4(new_n917), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT121), .ZN(new_n935));
  OR2_X1    g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n934), .A2(new_n935), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n808), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n927), .A2(new_n933), .A3(KEYINPUT51), .A4(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT48), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n826), .B1(KEYINPUT122), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n942), .B1(new_n936), .B2(new_n937), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n941), .A2(KEYINPUT122), .ZN(new_n944));
  OR2_X1    g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n796), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n661), .A2(new_n669), .ZN(new_n947));
  OAI221_X1 g761(.A(new_n572), .B1(new_n925), .B2(new_n946), .C1(new_n947), .C2(new_n918), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n948), .B1(new_n943), .B2(new_n944), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n940), .A2(new_n945), .A3(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT120), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n933), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n930), .A2(KEYINPUT120), .A3(new_n932), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n952), .A2(new_n953), .A3(new_n939), .A4(new_n927), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT51), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n950), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n863), .B1(new_n916), .B2(new_n956), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n785), .A2(new_n786), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT49), .ZN(new_n959));
  OR3_X1    g773(.A1(new_n236), .A2(new_n354), .A3(new_n583), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n960), .A2(new_n659), .A3(new_n770), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n753), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n962), .A2(new_n764), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n963), .B(KEYINPUT112), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n862), .B1(new_n957), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n898), .A2(new_n899), .ZN(new_n966));
  AOI21_X1  g780(.A(KEYINPUT53), .B1(new_n912), .B2(new_n900), .ZN(new_n967));
  OAI21_X1  g781(.A(KEYINPUT54), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n914), .A2(new_n915), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n968), .A2(new_n969), .A3(new_n956), .ZN(new_n970));
  INV_X1    g784(.A(new_n863), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(new_n964), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n972), .A2(KEYINPUT123), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n965), .A2(new_n974), .ZN(G75));
  NOR2_X1   g789(.A1(new_n447), .A2(G952), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n914), .A2(new_n224), .ZN(new_n978));
  AOI21_X1  g792(.A(KEYINPUT56), .B1(new_n978), .B2(G210), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n412), .A2(new_n418), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n980), .A2(new_n439), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n981), .B(KEYINPUT55), .Z(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n977), .B1(new_n979), .B2(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n984), .B1(new_n979), .B2(new_n983), .ZN(G51));
  NAND2_X1  g799(.A1(new_n611), .A2(new_n617), .ZN(new_n986));
  AND2_X1   g800(.A1(new_n914), .A2(new_n915), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n914), .A2(new_n915), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n585), .B(KEYINPUT57), .Z(new_n990));
  OAI21_X1  g804(.A(new_n986), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n978), .A2(new_n845), .A3(new_n844), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n976), .B1(new_n991), .B2(new_n992), .ZN(G54));
  NAND3_X1  g807(.A1(new_n978), .A2(KEYINPUT58), .A3(G475), .ZN(new_n994));
  AND2_X1   g808(.A1(new_n994), .A2(new_n506), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n994), .A2(new_n506), .ZN(new_n996));
  NOR3_X1   g810(.A1(new_n995), .A2(new_n996), .A3(new_n976), .ZN(G60));
  INV_X1    g811(.A(new_n657), .ZN(new_n998));
  NAND2_X1  g812(.A1(G478), .A2(G902), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT59), .Z(new_n1000));
  OR2_X1    g814(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n977), .B1(new_n989), .B2(new_n1001), .ZN(new_n1002));
  OR2_X1    g816(.A1(new_n916), .A2(new_n1000), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n1002), .B1(new_n998), .B2(new_n1003), .ZN(G63));
  INV_X1    g818(.A(KEYINPUT61), .ZN(new_n1005));
  NAND2_X1  g819(.A1(G217), .A2(G902), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1006), .B(KEYINPUT60), .ZN(new_n1007));
  OAI21_X1  g821(.A(KEYINPUT124), .B1(new_n914), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n223), .A2(new_n225), .ZN(new_n1009));
  INV_X1    g823(.A(KEYINPUT124), .ZN(new_n1010));
  INV_X1    g824(.A(new_n1007), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n903), .A2(new_n890), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1012), .A2(new_n909), .ZN(new_n1013));
  AOI21_X1  g827(.A(KEYINPUT53), .B1(new_n1013), .B2(new_n900), .ZN(new_n1014));
  INV_X1    g828(.A(new_n889), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1015), .B1(new_n907), .B2(new_n909), .ZN(new_n1016));
  OAI211_X1 g830(.A(new_n1010), .B(new_n1011), .C1(new_n1014), .C2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n1008), .A2(new_n1009), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1018), .A2(new_n977), .ZN(new_n1019));
  INV_X1    g833(.A(new_n700), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n1020), .B1(new_n1008), .B2(new_n1017), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1005), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1008), .A2(new_n1017), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1023), .A2(new_n700), .ZN(new_n1024));
  NAND4_X1  g838(.A1(new_n1024), .A2(KEYINPUT61), .A3(new_n977), .A4(new_n1018), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1022), .A2(new_n1025), .ZN(G66));
  OAI21_X1  g840(.A(G953), .B1(new_n578), .B2(new_n415), .ZN(new_n1027));
  INV_X1    g841(.A(new_n887), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n1027), .B1(new_n1028), .B2(G953), .ZN(new_n1029));
  OAI211_X1 g843(.A(new_n408), .B(new_n411), .C1(G898), .C2(new_n447), .ZN(new_n1030));
  XNOR2_X1  g844(.A(new_n1030), .B(KEYINPUT126), .ZN(new_n1031));
  XOR2_X1   g845(.A(new_n1031), .B(KEYINPUT125), .Z(new_n1032));
  XNOR2_X1  g846(.A(new_n1029), .B(new_n1032), .ZN(G69));
  NAND2_X1  g847(.A1(new_n316), .A2(new_n318), .ZN(new_n1034));
  OR2_X1    g848(.A1(new_n484), .A2(new_n485), .ZN(new_n1035));
  XOR2_X1   g849(.A(new_n1034), .B(new_n1035), .Z(new_n1036));
  NOR2_X1   g850(.A1(new_n1036), .A2(G953), .ZN(new_n1037));
  INV_X1    g851(.A(new_n1037), .ZN(new_n1038));
  OR2_X1    g852(.A1(new_n904), .A2(new_n906), .ZN(new_n1039));
  NAND3_X1  g853(.A1(new_n1039), .A2(new_n765), .A3(new_n783), .ZN(new_n1040));
  INV_X1    g854(.A(KEYINPUT62), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND4_X1  g856(.A1(new_n1039), .A2(KEYINPUT62), .A3(new_n765), .A4(new_n783), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g858(.A1(new_n853), .A2(new_n860), .ZN(new_n1045));
  OAI21_X1  g859(.A(new_n880), .B1(new_n660), .B2(new_n659), .ZN(new_n1046));
  NOR3_X1   g860(.A1(new_n761), .A2(new_n352), .A3(new_n811), .ZN(new_n1047));
  AOI21_X1  g861(.A(new_n1045), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g862(.A(new_n1038), .B1(new_n1044), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g863(.A(new_n1049), .ZN(new_n1050));
  NAND2_X1  g864(.A1(new_n1036), .A2(new_n722), .ZN(new_n1051));
  NOR2_X1   g865(.A1(new_n851), .A2(new_n759), .ZN(new_n1052));
  NAND4_X1  g866(.A1(new_n1052), .A2(new_n680), .A3(new_n755), .A4(new_n826), .ZN(new_n1053));
  NAND4_X1  g867(.A1(new_n1053), .A2(new_n829), .A3(new_n823), .A4(new_n832), .ZN(new_n1054));
  NOR2_X1   g868(.A1(new_n1045), .A2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g869(.A1(new_n1055), .A2(new_n783), .A3(new_n1039), .ZN(new_n1056));
  AOI21_X1  g870(.A(new_n1051), .B1(new_n1056), .B2(new_n447), .ZN(new_n1057));
  INV_X1    g871(.A(new_n1057), .ZN(new_n1058));
  INV_X1    g872(.A(G900), .ZN(new_n1059));
  OAI21_X1  g873(.A(G953), .B1(new_n605), .B2(new_n1059), .ZN(new_n1060));
  NAND4_X1  g874(.A1(new_n1050), .A2(new_n1058), .A3(KEYINPUT127), .A4(new_n1060), .ZN(new_n1061));
  NAND2_X1  g875(.A1(new_n1060), .A2(KEYINPUT127), .ZN(new_n1062));
  OR2_X1    g876(.A1(new_n1060), .A2(KEYINPUT127), .ZN(new_n1063));
  OAI211_X1 g877(.A(new_n1062), .B(new_n1063), .C1(new_n1049), .C2(new_n1057), .ZN(new_n1064));
  AND2_X1   g878(.A1(new_n1061), .A2(new_n1064), .ZN(G72));
  NAND2_X1  g879(.A1(G472), .A2(G902), .ZN(new_n1066));
  XOR2_X1   g880(.A(new_n1066), .B(KEYINPUT63), .Z(new_n1067));
  OAI21_X1  g881(.A(new_n1067), .B1(new_n1056), .B2(new_n887), .ZN(new_n1068));
  NOR2_X1   g882(.A1(new_n745), .A2(new_n313), .ZN(new_n1069));
  AOI21_X1  g883(.A(new_n976), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g884(.A(new_n911), .ZN(new_n1071));
  INV_X1    g885(.A(new_n320), .ZN(new_n1072));
  OAI21_X1  g886(.A(new_n1067), .B1(new_n1072), .B2(new_n340), .ZN(new_n1073));
  OAI21_X1  g887(.A(new_n1070), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g888(.A1(new_n1044), .A2(new_n1028), .A3(new_n1048), .ZN(new_n1075));
  AOI21_X1  g889(.A(new_n746), .B1(new_n1075), .B2(new_n1067), .ZN(new_n1076));
  NOR2_X1   g890(.A1(new_n1074), .A2(new_n1076), .ZN(G57));
endmodule


