//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 0 0 0 0 1 1 0 0 1 0 1 1 0 0 1 0 0 0 0 1 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 0 0 0 1 0 0 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n755, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n819, new_n821,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n862, new_n863, new_n864, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n874, new_n876, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928;
  XNOR2_X1  g000(.A(G127gat), .B(G155gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(G231gat), .A2(G233gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(G57gat), .B(G64gat), .Z(new_n206));
  INV_X1    g005(.A(KEYINPUT99), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G71gat), .ZN(new_n209));
  INV_X1    g008(.A(G78gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n209), .A2(new_n210), .A3(KEYINPUT9), .ZN(new_n211));
  NAND2_X1  g010(.A1(G71gat), .A2(G78gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G57gat), .B(G64gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT99), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n208), .A2(new_n213), .A3(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT100), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n216), .B(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n212), .B(KEYINPUT98), .ZN(new_n219));
  AOI21_X1  g018(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n220));
  OAI221_X1 g019(.A(new_n219), .B1(G71gat), .B2(G78gat), .C1(new_n214), .C2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n222), .B(KEYINPUT101), .ZN(new_n223));
  OR2_X1    g022(.A1(new_n223), .A2(KEYINPUT21), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n224), .B(G211gat), .ZN(new_n225));
  XNOR2_X1  g024(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n223), .A2(KEYINPUT21), .ZN(new_n227));
  XNOR2_X1  g026(.A(G15gat), .B(G22gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT16), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n228), .B1(new_n229), .B2(G1gat), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n230), .B1(G1gat), .B2(new_n228), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n231), .B(G8gat), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n227), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(G183gat), .ZN(new_n235));
  INV_X1    g034(.A(G183gat), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n227), .A2(new_n236), .A3(new_n233), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n226), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n235), .A2(new_n237), .A3(new_n226), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n225), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n240), .ZN(new_n242));
  INV_X1    g041(.A(G211gat), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n224), .B(new_n243), .ZN(new_n244));
  NOR3_X1   g043(.A1(new_n242), .A2(new_n238), .A3(new_n244), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n205), .B1(new_n241), .B2(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n244), .B1(new_n242), .B2(new_n238), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n239), .A2(new_n240), .A3(new_n225), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n247), .A2(new_n248), .A3(new_n204), .ZN(new_n249));
  AND2_X1   g048(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(G190gat), .B(G218gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n251), .B(G162gat), .ZN(new_n252));
  AND2_X1   g051(.A1(G232gat), .A2(G233gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(G85gat), .A2(G92gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n254), .B(KEYINPUT103), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n255), .B(KEYINPUT7), .ZN(new_n256));
  XNOR2_X1  g055(.A(KEYINPUT104), .B(G92gat), .ZN(new_n257));
  INV_X1    g056(.A(G85gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(G99gat), .A2(G106gat), .ZN(new_n259));
  AOI22_X1  g058(.A1(new_n257), .A2(new_n258), .B1(KEYINPUT8), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n256), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(G99gat), .B(G106gat), .ZN(new_n262));
  XOR2_X1   g061(.A(new_n261), .B(new_n262), .Z(new_n263));
  INV_X1    g062(.A(G29gat), .ZN(new_n264));
  INV_X1    g063(.A(G36gat), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NOR2_X1   g065(.A1(G29gat), .A2(G36gat), .ZN(new_n267));
  AND2_X1   g066(.A1(KEYINPUT93), .A2(KEYINPUT14), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G43gat), .B(G50gat), .ZN(new_n270));
  OAI22_X1  g069(.A1(KEYINPUT93), .A2(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n271));
  OAI221_X1 g070(.A(new_n269), .B1(KEYINPUT15), .B2(new_n270), .C1(new_n268), .C2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n270), .A2(KEYINPUT15), .ZN(new_n273));
  XOR2_X1   g072(.A(new_n272), .B(new_n273), .Z(new_n274));
  INV_X1    g073(.A(KEYINPUT17), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n272), .B(new_n273), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT17), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n263), .A2(new_n276), .A3(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n261), .B(new_n262), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(new_n274), .ZN(new_n281));
  AOI211_X1 g080(.A(KEYINPUT41), .B(new_n253), .C1(new_n279), .C2(new_n281), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n253), .A2(KEYINPUT41), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n253), .A2(KEYINPUT41), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n279), .A2(new_n284), .A3(new_n285), .A4(new_n281), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n252), .B1(new_n282), .B2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(KEYINPUT102), .B(G134gat), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n279), .A2(new_n285), .A3(new_n281), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(new_n283), .ZN(new_n291));
  INV_X1    g090(.A(new_n252), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n291), .A2(new_n292), .A3(new_n286), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n288), .A2(new_n289), .A3(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n289), .B1(new_n288), .B2(new_n293), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n250), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT101), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n222), .B(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(new_n263), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n280), .A2(new_n218), .A3(new_n221), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(G230gat), .A2(G233gat), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  XOR2_X1   g106(.A(new_n307), .B(KEYINPUT106), .Z(new_n308));
  INV_X1    g107(.A(KEYINPUT10), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n302), .A2(new_n309), .A3(new_n303), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n223), .A2(KEYINPUT10), .A3(new_n280), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT105), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT105), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n310), .A2(new_n314), .A3(new_n311), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n313), .A2(new_n305), .A3(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(KEYINPUT107), .B(G120gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n317), .B(G148gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(G176gat), .B(G204gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n318), .B(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n308), .A2(new_n316), .A3(new_n320), .ZN(new_n321));
  XOR2_X1   g120(.A(new_n320), .B(KEYINPUT108), .Z(new_n322));
  INV_X1    g121(.A(new_n307), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n306), .B1(new_n310), .B2(new_n311), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n299), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n276), .A2(new_n233), .A3(new_n278), .ZN(new_n329));
  NAND2_X1  g128(.A1(G229gat), .A2(G233gat), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n233), .A2(new_n277), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n329), .A2(KEYINPUT18), .A3(new_n330), .A4(new_n332), .ZN(new_n333));
  XOR2_X1   g132(.A(new_n330), .B(KEYINPUT13), .Z(new_n334));
  NOR2_X1   g133(.A1(new_n274), .A2(new_n232), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n334), .B1(new_n335), .B2(new_n331), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT95), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  OAI211_X1 g137(.A(KEYINPUT95), .B(new_n334), .C1(new_n335), .C2(new_n331), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n333), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT96), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n329), .A2(new_n330), .A3(new_n332), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT18), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT94), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n343), .A2(KEYINPUT94), .A3(new_n344), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n333), .A2(new_n338), .A3(KEYINPUT96), .A4(new_n339), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n342), .A2(new_n347), .A3(new_n348), .A4(new_n349), .ZN(new_n350));
  XOR2_X1   g149(.A(G113gat), .B(G141gat), .Z(new_n351));
  XNOR2_X1  g150(.A(new_n351), .B(G197gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(KEYINPUT11), .B(G169gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n352), .B(new_n353), .ZN(new_n354));
  XOR2_X1   g153(.A(new_n354), .B(KEYINPUT12), .Z(new_n355));
  NAND2_X1  g154(.A1(new_n350), .A2(new_n355), .ZN(new_n356));
  AND2_X1   g155(.A1(new_n343), .A2(new_n344), .ZN(new_n357));
  OR3_X1    g156(.A1(new_n340), .A2(new_n357), .A3(new_n355), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT35), .ZN(new_n360));
  INV_X1    g159(.A(G190gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(KEYINPUT65), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT65), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(G190gat), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT27), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(new_n236), .ZN(new_n366));
  NAND2_X1  g165(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n367));
  AOI22_X1  g166(.A1(new_n362), .A2(new_n364), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(KEYINPUT66), .B(KEYINPUT28), .ZN(new_n369));
  OAI21_X1  g168(.A(KEYINPUT67), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(KEYINPUT65), .B(G190gat), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n367), .ZN(new_n373));
  NOR2_X1   g172(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT68), .ZN(new_n375));
  NOR3_X1   g174(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(KEYINPUT68), .B1(new_n366), .B2(new_n367), .ZN(new_n377));
  OAI211_X1 g176(.A(KEYINPUT28), .B(new_n372), .C1(new_n376), .C2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n369), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT67), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n373), .A2(new_n374), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n379), .B(new_n380), .C1(new_n381), .C2(new_n371), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n370), .A2(new_n378), .A3(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(G169gat), .ZN(new_n384));
  INV_X1    g183(.A(G176gat), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n384), .A2(new_n385), .A3(KEYINPUT26), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT26), .B1(new_n384), .B2(new_n385), .ZN(new_n387));
  NAND2_X1  g186(.A1(G169gat), .A2(G176gat), .ZN(new_n388));
  AOI22_X1  g187(.A1(new_n387), .A2(new_n388), .B1(G183gat), .B2(G190gat), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n383), .A2(new_n386), .A3(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n384), .A2(new_n385), .A3(KEYINPUT23), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT23), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n392), .B1(G169gat), .B2(G176gat), .ZN(new_n393));
  AND3_X1   g192(.A1(new_n391), .A2(new_n393), .A3(new_n388), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT64), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n397), .B1(new_n371), .B2(G183gat), .ZN(new_n398));
  NAND3_X1  g197(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n399), .B1(new_n395), .B2(new_n396), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n394), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  NOR2_X1   g200(.A1(G183gat), .A2(G190gat), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n395), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(KEYINPUT25), .B1(new_n403), .B2(new_n399), .ZN(new_n404));
  AOI22_X1  g203(.A1(new_n401), .A2(KEYINPUT25), .B1(new_n394), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(G113gat), .B(G120gat), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT69), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT1), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(KEYINPUT69), .B1(new_n407), .B2(KEYINPUT1), .ZN(new_n412));
  XNOR2_X1  g211(.A(G127gat), .B(G134gat), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n413), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n408), .A2(new_n415), .A3(new_n409), .A4(new_n410), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n406), .B(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(G227gat), .ZN(new_n419));
  INV_X1    g218(.A(G233gat), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT33), .ZN(new_n423));
  OAI22_X1  g222(.A1(new_n418), .A2(new_n422), .B1(KEYINPUT32), .B2(new_n423), .ZN(new_n424));
  XOR2_X1   g223(.A(G15gat), .B(G43gat), .Z(new_n425));
  XNOR2_X1  g224(.A(G71gat), .B(G99gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n425), .B(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT32), .ZN(new_n429));
  INV_X1    g228(.A(new_n418), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n429), .B1(new_n430), .B2(new_n421), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n427), .A2(KEYINPUT33), .ZN(new_n432));
  AND3_X1   g231(.A1(new_n431), .A2(KEYINPUT70), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(KEYINPUT70), .B1(new_n431), .B2(new_n432), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n428), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n418), .A2(new_n422), .ZN(new_n436));
  XOR2_X1   g235(.A(new_n436), .B(KEYINPUT34), .Z(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n437), .B(new_n428), .C1(new_n433), .C2(new_n434), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(G162gat), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT80), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT80), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(G162gat), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n443), .A2(new_n445), .A3(G155gat), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT2), .ZN(new_n447));
  INV_X1    g246(.A(G141gat), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n448), .A2(G148gat), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  AND3_X1   g249(.A1(new_n448), .A2(KEYINPUT79), .A3(G148gat), .ZN(new_n451));
  AOI21_X1  g250(.A(KEYINPUT79), .B1(new_n448), .B2(G148gat), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  XNOR2_X1  g252(.A(G155gat), .B(G162gat), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n447), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  NOR2_X1   g254(.A1(G155gat), .A2(G162gat), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT78), .ZN(new_n457));
  XNOR2_X1  g256(.A(new_n456), .B(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(G155gat), .A2(G162gat), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT2), .ZN(new_n460));
  INV_X1    g259(.A(G148gat), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n461), .A2(G141gat), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n460), .B1(new_n449), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n458), .A2(new_n459), .A3(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT3), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n455), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT29), .ZN(new_n467));
  AND2_X1   g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT73), .ZN(new_n469));
  XNOR2_X1  g268(.A(G211gat), .B(G218gat), .ZN(new_n470));
  XNOR2_X1  g269(.A(G197gat), .B(G204gat), .ZN(new_n471));
  NAND2_X1  g270(.A1(G211gat), .A2(G218gat), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT22), .ZN(new_n473));
  AND3_X1   g272(.A1(new_n472), .A2(KEYINPUT71), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(KEYINPUT71), .B1(new_n472), .B2(new_n473), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n470), .B(new_n471), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT72), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n472), .A2(new_n473), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT71), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n472), .A2(KEYINPUT71), .A3(new_n473), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n470), .B1(new_n483), .B2(new_n471), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n478), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n471), .B1(new_n474), .B2(new_n475), .ZN(new_n486));
  INV_X1    g285(.A(new_n470), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n486), .A2(KEYINPUT72), .A3(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n469), .B1(new_n485), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n486), .A2(new_n487), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n491), .A2(new_n477), .A3(new_n476), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n492), .A2(KEYINPUT73), .A3(new_n488), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n468), .B1(new_n490), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n455), .A2(new_n464), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n491), .A2(KEYINPUT84), .A3(new_n476), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n497), .B(new_n467), .C1(KEYINPUT84), .C2(new_n491), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n496), .B1(new_n498), .B2(new_n465), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT83), .B1(new_n494), .B2(new_n499), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n492), .A2(new_n495), .A3(new_n467), .A4(new_n488), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n495), .A2(KEYINPUT3), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT85), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n466), .A2(new_n467), .ZN(new_n506));
  AND3_X1   g305(.A1(new_n492), .A2(KEYINPUT73), .A3(new_n488), .ZN(new_n507));
  AOI21_X1  g306(.A(KEYINPUT73), .B1(new_n492), .B2(new_n488), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n501), .A2(KEYINPUT85), .A3(new_n502), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n505), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(G228gat), .A2(G233gat), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n500), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT83), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n515), .B1(new_n494), .B2(new_n499), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(new_n512), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(G22gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT86), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n514), .A2(G22gat), .A3(new_n517), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(G78gat), .B(G106gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(KEYINPUT31), .B(G50gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n524), .B(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  OR2_X1    g326(.A1(new_n522), .A2(new_n521), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n523), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT87), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n520), .A2(new_n530), .A3(new_n526), .A4(new_n522), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n520), .A2(new_n526), .A3(new_n522), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(KEYINPUT87), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n529), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT88), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n529), .A2(new_n533), .A3(KEYINPUT88), .A4(new_n531), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n441), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n502), .A2(new_n414), .A3(new_n416), .A4(new_n466), .ZN(new_n539));
  NAND2_X1  g338(.A1(G225gat), .A2(G233gat), .ZN(new_n540));
  AOI211_X1 g339(.A(KEYINPUT4), .B(new_n495), .C1(new_n414), .C2(new_n416), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT4), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n542), .B1(new_n496), .B2(new_n417), .ZN(new_n543));
  OAI211_X1 g342(.A(new_n539), .B(new_n540), .C1(new_n541), .C2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT5), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n417), .B(new_n495), .ZN(new_n548));
  OR2_X1    g347(.A1(new_n548), .A2(new_n540), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n545), .B1(new_n549), .B2(new_n544), .ZN(new_n550));
  XNOR2_X1  g349(.A(G1gat), .B(G29gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(new_n258), .ZN(new_n552));
  XNOR2_X1  g351(.A(KEYINPUT0), .B(G57gat), .ZN(new_n553));
  XOR2_X1   g352(.A(new_n552), .B(new_n553), .Z(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NOR3_X1   g354(.A1(new_n547), .A2(new_n550), .A3(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT82), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n556), .A2(new_n557), .A3(KEYINPUT6), .ZN(new_n558));
  AND2_X1   g357(.A1(new_n549), .A2(new_n544), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n554), .B(new_n546), .C1(new_n559), .C2(new_n545), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n555), .B1(new_n547), .B2(new_n550), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT6), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT81), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(KEYINPUT82), .B1(new_n560), .B2(new_n562), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n560), .A2(new_n561), .A3(KEYINPUT81), .A4(new_n562), .ZN(new_n567));
  AND4_X1   g366(.A1(new_n558), .A2(new_n565), .A3(new_n566), .A4(new_n567), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n507), .A2(new_n508), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT74), .ZN(new_n570));
  AND3_X1   g369(.A1(new_n390), .A2(new_n570), .A3(new_n405), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n570), .B1(new_n390), .B2(new_n405), .ZN(new_n572));
  INV_X1    g371(.A(G226gat), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n573), .A2(new_n420), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NOR3_X1   g374(.A1(new_n571), .A2(new_n572), .A3(new_n575), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n574), .A2(KEYINPUT29), .ZN(new_n577));
  AND2_X1   g376(.A1(new_n406), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n569), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n577), .B1(new_n571), .B2(new_n572), .ZN(new_n580));
  INV_X1    g379(.A(new_n406), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(new_n574), .ZN(new_n582));
  INV_X1    g381(.A(new_n569), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n580), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(KEYINPUT75), .B(G64gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(G92gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(G8gat), .B(G36gat), .ZN(new_n587));
  XOR2_X1   g386(.A(new_n586), .B(new_n587), .Z(new_n588));
  NAND3_X1  g387(.A1(new_n579), .A2(new_n584), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(KEYINPUT76), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(KEYINPUT30), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT77), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT76), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n579), .A2(new_n584), .ZN(new_n597));
  INV_X1    g396(.A(new_n588), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(KEYINPUT76), .B1(new_n589), .B2(new_n592), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(KEYINPUT30), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n596), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n568), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n360), .B1(new_n538), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n536), .A2(new_n537), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n566), .A2(new_n558), .A3(new_n563), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(new_n360), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT89), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT30), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n609), .B1(new_n589), .B2(KEYINPUT76), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n599), .B1(new_n610), .B2(new_n600), .ZN(new_n611));
  AOI211_X1 g410(.A(KEYINPUT76), .B(new_n609), .C1(new_n589), .C2(new_n592), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n608), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n596), .A2(KEYINPUT89), .A3(new_n599), .A4(new_n601), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n607), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n441), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n605), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT92), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n538), .A2(KEYINPUT92), .A3(new_n615), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n604), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n605), .ZN(new_n622));
  OR2_X1    g421(.A1(new_n568), .A2(new_n602), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT91), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n539), .B1(new_n541), .B2(new_n543), .ZN(new_n626));
  INV_X1    g425(.A(new_n540), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(KEYINPUT90), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT90), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n626), .A2(new_n630), .A3(new_n627), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT39), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n554), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n633), .B1(new_n548), .B2(new_n540), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n629), .A2(new_n631), .A3(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n625), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT40), .ZN(new_n638));
  OR2_X1    g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n556), .B1(new_n637), .B2(new_n638), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n613), .A2(new_n614), .A3(new_n639), .A4(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n606), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n598), .B1(new_n597), .B2(KEYINPUT37), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n580), .A2(new_n569), .A3(new_n582), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n576), .A2(new_n578), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n644), .B1(new_n645), .B2(new_n569), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT37), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  OR3_X1    g447(.A1(new_n643), .A2(KEYINPUT38), .A3(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n647), .B1(new_n579), .B2(new_n584), .ZN(new_n650));
  OAI21_X1  g449(.A(KEYINPUT38), .B1(new_n643), .B2(new_n650), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n642), .A2(new_n649), .A3(new_n589), .A4(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n605), .A2(new_n641), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT36), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n441), .B(new_n654), .ZN(new_n655));
  AND3_X1   g454(.A1(new_n624), .A2(new_n653), .A3(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n359), .B1(new_n621), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(KEYINPUT97), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT97), .ZN(new_n659));
  OAI211_X1 g458(.A(new_n659), .B(new_n359), .C1(new_n621), .C2(new_n656), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n328), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(new_n568), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g462(.A1(new_n613), .A2(new_n614), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT42), .ZN(new_n667));
  XNOR2_X1  g466(.A(KEYINPUT16), .B(G8gat), .ZN(new_n668));
  OR3_X1    g467(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n666), .A2(G8gat), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n667), .B1(new_n666), .B2(new_n668), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(G1325gat));
  AOI21_X1  g471(.A(G15gat), .B1(new_n661), .B2(new_n616), .ZN(new_n673));
  INV_X1    g472(.A(new_n655), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n674), .A2(G15gat), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n673), .B1(new_n661), .B2(new_n675), .ZN(G1326gat));
  XNOR2_X1  g475(.A(KEYINPUT43), .B(G22gat), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT109), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n661), .A2(new_n679), .A3(new_n622), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n679), .B1(new_n661), .B2(new_n622), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n678), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n682), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n684), .A2(new_n680), .A3(new_n677), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n683), .A2(new_n685), .ZN(G1327gat));
  NAND2_X1  g485(.A1(new_n246), .A2(new_n249), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n687), .A2(new_n326), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(new_n298), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n689), .B1(new_n658), .B2(new_n660), .ZN(new_n690));
  AND3_X1   g489(.A1(new_n690), .A2(new_n264), .A3(new_n568), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(KEYINPUT45), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT45), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n605), .A2(new_n603), .A3(new_n616), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(KEYINPUT35), .ZN(new_n695));
  AND4_X1   g494(.A1(KEYINPUT92), .A2(new_n605), .A3(new_n615), .A4(new_n616), .ZN(new_n696));
  AOI21_X1  g495(.A(KEYINPUT92), .B1(new_n538), .B2(new_n615), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n695), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT110), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n622), .A2(new_n699), .A3(new_n623), .ZN(new_n700));
  OAI21_X1  g499(.A(KEYINPUT110), .B1(new_n605), .B2(new_n603), .ZN(new_n701));
  NAND4_X1  g500(.A1(new_n700), .A2(new_n701), .A3(new_n655), .A4(new_n653), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n297), .B1(new_n698), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n298), .B1(new_n621), .B2(new_n656), .ZN(new_n704));
  MUX2_X1   g503(.A(new_n703), .B(new_n704), .S(KEYINPUT44), .Z(new_n705));
  NAND4_X1  g504(.A1(new_n705), .A2(new_n568), .A3(new_n359), .A4(new_n688), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n693), .B1(new_n706), .B2(G29gat), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n692), .B1(new_n707), .B2(new_n691), .ZN(G1328gat));
  NAND3_X1  g507(.A1(new_n690), .A2(new_n265), .A3(new_n665), .ZN(new_n709));
  OR2_X1    g508(.A1(new_n709), .A2(KEYINPUT46), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n698), .A2(new_n702), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n298), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT44), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  OAI211_X1 g513(.A(KEYINPUT44), .B(new_n298), .C1(new_n621), .C2(new_n656), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n714), .A2(new_n359), .A3(new_n688), .A4(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(G36gat), .B1(new_n716), .B2(new_n664), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n709), .A2(KEYINPUT46), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n710), .A2(new_n717), .A3(new_n718), .ZN(G1329gat));
  OAI21_X1  g518(.A(G43gat), .B1(new_n716), .B2(new_n655), .ZN(new_n720));
  INV_X1    g519(.A(G43gat), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n690), .A2(new_n721), .A3(new_n616), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT111), .ZN(new_n724));
  AOI21_X1  g523(.A(KEYINPUT47), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  OAI211_X1 g525(.A(new_n720), .B(new_n722), .C1(new_n724), .C2(KEYINPUT47), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(G1330gat));
  INV_X1    g527(.A(G50gat), .ZN(new_n729));
  OR3_X1    g528(.A1(new_n716), .A2(new_n729), .A3(new_n605), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT48), .ZN(new_n731));
  AOI21_X1  g530(.A(G50gat), .B1(new_n690), .B2(new_n622), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n730), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n716), .A2(new_n729), .A3(new_n605), .ZN(new_n735));
  OAI21_X1  g534(.A(KEYINPUT48), .B1(new_n735), .B2(new_n732), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n736), .ZN(G1331gat));
  AOI21_X1  g536(.A(new_n359), .B1(new_n698), .B2(new_n702), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n250), .A2(new_n298), .A3(new_n327), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n738), .A2(new_n568), .A3(new_n739), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g540(.A1(new_n738), .A2(new_n739), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n742), .A2(new_n664), .ZN(new_n743));
  NOR2_X1   g542(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n744));
  AND2_X1   g543(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n743), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n746), .B1(new_n743), .B2(new_n744), .ZN(G1333gat));
  OAI21_X1  g546(.A(new_n209), .B1(new_n742), .B2(new_n441), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n738), .A2(G71gat), .A3(new_n674), .A4(new_n739), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT112), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n749), .A2(new_n750), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n748), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g553(.A1(new_n742), .A2(new_n605), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(new_n210), .ZN(G1335gat));
  NOR2_X1   g555(.A1(new_n687), .A2(new_n359), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n711), .A2(new_n298), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(KEYINPUT51), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT51), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n703), .A2(new_n760), .A3(new_n757), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n762), .A2(new_n568), .A3(new_n326), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n687), .A2(new_n327), .A3(new_n359), .ZN(new_n764));
  OAI211_X1 g563(.A(new_n715), .B(new_n764), .C1(KEYINPUT44), .C2(new_n703), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n765), .A2(new_n258), .ZN(new_n766));
  AOI22_X1  g565(.A1(new_n763), .A2(new_n258), .B1(new_n568), .B2(new_n766), .ZN(G1336gat));
  NOR2_X1   g566(.A1(new_n664), .A2(G92gat), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n759), .A2(new_n326), .A3(new_n761), .A4(new_n768), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n765), .A2(new_n664), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n769), .B1(new_n770), .B2(new_n257), .ZN(new_n771));
  XNOR2_X1  g570(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n771), .B(new_n772), .ZN(G1337gat));
  OAI21_X1  g572(.A(G99gat), .B1(new_n765), .B2(new_n655), .ZN(new_n774));
  INV_X1    g573(.A(G99gat), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n762), .A2(new_n775), .A3(new_n326), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n774), .B1(new_n776), .B2(new_n441), .ZN(G1338gat));
  OAI21_X1  g576(.A(G106gat), .B1(new_n765), .B2(new_n605), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT114), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n605), .A2(G106gat), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n759), .A2(new_n326), .A3(new_n761), .A4(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n778), .A2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT53), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n780), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  OAI211_X1 g584(.A(new_n778), .B(new_n782), .C1(new_n779), .C2(KEYINPUT53), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n785), .A2(new_n786), .ZN(G1339gat));
  INV_X1    g586(.A(new_n289), .ZN(new_n788));
  INV_X1    g587(.A(new_n293), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n292), .B1(new_n291), .B2(new_n286), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n356), .A2(new_n358), .A3(new_n791), .A4(new_n294), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n330), .B1(new_n329), .B2(new_n332), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n335), .A2(new_n331), .A3(new_n334), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n354), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n358), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n796), .B1(new_n295), .B2(new_n296), .ZN(new_n797));
  AND3_X1   g596(.A1(new_n792), .A2(new_n797), .A3(new_n321), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT115), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n310), .A2(new_n306), .A3(new_n311), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n316), .A2(KEYINPUT54), .A3(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT54), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n320), .B1(new_n324), .B2(new_n803), .ZN(new_n804));
  AOI211_X1 g603(.A(new_n799), .B(new_n800), .C1(new_n802), .C2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n799), .A2(new_n800), .ZN(new_n806));
  NAND2_X1  g605(.A1(KEYINPUT115), .A2(KEYINPUT55), .ZN(new_n807));
  AND4_X1   g606(.A1(new_n804), .A2(new_n802), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n798), .B1(new_n805), .B2(new_n808), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n326), .A2(new_n358), .A3(new_n297), .A4(new_n795), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n250), .ZN(new_n812));
  INV_X1    g611(.A(new_n359), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n299), .A2(new_n813), .A3(new_n327), .ZN(new_n814));
  AOI211_X1 g613(.A(new_n622), .B(new_n441), .C1(new_n812), .C2(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n815), .A2(new_n568), .A3(new_n664), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n816), .A2(new_n813), .ZN(new_n817));
  XOR2_X1   g616(.A(new_n817), .B(G113gat), .Z(G1340gat));
  NOR2_X1   g617(.A1(new_n816), .A2(new_n327), .ZN(new_n819));
  XOR2_X1   g618(.A(new_n819), .B(G120gat), .Z(G1341gat));
  NOR2_X1   g619(.A1(new_n816), .A2(new_n250), .ZN(new_n821));
  XOR2_X1   g620(.A(new_n821), .B(G127gat), .Z(G1342gat));
  INV_X1    g621(.A(G134gat), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n815), .A2(new_n823), .A3(new_n568), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n664), .A2(new_n298), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(KEYINPUT116), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g626(.A(new_n827), .B(KEYINPUT56), .ZN(new_n828));
  OAI21_X1  g627(.A(G134gat), .B1(new_n816), .B2(new_n297), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n829), .A2(KEYINPUT117), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT117), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n831), .B(G134gat), .C1(new_n816), .C2(new_n297), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n828), .B1(new_n830), .B2(new_n833), .ZN(G1343gat));
  AOI21_X1  g633(.A(new_n687), .B1(new_n809), .B2(new_n810), .ZN(new_n835));
  NOR4_X1   g634(.A1(new_n250), .A2(new_n359), .A3(new_n298), .A4(new_n326), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n622), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(KEYINPUT57), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT57), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n839), .B(new_n622), .C1(new_n835), .C2(new_n836), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n655), .A2(new_n568), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n841), .A2(new_n665), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n838), .A2(new_n359), .A3(new_n840), .A4(new_n842), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n843), .A2(KEYINPUT118), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n843), .A2(KEYINPUT118), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n844), .A2(new_n845), .A3(new_n448), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n837), .A2(new_n665), .A3(new_n841), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n847), .A2(new_n448), .A3(new_n359), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT58), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n843), .A2(G141gat), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n851), .A2(new_n848), .ZN(new_n852));
  OAI22_X1  g651(.A1(new_n846), .A2(new_n850), .B1(new_n849), .B2(new_n852), .ZN(G1344gat));
  NAND3_X1  g652(.A1(new_n847), .A2(new_n461), .A3(new_n326), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n838), .A2(new_n840), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n855), .A2(new_n326), .A3(new_n842), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT119), .ZN(new_n857));
  OAI21_X1  g656(.A(KEYINPUT59), .B1(new_n857), .B2(new_n461), .ZN(new_n858));
  AND3_X1   g657(.A1(new_n856), .A2(G148gat), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n858), .B1(new_n856), .B2(G148gat), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n854), .B1(new_n859), .B2(new_n860), .ZN(G1345gat));
  AOI21_X1  g660(.A(G155gat), .B1(new_n847), .B2(new_n687), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n855), .A2(new_n842), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n863), .A2(new_n250), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n862), .B1(new_n864), .B2(G155gat), .ZN(G1346gat));
  OAI211_X1 g664(.A(new_n443), .B(new_n445), .C1(new_n863), .C2(new_n297), .ZN(new_n866));
  INV_X1    g665(.A(new_n837), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n826), .B1(new_n443), .B2(new_n445), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n867), .A2(new_n568), .A3(new_n655), .A4(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n866), .A2(new_n869), .ZN(G1347gat));
  NOR2_X1   g669(.A1(new_n664), .A2(new_n568), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n815), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n872), .A2(new_n813), .ZN(new_n873));
  XOR2_X1   g672(.A(KEYINPUT120), .B(G169gat), .Z(new_n874));
  XNOR2_X1  g673(.A(new_n873), .B(new_n874), .ZN(G1348gat));
  NOR2_X1   g674(.A1(new_n872), .A2(new_n327), .ZN(new_n876));
  XNOR2_X1  g675(.A(new_n876), .B(new_n385), .ZN(G1349gat));
  NAND3_X1  g676(.A1(new_n815), .A2(new_n687), .A3(new_n871), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(G183gat), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n376), .A2(new_n377), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n879), .B1(new_n880), .B2(new_n878), .ZN(new_n881));
  XNOR2_X1  g680(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  XNOR2_X1  g682(.A(new_n881), .B(new_n883), .ZN(G1350gat));
  OAI21_X1  g683(.A(G190gat), .B1(new_n872), .B2(new_n297), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n885), .A2(KEYINPUT61), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT61), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n872), .A2(new_n297), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n887), .B1(new_n888), .B2(new_n372), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n886), .B1(new_n885), .B2(new_n889), .ZN(G1351gat));
  NAND2_X1  g689(.A1(new_n655), .A2(new_n871), .ZN(new_n891));
  XOR2_X1   g690(.A(new_n891), .B(KEYINPUT122), .Z(new_n892));
  INV_X1    g691(.A(KEYINPUT123), .ZN(new_n893));
  OR2_X1    g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n892), .A2(new_n893), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n855), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  OAI21_X1  g695(.A(KEYINPUT124), .B1(new_n896), .B2(new_n813), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n894), .A2(new_n895), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT124), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n898), .A2(new_n899), .A3(new_n359), .A4(new_n855), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n897), .A2(new_n900), .A3(G197gat), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n837), .A2(new_n891), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  OR3_X1    g702(.A1(new_n903), .A2(G197gat), .A3(new_n813), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n901), .A2(new_n904), .ZN(G1352gat));
  XNOR2_X1  g704(.A(KEYINPUT125), .B(G204gat), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n903), .A2(new_n327), .A3(new_n906), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n907), .B(KEYINPUT62), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n906), .B1(new_n896), .B2(new_n327), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(G1353gat));
  NAND4_X1  g709(.A1(new_n838), .A2(new_n687), .A3(new_n840), .A4(new_n892), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(G211gat), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(KEYINPUT63), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT63), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n911), .A2(new_n914), .A3(G211gat), .ZN(new_n915));
  INV_X1    g714(.A(new_n891), .ZN(new_n916));
  NAND4_X1  g715(.A1(new_n867), .A2(new_n243), .A3(new_n687), .A4(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT126), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n902), .A2(KEYINPUT126), .A3(new_n243), .A4(new_n687), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n913), .A2(new_n915), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(KEYINPUT127), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT127), .ZN(new_n924));
  NAND4_X1  g723(.A1(new_n913), .A2(new_n921), .A3(new_n924), .A4(new_n915), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n923), .A2(new_n925), .ZN(G1354gat));
  AOI21_X1  g725(.A(G218gat), .B1(new_n902), .B2(new_n298), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n896), .A2(new_n297), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n927), .B1(new_n928), .B2(G218gat), .ZN(G1355gat));
endmodule


