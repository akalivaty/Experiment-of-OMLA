//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 1 1 0 1 0 0 1 0 1 1 1 0 0 0 0 0 1 1 1 0 0 0 1 0 0 1 0 1 0 1 1 0 0 0 0 0 1 1 1 0 0 0 1 0 1 0 1 0 1 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:33 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n569, new_n570, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n631, new_n633,
    new_n634, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1175;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(G220));
  XOR2_X1   g012(.A(KEYINPUT66), .B(G96), .Z(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XOR2_X1   g016(.A(KEYINPUT67), .B(G108), .Z(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G219), .A4(G221), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G125), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AND2_X1   g042(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n468));
  NOR2_X1   g043(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n470), .A2(new_n473), .A3(G137), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT70), .ZN(new_n475));
  INV_X1    g050(.A(G2105), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n476), .A2(G101), .A3(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(KEYINPUT69), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT69), .ZN(new_n479));
  NAND4_X1  g054(.A1(new_n479), .A2(new_n476), .A3(G101), .A4(G2104), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  AND3_X1   g056(.A1(new_n474), .A2(new_n475), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n475), .B1(new_n474), .B2(new_n481), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n472), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G160));
  NAND2_X1  g060(.A1(new_n471), .A2(new_n473), .ZN(new_n486));
  INV_X1    g061(.A(G124), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n470), .A2(G112), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n489));
  OAI22_X1  g064(.A1(new_n486), .A2(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n465), .A2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(G136), .ZN(new_n493));
  OR3_X1    g068(.A1(new_n492), .A2(KEYINPUT71), .A3(new_n493), .ZN(new_n494));
  OAI21_X1  g069(.A(KEYINPUT71), .B1(new_n492), .B2(new_n493), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n490), .B1(new_n494), .B2(new_n495), .ZN(G162));
  NAND2_X1  g071(.A1(G126), .A2(G2105), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n476), .A2(G114), .ZN(new_n498));
  OAI21_X1  g073(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n499));
  OAI22_X1  g074(.A1(new_n465), .A2(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT68), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(new_n476), .ZN(new_n502));
  NAND2_X1  g077(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n503));
  OAI211_X1 g078(.A(new_n502), .B(new_n503), .C1(new_n463), .C2(new_n464), .ZN(new_n504));
  INV_X1    g079(.A(G138), .ZN(new_n505));
  OAI21_X1  g080(.A(KEYINPUT4), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT4), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n470), .A2(new_n473), .A3(new_n507), .A4(G138), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n500), .B1(new_n506), .B2(new_n508), .ZN(G164));
  NOR2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT72), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(KEYINPUT72), .A2(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n510), .B1(new_n515), .B2(KEYINPUT6), .ZN(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G50), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT5), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G543), .ZN(new_n521));
  AND3_X1   g096(.A1(new_n517), .A2(KEYINPUT73), .A3(KEYINPUT5), .ZN(new_n522));
  AOI21_X1  g097(.A(KEYINPUT73), .B1(new_n517), .B2(KEYINPUT5), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n516), .A2(new_n524), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT74), .B(G88), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT73), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n528), .B1(new_n520), .B2(G543), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n517), .A2(KEYINPUT73), .A3(KEYINPUT5), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n529), .A2(new_n530), .B1(new_n520), .B2(G543), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n531), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n532));
  INV_X1    g107(.A(new_n515), .ZN(new_n533));
  OAI211_X1 g108(.A(new_n519), .B(new_n527), .C1(new_n532), .C2(new_n533), .ZN(G303));
  INV_X1    g109(.A(G303), .ZN(G166));
  AND2_X1   g110(.A1(G63), .A2(G651), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(KEYINPUT7), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n537), .A2(KEYINPUT7), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n531), .A2(new_n536), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AND2_X1   g115(.A1(KEYINPUT72), .A2(G651), .ZN(new_n541));
  NOR2_X1   g116(.A1(KEYINPUT72), .A2(G651), .ZN(new_n542));
  OAI21_X1  g117(.A(KEYINPUT6), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(new_n510), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G543), .ZN(new_n546));
  XNOR2_X1  g121(.A(KEYINPUT75), .B(G51), .ZN(new_n547));
  INV_X1    g122(.A(G89), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n545), .A2(new_n531), .ZN(new_n549));
  OAI221_X1 g124(.A(new_n540), .B1(new_n546), .B2(new_n547), .C1(new_n548), .C2(new_n549), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n550), .A2(KEYINPUT76), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(KEYINPUT76), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(G168));
  INV_X1    g128(.A(G52), .ZN(new_n554));
  INV_X1    g129(.A(G90), .ZN(new_n555));
  OAI22_X1  g130(.A1(new_n554), .A2(new_n546), .B1(new_n549), .B2(new_n555), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n531), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n557), .A2(new_n533), .ZN(new_n558));
  OR2_X1    g133(.A1(new_n556), .A2(new_n558), .ZN(G301));
  INV_X1    g134(.A(G301), .ZN(G171));
  AOI22_X1  g135(.A1(G43), .A2(new_n518), .B1(new_n525), .B2(G81), .ZN(new_n561));
  NAND2_X1  g136(.A1(G68), .A2(G543), .ZN(new_n562));
  INV_X1    g137(.A(G56), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n524), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(new_n515), .ZN(new_n565));
  AND2_X1   g140(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(G153));
  NAND4_X1  g142(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND4_X1  g145(.A1(G319), .A2(G483), .A3(G661), .A4(new_n570), .ZN(G188));
  NAND3_X1  g146(.A1(new_n545), .A2(G91), .A3(new_n531), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(KEYINPUT79), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT79), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n545), .A2(new_n531), .A3(new_n574), .A4(G91), .ZN(new_n575));
  NAND2_X1  g150(.A1(G78), .A2(G543), .ZN(new_n576));
  INV_X1    g151(.A(G65), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n524), .B2(new_n577), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n573), .A2(new_n575), .B1(G651), .B2(new_n578), .ZN(new_n579));
  AND2_X1   g154(.A1(KEYINPUT77), .A2(G53), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT6), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n581), .B1(new_n513), .B2(new_n514), .ZN(new_n582));
  OAI211_X1 g157(.A(G543), .B(new_n580), .C1(new_n582), .C2(new_n510), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(KEYINPUT9), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT9), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n545), .A2(new_n585), .A3(G543), .A4(new_n580), .ZN(new_n586));
  AND3_X1   g161(.A1(new_n584), .A2(KEYINPUT78), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g162(.A(KEYINPUT78), .B1(new_n584), .B2(new_n586), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n579), .B1(new_n587), .B2(new_n588), .ZN(G299));
  INV_X1    g164(.A(G168), .ZN(G286));
  OAI21_X1  g165(.A(G651), .B1(new_n531), .B2(G74), .ZN(new_n591));
  INV_X1    g166(.A(G49), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n546), .B2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(G87), .ZN(new_n594));
  OR3_X1    g169(.A1(new_n549), .A2(KEYINPUT80), .A3(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(KEYINPUT80), .B1(new_n549), .B2(new_n594), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n593), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G288));
  INV_X1    g173(.A(KEYINPUT82), .ZN(new_n599));
  NAND2_X1  g174(.A1(G48), .A2(G543), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n516), .B2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n600), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n545), .A2(KEYINPUT82), .A3(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n601), .A2(new_n603), .B1(new_n525), .B2(G86), .ZN(new_n604));
  OAI211_X1 g179(.A(G61), .B(new_n521), .C1(new_n522), .C2(new_n523), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT81), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n605), .A2(new_n606), .B1(G73), .B2(G543), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n531), .A2(KEYINPUT81), .A3(G61), .ZN(new_n608));
  AND2_X1   g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n604), .B1(new_n609), .B2(new_n533), .ZN(G305));
  INV_X1    g185(.A(G47), .ZN(new_n611));
  INV_X1    g186(.A(G85), .ZN(new_n612));
  OAI22_X1  g187(.A1(new_n611), .A2(new_n546), .B1(new_n549), .B2(new_n612), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT83), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n531), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n615));
  OR2_X1    g190(.A1(new_n615), .A2(new_n533), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n614), .A2(new_n616), .ZN(G290));
  NAND2_X1  g192(.A1(G301), .A2(G868), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n525), .A2(G92), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(KEYINPUT10), .Z(new_n620));
  NAND2_X1  g195(.A1(G79), .A2(G543), .ZN(new_n621));
  INV_X1    g196(.A(G66), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n524), .B2(new_n622), .ZN(new_n623));
  AOI22_X1  g198(.A1(G54), .A2(new_n518), .B1(new_n623), .B2(G651), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n618), .B1(new_n626), .B2(G868), .ZN(G284));
  OAI21_X1  g202(.A(new_n618), .B1(new_n626), .B2(G868), .ZN(G321));
  MUX2_X1   g203(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g204(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g205(.A(G559), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n626), .B1(new_n631), .B2(G860), .ZN(G148));
  NAND2_X1  g207(.A1(new_n626), .A2(new_n631), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(G868), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(G868), .B2(new_n566), .ZN(G323));
  XNOR2_X1  g210(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g211(.A(G111), .ZN(new_n637));
  INV_X1    g212(.A(KEYINPUT85), .ZN(new_n638));
  OAI21_X1  g213(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n639));
  AOI22_X1  g214(.A1(new_n471), .A2(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n640), .B1(new_n638), .B2(new_n639), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n491), .A2(G135), .ZN(new_n642));
  INV_X1    g217(.A(G123), .ZN(new_n643));
  OAI211_X1 g218(.A(new_n641), .B(new_n642), .C1(new_n643), .C2(new_n486), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT86), .B(G2096), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n476), .A2(G2104), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n473), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT13), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n652), .A2(G2100), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(G2100), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n646), .A2(new_n653), .A3(new_n654), .ZN(G156));
  XNOR2_X1  g230(.A(KEYINPUT15), .B(G2435), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(G2438), .Z(new_n657));
  XNOR2_X1  g232(.A(G2427), .B(G2430), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g234(.A(KEYINPUT14), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(KEYINPUT87), .Z(new_n661));
  INV_X1    g236(.A(new_n657), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n661), .B1(new_n662), .B2(new_n658), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2443), .B(G2446), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1341), .B(G1348), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n665), .B(new_n666), .Z(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G2451), .B(G2454), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT16), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT88), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  OAI21_X1  g247(.A(G14), .B1(new_n668), .B2(new_n672), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(new_n672), .B2(new_n668), .ZN(G401));
  INV_X1    g249(.A(KEYINPUT18), .ZN(new_n675));
  XOR2_X1   g250(.A(G2084), .B(G2090), .Z(new_n676));
  XNOR2_X1  g251(.A(G2067), .B(G2678), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n678), .A2(KEYINPUT17), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n676), .A2(new_n677), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n675), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(G2100), .ZN(new_n682));
  XOR2_X1   g257(.A(G2072), .B(G2078), .Z(new_n683));
  AOI21_X1  g258(.A(new_n683), .B1(new_n678), .B2(KEYINPUT18), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(G2096), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n682), .B(new_n685), .ZN(G227));
  XOR2_X1   g261(.A(G1956), .B(G2474), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT89), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1961), .B(G1966), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1971), .B(G1976), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT19), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(KEYINPUT20), .Z(new_n695));
  NOR2_X1   g270(.A1(new_n688), .A2(new_n690), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n697), .A2(new_n693), .A3(new_n691), .ZN(new_n698));
  OAI211_X1 g273(.A(new_n695), .B(new_n698), .C1(new_n693), .C2(new_n697), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1991), .B(G1996), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XOR2_X1   g278(.A(G1981), .B(G1986), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(G229));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G24), .ZN(new_n708));
  INV_X1    g283(.A(G290), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n708), .B1(new_n709), .B2(new_n707), .ZN(new_n710));
  INV_X1    g285(.A(G1986), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  AND2_X1   g287(.A1(new_n712), .A2(KEYINPUT90), .ZN(new_n713));
  OAI221_X1 g288(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n470), .C2(G107), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n491), .A2(G131), .ZN(new_n715));
  INV_X1    g290(.A(G119), .ZN(new_n716));
  OAI211_X1 g291(.A(new_n714), .B(new_n715), .C1(new_n716), .C2(new_n486), .ZN(new_n717));
  MUX2_X1   g292(.A(G25), .B(new_n717), .S(G29), .Z(new_n718));
  XOR2_X1   g293(.A(KEYINPUT35), .B(G1991), .Z(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n718), .B(new_n720), .ZN(new_n721));
  NOR3_X1   g296(.A1(new_n713), .A2(KEYINPUT91), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n707), .A2(G22), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G166), .B2(new_n707), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(G1971), .Z(new_n725));
  NOR2_X1   g300(.A1(new_n597), .A2(new_n707), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(new_n707), .B2(G23), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT33), .B(G1976), .Z(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n727), .A2(new_n729), .ZN(new_n731));
  NOR2_X1   g306(.A1(G6), .A2(G16), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n533), .B1(new_n607), .B2(new_n608), .ZN(new_n733));
  AOI21_X1  g308(.A(KEYINPUT82), .B1(new_n545), .B2(new_n602), .ZN(new_n734));
  AOI211_X1 g309(.A(new_n599), .B(new_n600), .C1(new_n543), .C2(new_n544), .ZN(new_n735));
  INV_X1    g310(.A(G86), .ZN(new_n736));
  OAI22_X1  g311(.A1(new_n734), .A2(new_n735), .B1(new_n736), .B2(new_n549), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n733), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n732), .B1(new_n738), .B2(G16), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT32), .B(G1981), .Z(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NAND4_X1  g316(.A1(new_n725), .A2(new_n730), .A3(new_n731), .A4(new_n741), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT34), .Z(new_n743));
  OAI211_X1 g318(.A(new_n722), .B(new_n743), .C1(KEYINPUT90), .C2(new_n712), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT36), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n744), .A2(new_n745), .ZN(new_n747));
  INV_X1    g322(.A(G29), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(G32), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n648), .A2(G105), .ZN(new_n750));
  NAND3_X1  g325(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT26), .Z(new_n752));
  INV_X1    g327(.A(G129), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n752), .B1(new_n486), .B2(new_n753), .ZN(new_n754));
  AOI211_X1 g329(.A(new_n750), .B(new_n754), .C1(G141), .C2(new_n491), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n749), .B1(new_n755), .B2(new_n748), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT27), .ZN(new_n757));
  INV_X1    g332(.A(G1996), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  AND2_X1   g334(.A1(new_n748), .A2(G33), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT25), .Z(new_n762));
  NAND2_X1  g337(.A1(new_n491), .A2(G139), .ZN(new_n763));
  AOI22_X1  g338(.A1(new_n473), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n764));
  OAI211_X1 g339(.A(new_n762), .B(new_n763), .C1(new_n470), .C2(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n760), .B1(new_n765), .B2(G29), .ZN(new_n766));
  INV_X1    g341(.A(G2072), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT94), .Z(new_n769));
  NOR2_X1   g344(.A1(new_n759), .A2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(G34), .ZN(new_n771));
  AOI21_X1  g346(.A(G29), .B1(new_n771), .B2(KEYINPUT24), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(KEYINPUT24), .B2(new_n771), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(new_n484), .B2(new_n748), .ZN(new_n774));
  INV_X1    g349(.A(G2084), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n748), .A2(G26), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT28), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n471), .A2(new_n473), .A3(G128), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT93), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n470), .A2(G116), .ZN(new_n781));
  OAI21_X1  g356(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  AOI22_X1  g358(.A1(new_n781), .A2(new_n783), .B1(new_n491), .B2(G140), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n780), .A2(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n778), .B1(new_n786), .B2(new_n748), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G2067), .ZN(new_n788));
  INV_X1    g363(.A(G1961), .ZN(new_n789));
  NOR2_X1   g364(.A1(G171), .A2(new_n707), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G5), .B2(new_n707), .ZN(new_n791));
  AOI211_X1 g366(.A(new_n776), .B(new_n788), .C1(new_n789), .C2(new_n791), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT31), .B(G11), .Z(new_n793));
  NOR2_X1   g368(.A1(new_n644), .A2(new_n748), .ZN(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT30), .B(G28), .ZN(new_n795));
  AOI211_X1 g370(.A(new_n793), .B(new_n794), .C1(new_n748), .C2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n766), .A2(new_n767), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n748), .A2(G27), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G164), .B2(new_n748), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n799), .A2(G2078), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(G2078), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n796), .A2(new_n797), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(G2090), .ZN(new_n803));
  INV_X1    g378(.A(G35), .ZN(new_n804));
  OR3_X1    g379(.A1(new_n804), .A2(KEYINPUT95), .A3(G29), .ZN(new_n805));
  OAI21_X1  g380(.A(KEYINPUT95), .B1(new_n804), .B2(G29), .ZN(new_n806));
  OAI211_X1 g381(.A(new_n805), .B(new_n806), .C1(G162), .C2(new_n748), .ZN(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT96), .B(KEYINPUT29), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n802), .B1(new_n803), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n566), .A2(new_n707), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n707), .B2(G19), .ZN(new_n813));
  INV_X1    g388(.A(G1341), .ZN(new_n814));
  OAI22_X1  g389(.A1(new_n791), .A2(new_n789), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(new_n814), .B2(new_n813), .ZN(new_n816));
  NAND4_X1  g391(.A1(new_n770), .A2(new_n792), .A3(new_n811), .A4(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n626), .A2(G16), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(G4), .B2(G16), .ZN(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT92), .B(G1348), .ZN(new_n820));
  AOI22_X1  g395(.A1(new_n819), .A2(new_n820), .B1(G2090), .B2(new_n809), .ZN(new_n821));
  NOR2_X1   g396(.A1(G16), .A2(G21), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(G168), .B2(G16), .ZN(new_n823));
  INV_X1    g398(.A(G1966), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  OAI211_X1 g400(.A(new_n821), .B(new_n825), .C1(new_n819), .C2(new_n820), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n707), .A2(G20), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT23), .ZN(new_n828));
  INV_X1    g403(.A(G299), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n828), .B1(new_n829), .B2(new_n707), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(G1956), .ZN(new_n831));
  NOR3_X1   g406(.A1(new_n817), .A2(new_n826), .A3(new_n831), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n746), .A2(new_n747), .A3(new_n832), .ZN(G150));
  INV_X1    g408(.A(G150), .ZN(G311));
  NOR2_X1   g409(.A1(new_n625), .A2(new_n631), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT38), .ZN(new_n836));
  AOI22_X1  g411(.A1(G55), .A2(new_n518), .B1(new_n525), .B2(G93), .ZN(new_n837));
  AOI22_X1  g412(.A1(new_n531), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n838));
  OR2_X1    g413(.A1(new_n838), .A2(new_n533), .ZN(new_n839));
  AND2_X1   g414(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n566), .B(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n836), .B(new_n841), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n842), .A2(KEYINPUT39), .ZN(new_n843));
  INV_X1    g418(.A(G860), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n842), .A2(KEYINPUT39), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n840), .A2(new_n844), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT37), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(new_n848), .ZN(G145));
  NAND2_X1  g424(.A1(new_n506), .A2(new_n508), .ZN(new_n850));
  INV_X1    g425(.A(new_n500), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT97), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(new_n765), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n717), .B(new_n651), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n786), .B(new_n755), .ZN(new_n857));
  OAI221_X1 g432(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n470), .C2(G118), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n491), .A2(G142), .ZN(new_n859));
  INV_X1    g434(.A(G130), .ZN(new_n860));
  OAI211_X1 g435(.A(new_n858), .B(new_n859), .C1(new_n860), .C2(new_n486), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n857), .B(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n856), .B(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(G160), .B(new_n644), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(G162), .ZN(new_n865));
  AOI21_X1  g440(.A(G37), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n866), .B1(new_n865), .B2(new_n863), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g443(.A1(new_n625), .A2(G299), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n625), .A2(G299), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  OR2_X1    g448(.A1(new_n873), .A2(KEYINPUT41), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n633), .B(new_n841), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n873), .A2(KEYINPUT41), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n874), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n878), .A2(KEYINPUT99), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(KEYINPUT99), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT98), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n872), .B(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(new_n875), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n879), .A2(new_n880), .A3(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n597), .B(KEYINPUT100), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(G305), .ZN(new_n886));
  XNOR2_X1  g461(.A(G290), .B(G166), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n886), .B(new_n887), .ZN(new_n888));
  XOR2_X1   g463(.A(new_n888), .B(KEYINPUT42), .Z(new_n889));
  XNOR2_X1  g464(.A(new_n884), .B(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(G868), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n891), .B1(G868), .B2(new_n840), .ZN(G295));
  OAI21_X1  g467(.A(new_n891), .B1(G868), .B2(new_n840), .ZN(G331));
  XNOR2_X1  g468(.A(G168), .B(G301), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(new_n841), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n896), .A2(new_n874), .A3(new_n877), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n895), .A2(new_n873), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n897), .A2(new_n888), .A3(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(G37), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n888), .B1(new_n897), .B2(new_n898), .ZN(new_n902));
  OAI21_X1  g477(.A(KEYINPUT43), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT101), .ZN(new_n904));
  OR2_X1    g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI22_X1  g480(.A1(new_n897), .A2(KEYINPUT102), .B1(new_n882), .B2(new_n895), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n906), .B1(KEYINPUT102), .B2(new_n897), .ZN(new_n907));
  INV_X1    g482(.A(new_n888), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n901), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT43), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n903), .A2(new_n904), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n905), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI211_X1 g490(.A(new_n910), .B(new_n901), .C1(new_n907), .C2(new_n908), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n901), .A2(new_n902), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n917), .A2(KEYINPUT43), .ZN(new_n918));
  OAI21_X1  g493(.A(KEYINPUT44), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n915), .A2(new_n919), .ZN(G397));
  INV_X1    g495(.A(G1384), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n852), .A2(new_n921), .ZN(new_n922));
  OAI211_X1 g497(.A(G40), .B(new_n472), .C1(new_n482), .C2(new_n483), .ZN(new_n923));
  OAI21_X1  g498(.A(G8), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(G305), .A2(G1981), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT108), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT107), .ZN(new_n928));
  OR2_X1    g503(.A1(new_n928), .A2(G1981), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(G1981), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n927), .B1(new_n738), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n931), .ZN(new_n933));
  NOR4_X1   g508(.A1(new_n733), .A2(new_n737), .A3(KEYINPUT108), .A4(new_n933), .ZN(new_n934));
  OAI211_X1 g509(.A(KEYINPUT49), .B(new_n926), .C1(new_n932), .C2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(KEYINPUT109), .ZN(new_n936));
  OAI21_X1  g511(.A(KEYINPUT108), .B1(G305), .B2(new_n933), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n738), .A2(new_n927), .A3(new_n931), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT109), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n939), .A2(new_n940), .A3(KEYINPUT49), .A4(new_n926), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n936), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n939), .A2(new_n926), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT49), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n924), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  AOI211_X1 g520(.A(G1976), .B(G288), .C1(new_n942), .C2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n939), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n925), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT52), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n949), .B1(new_n597), .B2(G1976), .ZN(new_n950));
  INV_X1    g525(.A(G1976), .ZN(new_n951));
  OAI211_X1 g526(.A(new_n950), .B(new_n925), .C1(new_n951), .C2(G288), .ZN(new_n952));
  AOI211_X1 g527(.A(new_n951), .B(new_n593), .C1(new_n595), .C2(new_n596), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n949), .B1(new_n953), .B2(new_n924), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n956), .B1(new_n942), .B2(new_n945), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(G8), .ZN(new_n959));
  XNOR2_X1  g534(.A(KEYINPUT103), .B(KEYINPUT45), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n852), .A2(new_n921), .A3(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT112), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n852), .A2(KEYINPUT112), .A3(new_n921), .A4(new_n961), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n923), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT45), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n968), .B1(G164), .B2(G1384), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n967), .A2(KEYINPUT111), .A3(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT111), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT45), .B1(new_n852), .B2(new_n921), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n971), .B1(new_n972), .B2(new_n923), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n966), .A2(new_n970), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(new_n824), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT50), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n852), .A2(new_n976), .A3(new_n921), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT105), .ZN(new_n978));
  OAI21_X1  g553(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n977), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n922), .A2(KEYINPUT105), .A3(KEYINPUT50), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n923), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n775), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n959), .B1(new_n975), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(G303), .A2(G8), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT55), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n980), .A2(new_n981), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n967), .A2(new_n803), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n960), .B1(G164), .B2(G1384), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n852), .A2(KEYINPUT45), .A3(new_n921), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n967), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  XOR2_X1   g571(.A(KEYINPUT104), .B(G1971), .Z(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n959), .B1(new_n993), .B2(new_n999), .ZN(new_n1000));
  OAI211_X1 g575(.A(new_n984), .B(G168), .C1(new_n989), .C2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(KEYINPUT63), .B1(new_n958), .B2(new_n1001), .ZN(new_n1002));
  NOR3_X1   g577(.A1(new_n972), .A2(new_n971), .A3(new_n923), .ZN(new_n1003));
  AOI21_X1  g578(.A(KEYINPUT111), .B1(new_n967), .B2(new_n969), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(G1966), .B1(new_n1005), .B2(new_n966), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n982), .A2(new_n775), .ZN(new_n1007));
  OAI21_X1  g582(.A(G8), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1008), .A2(G286), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT110), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n967), .A2(new_n977), .A3(new_n803), .A4(new_n979), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n959), .B1(new_n999), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1010), .B1(new_n1012), .B2(new_n989), .ZN(new_n1013));
  AND2_X1   g588(.A1(new_n987), .A2(new_n988), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n976), .B1(new_n852), .B2(new_n921), .ZN(new_n1015));
  NOR3_X1   g590(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1016));
  NOR3_X1   g591(.A1(new_n1015), .A2(new_n1016), .A3(new_n923), .ZN(new_n1017));
  AOI22_X1  g592(.A1(new_n1017), .A2(new_n803), .B1(new_n996), .B2(new_n998), .ZN(new_n1018));
  OAI211_X1 g593(.A(KEYINPUT110), .B(new_n1014), .C1(new_n1018), .C2(new_n959), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT63), .B1(new_n1013), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n991), .B1(new_n981), .B2(new_n980), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n923), .B1(new_n922), .B2(new_n960), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n997), .B1(new_n1022), .B2(new_n995), .ZN(new_n1023));
  OAI211_X1 g598(.A(G8), .B(new_n989), .C1(new_n1021), .C2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT106), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n993), .A2(new_n999), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1027), .A2(KEYINPUT106), .A3(G8), .A4(new_n989), .ZN(new_n1028));
  AOI22_X1  g603(.A1(new_n1009), .A2(new_n1020), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n948), .B(new_n1002), .C1(new_n958), .C2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n967), .A2(new_n979), .A3(new_n977), .ZN(new_n1031));
  INV_X1    g606(.A(G1956), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g608(.A(KEYINPUT56), .B(G2072), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n967), .A2(new_n995), .A3(new_n994), .A4(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1036));
  AOI21_X1  g611(.A(KEYINPUT57), .B1(new_n584), .B2(new_n586), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n579), .A2(new_n1037), .ZN(new_n1038));
  AOI22_X1  g613(.A1(new_n1033), .A2(new_n1035), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n990), .A2(new_n967), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(KEYINPUT114), .ZN(new_n1042));
  INV_X1    g617(.A(G1348), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT114), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n982), .A2(new_n1044), .ZN(new_n1045));
  AND3_X1   g620(.A1(new_n1042), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n922), .A2(new_n923), .ZN(new_n1047));
  INV_X1    g622(.A(G2067), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g624(.A(new_n1049), .B(KEYINPUT113), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1046), .A2(new_n1051), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1033), .A2(new_n1036), .A3(new_n1038), .A4(new_n1035), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(new_n626), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1040), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  XOR2_X1   g630(.A(KEYINPUT115), .B(KEYINPUT61), .Z(new_n1056));
  INV_X1    g631(.A(KEYINPUT116), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1039), .B1(new_n1057), .B2(new_n1053), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1060));
  AND3_X1   g635(.A1(new_n1059), .A2(new_n1057), .A3(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1056), .B1(new_n1058), .B2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1042), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1063), .A2(KEYINPUT60), .A3(new_n625), .A4(new_n1050), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT61), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1039), .A2(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g641(.A(KEYINPUT58), .B(G1341), .ZN(new_n1067));
  OAI22_X1  g642(.A1(new_n996), .A2(G1996), .B1(new_n1047), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(new_n566), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(KEYINPUT59), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT59), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1068), .A2(new_n1071), .A3(new_n566), .ZN(new_n1072));
  AOI22_X1  g647(.A1(new_n1066), .A2(new_n1053), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1073));
  AND3_X1   g648(.A1(new_n1062), .A2(new_n1064), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT60), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1075), .B1(new_n1046), .B2(new_n1051), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1063), .A2(KEYINPUT60), .A3(new_n1050), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1076), .A2(new_n626), .A3(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1055), .B1(new_n1074), .B2(new_n1078), .ZN(new_n1079));
  AOI22_X1  g654(.A1(new_n1028), .A2(new_n1026), .B1(new_n1013), .B2(new_n1019), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(new_n957), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(KEYINPUT121), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT121), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1080), .A2(new_n957), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1079), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT118), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n551), .A2(G8), .A3(new_n552), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT117), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT51), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1088), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n551), .A2(KEYINPUT117), .A3(G8), .A4(new_n552), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  AOI22_X1  g668(.A1(new_n974), .A2(new_n824), .B1(new_n982), .B2(new_n775), .ZN(new_n1094));
  OAI22_X1  g669(.A1(new_n984), .A2(new_n1093), .B1(new_n1088), .B2(new_n1094), .ZN(new_n1095));
  AOI211_X1 g670(.A(KEYINPUT51), .B(new_n959), .C1(new_n1094), .C2(G168), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1087), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1093), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1008), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n975), .A2(new_n983), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1090), .B(G8), .C1(new_n1100), .C2(G286), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1088), .B1(new_n975), .B2(new_n983), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1099), .A2(new_n1101), .A3(KEYINPUT118), .A4(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1097), .A2(new_n1104), .ZN(new_n1105));
  XOR2_X1   g680(.A(KEYINPUT119), .B(KEYINPUT54), .Z(new_n1106));
  INV_X1    g681(.A(new_n996), .ZN(new_n1107));
  INV_X1    g682(.A(G2078), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  XNOR2_X1  g684(.A(KEYINPUT120), .B(KEYINPUT53), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n982), .B(KEYINPUT114), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1112), .B1(new_n1113), .B2(new_n789), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1005), .A2(KEYINPUT53), .A3(new_n1108), .A4(new_n966), .ZN(new_n1115));
  AOI21_X1  g690(.A(G301), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1042), .A2(new_n789), .A3(new_n1045), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1107), .A2(KEYINPUT53), .A3(new_n1108), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1117), .A2(new_n1111), .A3(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1119), .A2(G171), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1106), .B1(new_n1116), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1119), .A2(G171), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1123));
  OAI211_X1 g698(.A(KEYINPUT54), .B(new_n1122), .C1(new_n1123), .C2(G171), .ZN(new_n1124));
  AND3_X1   g699(.A1(new_n1105), .A2(new_n1121), .A3(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1030), .B1(new_n1086), .B2(new_n1125), .ZN(new_n1126));
  AND3_X1   g701(.A1(new_n1080), .A2(new_n957), .A3(new_n1083), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1083), .B1(new_n1080), .B2(new_n957), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1123), .A2(G171), .ZN(new_n1129));
  NOR3_X1   g704(.A1(new_n1127), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  NOR3_X1   g705(.A1(new_n1095), .A2(new_n1096), .A3(new_n1087), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1102), .B1(new_n1008), .B2(new_n1098), .ZN(new_n1132));
  AOI21_X1  g707(.A(KEYINPUT118), .B1(new_n1132), .B2(new_n1101), .ZN(new_n1133));
  OAI21_X1  g708(.A(KEYINPUT62), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT62), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1097), .A2(new_n1135), .A3(new_n1104), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1130), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(KEYINPUT122), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT122), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1130), .A2(new_n1134), .A3(new_n1139), .A4(new_n1136), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1126), .A2(new_n1138), .A3(new_n1140), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n994), .A2(new_n923), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n709), .A2(new_n711), .ZN(new_n1143));
  XNOR2_X1  g718(.A(new_n755), .B(G1996), .ZN(new_n1144));
  XNOR2_X1  g719(.A(new_n785), .B(new_n1048), .ZN(new_n1145));
  AND2_X1   g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  OR2_X1    g721(.A1(new_n717), .A2(new_n720), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n717), .A2(new_n720), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1143), .A2(new_n1146), .A3(new_n1147), .A4(new_n1148), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n709), .A2(new_n711), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1142), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1141), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1142), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1153), .B1(new_n1145), .B2(new_n755), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1154), .B(KEYINPUT124), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1142), .A2(new_n758), .ZN(new_n1156));
  XNOR2_X1  g731(.A(new_n1156), .B(KEYINPUT46), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  XNOR2_X1  g733(.A(new_n1158), .B(KEYINPUT47), .ZN(new_n1159));
  XOR2_X1   g734(.A(new_n1147), .B(KEYINPUT123), .Z(new_n1160));
  AOI22_X1  g735(.A1(new_n1146), .A2(new_n1160), .B1(new_n1048), .B2(new_n786), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1143), .A2(new_n1153), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1162), .B(KEYINPUT48), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1146), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(new_n1142), .ZN(new_n1165));
  XNOR2_X1  g740(.A(new_n1165), .B(KEYINPUT125), .ZN(new_n1166));
  OAI221_X1 g741(.A(new_n1159), .B1(new_n1153), .B2(new_n1161), .C1(new_n1163), .C2(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1167), .B(KEYINPUT126), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1152), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT127), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1152), .A2(KEYINPUT127), .A3(new_n1168), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1171), .A2(new_n1172), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g748(.A1(G401), .A2(G229), .A3(new_n460), .A4(G227), .ZN(new_n1175));
  NAND3_X1  g749(.A1(new_n913), .A2(new_n867), .A3(new_n1175), .ZN(G225));
  INV_X1    g750(.A(G225), .ZN(G308));
endmodule


