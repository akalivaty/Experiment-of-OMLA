//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 1 1 1 1 0 1 0 0 0 0 0 0 0 0 0 1 1 1 1 1 0 1 1 0 1 0 1 0 0 0 0 0 1 0 0 1 1 1 1 1 0 0 0 0 1 1 1 0 1 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:46 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G87), .ZN(new_n207));
  INV_X1    g0007(.A(G250), .ZN(new_n208));
  INV_X1    g0008(.A(G97), .ZN(new_n209));
  INV_X1    g0009(.A(G257), .ZN(new_n210));
  OAI22_X1  g0010(.A1(new_n207), .A2(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI21_X1  g0011(.A(new_n211), .B1(G68), .B2(G238), .ZN(new_n212));
  INV_X1    g0012(.A(G107), .ZN(new_n213));
  INV_X1    g0013(.A(G264), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AOI21_X1  g0015(.A(new_n215), .B1(G116), .B2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G50), .ZN(new_n217));
  INV_X1    g0017(.A(G226), .ZN(new_n218));
  INV_X1    g0018(.A(G77), .ZN(new_n219));
  INV_X1    g0019(.A(G244), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G58), .ZN(new_n222));
  INV_X1    g0022(.A(G232), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n206), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT1), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n204), .A2(KEYINPUT64), .ZN(new_n227));
  INV_X1    g0027(.A(KEYINPUT64), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G20), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  OAI21_X1  g0031(.A(G50), .B1(G58), .B2(G68), .ZN(new_n232));
  NOR3_X1   g0032(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n206), .A2(G13), .ZN(new_n234));
  OAI211_X1 g0034(.A(new_n234), .B(G250), .C1(G257), .C2(G264), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n235), .B(KEYINPUT0), .Z(new_n236));
  NOR3_X1   g0036(.A1(new_n226), .A2(new_n233), .A3(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(new_n214), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(G270), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G68), .B(G77), .Z(new_n246));
  XOR2_X1   g0046(.A(G50), .B(G58), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G97), .B(G107), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  AND2_X1   g0053(.A1(new_n253), .A2(new_n231), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  AND2_X1   g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT7), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n230), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  OR2_X1    g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n261), .A2(new_n204), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(KEYINPUT7), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n260), .A2(new_n264), .A3(G68), .ZN(new_n265));
  XNOR2_X1  g0065(.A(G58), .B(G68), .ZN(new_n266));
  NOR2_X1   g0066(.A1(G20), .A2(G33), .ZN(new_n267));
  AOI22_X1  g0067(.A1(new_n266), .A2(G20), .B1(G159), .B2(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n265), .A2(KEYINPUT16), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n268), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n230), .A2(new_n258), .A3(KEYINPUT7), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n263), .A2(new_n259), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n270), .B1(new_n273), .B2(G68), .ZN(new_n274));
  OAI211_X1 g0074(.A(new_n255), .B(new_n269), .C1(new_n274), .C2(KEYINPUT16), .ZN(new_n275));
  XOR2_X1   g0075(.A(KEYINPUT8), .B(G58), .Z(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n255), .B1(new_n203), .B2(G20), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n280), .B1(new_n282), .B2(new_n277), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G33), .ZN(new_n285));
  INV_X1    g0085(.A(G41), .ZN(new_n286));
  OAI211_X1 g0086(.A(G1), .B(G13), .C1(new_n285), .C2(new_n286), .ZN(new_n287));
  OR2_X1    g0087(.A1(G223), .A2(G1698), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n218), .A2(G1698), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n288), .B(new_n289), .C1(new_n256), .C2(new_n257), .ZN(new_n290));
  NAND2_X1  g0090(.A1(G33), .A2(G87), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n287), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n287), .A2(G232), .A3(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n293), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G274), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(G200), .B1(new_n292), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n297), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n290), .A2(new_n291), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n231), .B1(G33), .B2(G41), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n299), .A2(new_n302), .A3(G190), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n275), .A2(new_n284), .A3(new_n298), .A4(new_n303), .ZN(new_n304));
  XNOR2_X1  g0104(.A(new_n304), .B(KEYINPUT17), .ZN(new_n305));
  INV_X1    g0105(.A(G179), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n299), .A2(new_n302), .A3(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G169), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n308), .B1(new_n292), .B2(new_n297), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n307), .A2(KEYINPUT73), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT73), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n299), .A2(new_n302), .A3(new_n311), .A4(new_n306), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(KEYINPUT74), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT74), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n310), .A2(new_n315), .A3(new_n312), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n275), .A2(new_n284), .ZN(new_n318));
  AOI21_X1  g0118(.A(KEYINPUT18), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  AND3_X1   g0119(.A1(new_n310), .A2(new_n315), .A3(new_n312), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n315), .B1(new_n310), .B2(new_n312), .ZN(new_n321));
  OAI211_X1 g0121(.A(KEYINPUT18), .B(new_n318), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n305), .B1(new_n319), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n296), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n261), .A2(new_n262), .ZN(new_n326));
  NAND2_X1  g0126(.A1(G238), .A2(G1698), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n326), .B(new_n327), .C1(new_n223), .C2(G1698), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n287), .B1(new_n258), .B2(new_n213), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n325), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n301), .A2(new_n295), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G244), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(G190), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n335), .B1(G200), .B2(new_n333), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT65), .ZN(new_n338));
  XNOR2_X1  g0138(.A(KEYINPUT64), .B(G20), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n338), .B1(new_n339), .B2(new_n285), .ZN(new_n340));
  XOR2_X1   g0140(.A(KEYINPUT15), .B(G87), .Z(new_n341));
  NOR2_X1   g0141(.A1(new_n228), .A2(G20), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n204), .A2(KEYINPUT64), .ZN(new_n343));
  OAI211_X1 g0143(.A(KEYINPUT65), .B(G33), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n340), .A2(new_n341), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n339), .A2(G77), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n276), .A2(new_n267), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n255), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n281), .A2(G77), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n279), .A2(new_n219), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  OR2_X1    g0152(.A1(new_n337), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n333), .A2(new_n308), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(KEYINPUT67), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n330), .A2(new_n306), .A3(new_n332), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT67), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n352), .A2(new_n358), .A3(new_n354), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n356), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n353), .A2(new_n360), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n324), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(G68), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n279), .A2(KEYINPUT70), .A3(KEYINPUT12), .A4(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n279), .A2(new_n363), .ZN(new_n365));
  XOR2_X1   g0165(.A(KEYINPUT70), .B(KEYINPUT12), .Z(new_n366));
  AOI22_X1  g0166(.A1(new_n281), .A2(G68), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT11), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n340), .A2(G77), .A3(new_n344), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n267), .A2(G50), .B1(G20), .B2(new_n363), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n368), .B1(new_n371), .B2(new_n255), .ZN(new_n372));
  AOI211_X1 g0172(.A(KEYINPUT11), .B(new_n254), .C1(new_n369), .C2(new_n370), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n364), .B(new_n367), .C1(new_n372), .C2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(G1698), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n218), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n223), .A2(G1698), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n377), .B(new_n378), .C1(new_n256), .C2(new_n257), .ZN(new_n379));
  NAND2_X1  g0179(.A1(G33), .A2(G97), .ZN(new_n380));
  AND3_X1   g0180(.A1(new_n379), .A2(KEYINPUT69), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT69), .B1(new_n379), .B2(new_n380), .ZN(new_n382));
  NOR3_X1   g0182(.A1(new_n381), .A2(new_n382), .A3(new_n287), .ZN(new_n383));
  INV_X1    g0183(.A(new_n331), .ZN(new_n384));
  INV_X1    g0184(.A(G238), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n296), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(KEYINPUT13), .B1(new_n383), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n382), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n379), .A2(KEYINPUT69), .A3(new_n380), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(new_n301), .A3(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT13), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n325), .B1(new_n331), .B2(G238), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n387), .A2(new_n393), .A3(G179), .ZN(new_n394));
  XNOR2_X1  g0194(.A(new_n394), .B(KEYINPUT71), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT14), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n387), .A2(new_n393), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n396), .B1(new_n397), .B2(G169), .ZN(new_n398));
  AOI211_X1 g0198(.A(KEYINPUT14), .B(new_n308), .C1(new_n387), .C2(new_n393), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n375), .B1(new_n395), .B2(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n397), .A2(new_n334), .ZN(new_n402));
  INV_X1    g0202(.A(G200), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n403), .B1(new_n387), .B2(new_n393), .ZN(new_n404));
  NOR3_X1   g0204(.A1(new_n402), .A2(new_n374), .A3(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(KEYINPUT72), .B1(new_n401), .B2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT68), .ZN(new_n407));
  AND2_X1   g0207(.A1(new_n407), .A2(KEYINPUT10), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n376), .A2(G222), .ZN(new_n409));
  NAND2_X1  g0209(.A1(G223), .A2(G1698), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n326), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n411), .B(new_n301), .C1(G77), .C2(new_n326), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n331), .A2(G226), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n412), .A2(new_n296), .A3(new_n413), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n414), .A2(new_n334), .ZN(new_n415));
  AOI211_X1 g0215(.A(new_n408), .B(new_n415), .C1(G200), .C2(new_n414), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n282), .A2(new_n217), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n340), .A2(new_n344), .A3(new_n276), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n217), .A2(new_n222), .A3(new_n363), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n420), .A2(G20), .B1(G150), .B2(new_n267), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n422), .A2(new_n255), .B1(new_n217), .B2(new_n279), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n418), .A2(new_n423), .ZN(new_n424));
  AND2_X1   g0224(.A1(new_n424), .A2(KEYINPUT9), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n424), .A2(KEYINPUT9), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n416), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n407), .A2(KEYINPUT10), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  OAI221_X1 g0229(.A(new_n416), .B1(new_n407), .B2(KEYINPUT10), .C1(new_n425), .C2(new_n426), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n414), .A2(G179), .ZN(new_n431));
  XNOR2_X1  g0231(.A(new_n431), .B(KEYINPUT66), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n414), .A2(new_n308), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n432), .A2(new_n424), .A3(new_n433), .ZN(new_n434));
  AND3_X1   g0234(.A1(new_n429), .A2(new_n430), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n397), .A2(G169), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT14), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n397), .A2(new_n396), .A3(G169), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT71), .ZN(new_n440));
  XNOR2_X1  g0240(.A(new_n394), .B(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n374), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT72), .ZN(new_n443));
  INV_X1    g0243(.A(new_n405), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  AND4_X1   g0245(.A1(new_n362), .A2(new_n406), .A3(new_n435), .A4(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n203), .A2(G33), .ZN(new_n448));
  AND3_X1   g0248(.A1(new_n254), .A2(new_n448), .A3(new_n278), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(G107), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT23), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n227), .A2(new_n229), .A3(new_n452), .A4(new_n213), .ZN(new_n453));
  NAND2_X1  g0253(.A1(G33), .A2(G116), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(new_n452), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n204), .ZN(new_n456));
  NAND2_X1  g0256(.A1(KEYINPUT23), .A2(G107), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n453), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT22), .ZN(new_n460));
  AOI22_X1  g0260(.A1(new_n227), .A2(new_n229), .B1(new_n261), .B2(new_n262), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n460), .B1(new_n461), .B2(G87), .ZN(new_n462));
  AND4_X1   g0262(.A1(new_n460), .A2(new_n326), .A3(new_n230), .A4(G87), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n459), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT24), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n326), .A2(new_n230), .A3(G87), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(KEYINPUT22), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n326), .A2(new_n230), .A3(new_n460), .A4(G87), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT24), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n469), .A2(new_n470), .A3(new_n459), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n465), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n451), .B1(new_n472), .B2(new_n255), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n278), .A2(G107), .ZN(new_n474));
  XNOR2_X1  g0274(.A(new_n474), .B(KEYINPUT25), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT78), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n286), .A2(KEYINPUT5), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n203), .A2(G45), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT5), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(G41), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n481), .A2(KEYINPUT78), .A3(new_n203), .A4(G45), .ZN(new_n482));
  AND2_X1   g0282(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n286), .A2(KEYINPUT5), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n483), .A2(G274), .A3(new_n287), .A4(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n208), .A2(new_n376), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n210), .A2(G1698), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n486), .B(new_n487), .C1(new_n256), .C2(new_n257), .ZN(new_n488));
  INV_X1    g0288(.A(G294), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n488), .B1(new_n285), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n301), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n479), .A2(new_n484), .A3(new_n482), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n492), .A2(G264), .A3(new_n287), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n485), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G200), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n493), .A2(new_n491), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n479), .A2(new_n482), .A3(G274), .A4(new_n484), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n497), .A2(new_n301), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(G190), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n473), .A2(new_n475), .A3(new_n495), .A4(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(G169), .B1(new_n496), .B2(new_n498), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(KEYINPUT85), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n499), .A2(G179), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT85), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n494), .A2(new_n505), .A3(G169), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n503), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n470), .B1(new_n469), .B2(new_n459), .ZN(new_n508));
  AOI211_X1 g0308(.A(KEYINPUT24), .B(new_n458), .C1(new_n467), .C2(new_n468), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n255), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n510), .A2(new_n450), .A3(new_n475), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n501), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n492), .A2(G270), .A3(new_n287), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n376), .A2(G257), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n326), .B(new_n515), .C1(new_n214), .C2(new_n376), .ZN(new_n516));
  INV_X1    g0316(.A(G303), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n258), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n516), .A2(new_n301), .A3(new_n518), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n514), .B(new_n519), .C1(new_n301), .C2(new_n497), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n520), .A2(KEYINPUT21), .A3(G169), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n485), .A2(G179), .A3(new_n519), .A4(new_n514), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n449), .A2(G116), .ZN(new_n524));
  INV_X1    g0324(.A(G116), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n279), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(G33), .A2(G283), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n285), .A2(G97), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n527), .B(new_n528), .C1(new_n342), .C2(new_n343), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n253), .A2(new_n231), .B1(G20), .B2(new_n525), .ZN(new_n530));
  AND3_X1   g0330(.A1(new_n529), .A2(KEYINPUT20), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(KEYINPUT20), .B1(new_n529), .B2(new_n530), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n524), .B(new_n526), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n523), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n520), .A2(G200), .ZN(new_n535));
  INV_X1    g0335(.A(new_n533), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n535), .B(new_n536), .C1(new_n334), .C2(new_n520), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n520), .A2(new_n533), .A3(G169), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT21), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n538), .A2(KEYINPUT84), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(KEYINPUT84), .B1(new_n538), .B2(new_n539), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n534), .B(new_n537), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n513), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n340), .A2(G97), .A3(new_n344), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT19), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n230), .B1(new_n545), .B2(new_n380), .ZN(new_n547));
  XNOR2_X1  g0347(.A(KEYINPUT82), .B(G87), .ZN(new_n548));
  NOR2_X1   g0348(.A1(G97), .A2(G107), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n547), .A2(new_n550), .B1(new_n461), .B2(G68), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n546), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(KEYINPUT83), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT83), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n546), .A2(new_n554), .A3(new_n551), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n553), .A2(new_n255), .A3(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(new_n341), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n279), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n449), .A2(G87), .ZN(new_n559));
  AND3_X1   g0359(.A1(new_n556), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n385), .A2(new_n376), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n326), .B(new_n561), .C1(G244), .C2(new_n376), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n287), .B1(new_n562), .B2(new_n454), .ZN(new_n563));
  INV_X1    g0363(.A(G274), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n478), .A2(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n287), .A2(G250), .A3(new_n478), .ZN(new_n567));
  XOR2_X1   g0367(.A(new_n567), .B(KEYINPUT81), .Z(new_n568));
  NAND2_X1  g0368(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n403), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n566), .A2(new_n568), .A3(new_n334), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n449), .A2(new_n341), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n556), .A2(new_n573), .A3(new_n558), .ZN(new_n574));
  XNOR2_X1  g0374(.A(new_n567), .B(KEYINPUT81), .ZN(new_n575));
  NOR4_X1   g0375(.A1(new_n575), .A2(new_n563), .A3(G179), .A4(new_n565), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n576), .B1(new_n308), .B2(new_n569), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n560), .A2(new_n572), .B1(new_n574), .B2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT6), .ZN(new_n579));
  NOR3_X1   g0379(.A1(new_n579), .A2(new_n209), .A3(G107), .ZN(new_n580));
  XNOR2_X1  g0380(.A(G97), .B(G107), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n580), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(new_n267), .ZN(new_n583));
  OAI22_X1  g0383(.A1(new_n582), .A2(new_n230), .B1(new_n219), .B2(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n213), .B1(new_n271), .B2(new_n272), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n255), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n449), .A2(G97), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n278), .A2(G97), .ZN(new_n588));
  XNOR2_X1  g0388(.A(new_n588), .B(KEYINPUT75), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n586), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT76), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n586), .A2(KEYINPUT76), .A3(new_n587), .A4(new_n589), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT79), .ZN(new_n595));
  AND3_X1   g0395(.A1(new_n492), .A2(G257), .A3(new_n287), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n596), .A2(new_n498), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT4), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n598), .A2(G1698), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n599), .B(G244), .C1(new_n257), .C2(new_n256), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n220), .B1(new_n261), .B2(new_n262), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n600), .B(new_n527), .C1(new_n601), .C2(KEYINPUT4), .ZN(new_n602));
  OAI21_X1  g0402(.A(G250), .B1(new_n256), .B2(new_n257), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n376), .B1(new_n603), .B2(KEYINPUT4), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n301), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n595), .B1(new_n597), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n492), .A2(G257), .A3(new_n287), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n605), .A2(new_n485), .A3(new_n595), .A4(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(G190), .B1(new_n606), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n605), .A2(KEYINPUT77), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT77), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n612), .B(new_n301), .C1(new_n602), .C2(new_n604), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n611), .A2(new_n597), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(G200), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n594), .A2(new_n610), .A3(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT80), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n605), .A2(new_n607), .A3(new_n485), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(KEYINPUT79), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n619), .A2(new_n308), .A3(new_n608), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n611), .A2(new_n597), .A3(new_n306), .A4(new_n613), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n620), .A2(new_n621), .A3(new_n590), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n616), .A2(new_n617), .A3(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n617), .B1(new_n616), .B2(new_n622), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n543), .B(new_n578), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n447), .A2(new_n625), .ZN(G372));
  INV_X1    g0426(.A(new_n434), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT86), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n360), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n356), .A2(KEYINPUT86), .A3(new_n357), .A4(new_n359), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n442), .B1(new_n631), .B2(new_n405), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n305), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n633), .B1(new_n319), .B2(new_n323), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n429), .A2(new_n430), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n627), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n616), .A2(new_n622), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n572), .A2(new_n556), .A3(new_n558), .A4(new_n559), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n538), .A2(new_n539), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT84), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n538), .A2(KEYINPUT84), .A3(new_n539), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n644), .A2(new_n512), .A3(new_n534), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n638), .A2(new_n639), .A3(new_n501), .A4(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n574), .A2(new_n577), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT26), .ZN(new_n648));
  AND4_X1   g0448(.A1(new_n620), .A2(new_n621), .A3(new_n592), .A4(new_n593), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n578), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n620), .A2(new_n621), .A3(new_n590), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n651), .A2(new_n647), .A3(new_n639), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(KEYINPUT26), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n646), .A2(new_n647), .A3(new_n650), .A4(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n446), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n637), .A2(new_n655), .ZN(G369));
  XOR2_X1   g0456(.A(new_n542), .B(KEYINPUT88), .Z(new_n657));
  INV_X1    g0457(.A(G13), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n339), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(new_n203), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n660), .A2(KEYINPUT27), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(KEYINPUT27), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n661), .A2(G213), .A3(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(G343), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n533), .ZN(new_n666));
  XNOR2_X1  g0466(.A(new_n666), .B(KEYINPUT87), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n657), .A2(new_n667), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n644), .A2(new_n534), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n668), .B1(new_n669), .B2(new_n667), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(G330), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  AND3_X1   g0472(.A1(new_n511), .A2(KEYINPUT89), .A3(new_n665), .ZN(new_n673));
  AOI21_X1  g0473(.A(KEYINPUT89), .B1(new_n511), .B2(new_n665), .ZN(new_n674));
  OR3_X1    g0474(.A1(new_n513), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n665), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n675), .B1(new_n512), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n672), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n507), .A2(new_n511), .A3(new_n676), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n669), .A2(new_n665), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(new_n675), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n678), .A2(new_n679), .A3(new_n683), .ZN(G399));
  INV_X1    g0484(.A(new_n234), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(G41), .ZN(new_n686));
  INV_X1    g0486(.A(new_n550), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n525), .ZN(new_n688));
  NOR3_X1   g0488(.A1(new_n686), .A2(new_n203), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n232), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n689), .B1(new_n690), .B2(new_n686), .ZN(new_n691));
  XOR2_X1   g0491(.A(new_n691), .B(KEYINPUT28), .Z(new_n692));
  NAND2_X1  g0492(.A1(new_n652), .A2(new_n648), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT92), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n652), .A2(KEYINPUT92), .A3(new_n648), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n649), .A2(KEYINPUT26), .A3(new_n647), .A4(new_n639), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(KEYINPUT91), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT91), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n578), .A2(new_n699), .A3(KEYINPUT26), .A4(new_n649), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n695), .A2(new_n696), .A3(new_n698), .A4(new_n700), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n646), .A2(new_n647), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n703), .A2(KEYINPUT29), .A3(new_n676), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n654), .A2(new_n676), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT29), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n569), .A2(new_n496), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT90), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n522), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n619), .A2(new_n608), .ZN(new_n712));
  OAI21_X1  g0512(.A(KEYINPUT90), .B1(new_n569), .B2(new_n496), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT30), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n711), .A2(KEYINPUT30), .A3(new_n712), .A4(new_n713), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n614), .A2(new_n306), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n718), .A2(new_n569), .A3(new_n494), .A4(new_n520), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n716), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(new_n665), .ZN(new_n721));
  OAI211_X1 g0521(.A(KEYINPUT31), .B(new_n721), .C1(new_n625), .C2(new_n665), .ZN(new_n722));
  OR2_X1    g0522(.A1(new_n721), .A2(KEYINPUT31), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(G330), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n708), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n692), .B1(new_n727), .B2(G1), .ZN(G364));
  AOI21_X1  g0528(.A(new_n231), .B1(G20), .B2(new_n308), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(G179), .A2(G190), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n339), .A2(G200), .A3(new_n731), .ZN(new_n732));
  OR2_X1    g0532(.A1(new_n732), .A2(KEYINPUT97), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(KEYINPUT97), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(new_n213), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n230), .A2(new_n306), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(new_n334), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(G200), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n339), .A2(new_n403), .A3(new_n731), .ZN(new_n741));
  INV_X1    g0541(.A(G159), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  OAI22_X1  g0544(.A1(new_n740), .A2(new_n219), .B1(KEYINPUT32), .B2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n334), .A2(G200), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n737), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  AOI211_X1 g0548(.A(new_n736), .B(new_n745), .C1(G58), .C2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n746), .A2(new_n306), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(new_n339), .ZN(new_n751));
  AOI22_X1  g0551(.A1(new_n744), .A2(KEYINPUT32), .B1(G97), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n334), .A2(new_n403), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n753), .A2(G20), .A3(new_n306), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n738), .A2(new_n403), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  OAI221_X1 g0556(.A(new_n752), .B1(new_n548), .B2(new_n754), .C1(new_n363), .C2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(new_n258), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n737), .A2(new_n753), .ZN(new_n759));
  OAI211_X1 g0559(.A(new_n749), .B(new_n758), .C1(new_n217), .C2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n751), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n489), .ZN(new_n762));
  INV_X1    g0562(.A(G311), .ZN(new_n763));
  OAI22_X1  g0563(.A1(new_n740), .A2(new_n763), .B1(new_n517), .B2(new_n754), .ZN(new_n764));
  INV_X1    g0564(.A(new_n735), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n762), .B(new_n764), .C1(G283), .C2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n759), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G326), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n748), .A2(G322), .ZN(new_n769));
  XOR2_X1   g0569(.A(KEYINPUT33), .B(G317), .Z(new_n770));
  NOR2_X1   g0570(.A1(new_n756), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n741), .ZN(new_n772));
  AOI211_X1 g0572(.A(new_n326), .B(new_n771), .C1(G329), .C2(new_n772), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n766), .A2(new_n768), .A3(new_n769), .A4(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n730), .B1(new_n760), .B2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(G45), .ZN(new_n776));
  NOR3_X1   g0576(.A1(new_n339), .A2(new_n658), .A3(new_n776), .ZN(new_n777));
  OR2_X1    g0577(.A1(new_n777), .A2(KEYINPUT95), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(KEYINPUT95), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n778), .A2(G1), .A3(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n686), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(G13), .A2(G33), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(G20), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n729), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(KEYINPUT96), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n685), .A2(new_n326), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n789), .B1(new_n776), .B2(new_n690), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n248), .A2(G45), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n790), .A2(new_n791), .B1(new_n525), .B2(new_n685), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n234), .A2(G355), .A3(new_n326), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n787), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NOR3_X1   g0594(.A1(new_n775), .A2(new_n782), .A3(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n785), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n795), .B1(new_n670), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n670), .A2(G330), .ZN(new_n798));
  OR2_X1    g0598(.A1(new_n798), .A2(KEYINPUT93), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n798), .A2(KEYINPUT93), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n799), .A2(new_n782), .A3(new_n800), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n671), .B(KEYINPUT94), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n797), .B1(new_n801), .B2(new_n802), .ZN(G396));
  INV_X1    g0603(.A(new_n361), .ZN(new_n804));
  NAND4_X1  g0604(.A1(new_n645), .A2(new_n622), .A3(new_n616), .A4(new_n501), .ZN(new_n805));
  INV_X1    g0605(.A(new_n639), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n647), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n650), .A2(new_n653), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n804), .B(new_n676), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(KEYINPUT98), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND4_X1  g0611(.A1(new_n654), .A2(KEYINPUT98), .A3(new_n804), .A4(new_n676), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n352), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n361), .B1(new_n814), .B2(new_n676), .ZN(new_n815));
  NAND4_X1  g0615(.A1(new_n629), .A2(new_n352), .A3(new_n630), .A4(new_n665), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n705), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n813), .A2(new_n818), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(new_n726), .Z(new_n820));
  NOR2_X1   g0620(.A1(new_n820), .A2(new_n781), .ZN(new_n821));
  INV_X1    g0621(.A(new_n817), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n822), .A2(new_n784), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n729), .A2(new_n783), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n825), .A2(G77), .ZN(new_n826));
  INV_X1    g0626(.A(new_n754), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(G50), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n755), .A2(G150), .B1(new_n748), .B2(G143), .ZN(new_n829));
  INV_X1    g0629(.A(G137), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n829), .B1(new_n830), .B2(new_n759), .C1(new_n742), .C2(new_n740), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT34), .ZN(new_n832));
  OR2_X1    g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n831), .A2(new_n832), .B1(G68), .B2(new_n765), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n258), .B1(new_n772), .B2(G132), .ZN(new_n835));
  AND4_X1   g0635(.A1(new_n828), .A2(new_n833), .A3(new_n834), .A4(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(new_n222), .B2(new_n761), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n735), .A2(new_n207), .B1(new_n213), .B2(new_n754), .ZN(new_n838));
  INV_X1    g0638(.A(G283), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n756), .A2(new_n839), .B1(new_n209), .B2(new_n761), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n740), .A2(new_n525), .B1(new_n759), .B2(new_n517), .ZN(new_n841));
  NOR4_X1   g0641(.A1(new_n838), .A2(new_n326), .A3(new_n840), .A4(new_n841), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n842), .B1(new_n489), .B2(new_n747), .C1(new_n763), .C2(new_n741), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n730), .B1(new_n837), .B2(new_n843), .ZN(new_n844));
  NOR4_X1   g0644(.A1(new_n823), .A2(new_n782), .A3(new_n826), .A4(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n821), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(G384));
  INV_X1    g0647(.A(new_n663), .ZN(new_n848));
  OR3_X1    g0648(.A1(new_n319), .A2(new_n323), .A3(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n360), .A2(new_n665), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n851), .B1(new_n811), .B2(new_n812), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n374), .A2(new_n665), .ZN(new_n853));
  OR2_X1    g0653(.A1(new_n853), .A2(KEYINPUT99), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(KEYINPUT99), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n442), .A2(new_n854), .A3(new_n444), .A4(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n401), .A2(new_n665), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n852), .A2(new_n859), .ZN(new_n860));
  OR2_X1    g0660(.A1(KEYINPUT100), .A2(KEYINPUT16), .ZN(new_n861));
  AND3_X1   g0661(.A1(new_n265), .A2(new_n268), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n861), .B1(new_n265), .B2(new_n268), .ZN(new_n863));
  OR3_X1    g0663(.A1(new_n862), .A2(new_n863), .A3(new_n254), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n314), .A2(new_n316), .B1(new_n284), .B2(new_n864), .ZN(new_n865));
  NOR3_X1   g0665(.A1(new_n862), .A2(new_n863), .A3(new_n254), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n848), .B1(new_n866), .B2(new_n283), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n304), .ZN(new_n868));
  OAI21_X1  g0668(.A(KEYINPUT37), .B1(new_n865), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(KEYINPUT101), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n318), .B1(new_n317), .B2(new_n848), .ZN(new_n871));
  XOR2_X1   g0671(.A(KEYINPUT102), .B(KEYINPUT37), .Z(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n871), .A2(new_n304), .A3(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT101), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n875), .B(KEYINPUT37), .C1(new_n865), .C2(new_n868), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n870), .A2(new_n874), .A3(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n867), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n324), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT38), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n877), .A2(new_n879), .A3(KEYINPUT38), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n850), .B1(new_n860), .B2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n882), .A2(KEYINPUT39), .A3(new_n883), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT105), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n883), .A2(new_n887), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n877), .A2(new_n879), .A3(KEYINPUT105), .A4(KEYINPUT38), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n871), .A2(KEYINPUT104), .A3(new_n304), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n318), .B1(new_n320), .B2(new_n321), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n318), .A2(new_n848), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n891), .A2(new_n304), .A3(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT104), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n890), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT103), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n871), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n872), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n890), .A2(new_n895), .A3(new_n898), .A4(new_n872), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n324), .A2(new_n318), .A3(new_n848), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  AOI22_X1  g0703(.A1(new_n888), .A2(new_n889), .B1(new_n903), .B2(new_n881), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n886), .B1(new_n904), .B2(KEYINPUT39), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n442), .A2(new_n665), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n885), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n704), .A2(new_n446), .A3(new_n707), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n637), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n909), .B(new_n911), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n722), .A2(new_n723), .A3(new_n822), .A4(new_n858), .ZN(new_n913));
  OAI21_X1  g0713(.A(KEYINPUT40), .B1(new_n904), .B2(new_n913), .ZN(new_n914));
  AND4_X1   g0714(.A1(new_n722), .A2(new_n723), .A3(new_n822), .A4(new_n858), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT40), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n915), .A2(new_n916), .A3(new_n884), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n724), .A2(new_n447), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n919), .B(KEYINPUT106), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n918), .B(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(G330), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n912), .B(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n203), .B2(new_n659), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT35), .ZN(new_n925));
  AOI211_X1 g0725(.A(new_n231), .B(new_n230), .C1(new_n582), .C2(new_n925), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n926), .B(G116), .C1(new_n925), .C2(new_n582), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT36), .ZN(new_n928));
  OAI21_X1  g0728(.A(G77), .B1(new_n222), .B2(new_n363), .ZN(new_n929));
  OAI22_X1  g0729(.A1(new_n929), .A2(new_n232), .B1(G50), .B2(new_n363), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n930), .A2(G1), .A3(new_n658), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n924), .A2(new_n928), .A3(new_n931), .ZN(G367));
  NAND2_X1  g0732(.A1(new_n683), .A2(new_n679), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n638), .B1(new_n594), .B2(new_n676), .ZN(new_n934));
  INV_X1    g0734(.A(new_n594), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n935), .A2(new_n620), .A3(new_n621), .A4(new_n665), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n933), .A2(new_n938), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT45), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n933), .A2(new_n938), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT44), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n941), .B(new_n942), .ZN(new_n943));
  AND3_X1   g0743(.A1(new_n940), .A2(new_n678), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n678), .B1(new_n940), .B2(new_n943), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n683), .B1(new_n677), .B2(new_n680), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n671), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n802), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n948), .B1(new_n949), .B2(new_n947), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n946), .A2(new_n727), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n727), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n686), .B(KEYINPUT41), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n780), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n560), .A2(new_n676), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n647), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n578), .B2(new_n955), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n957), .B(KEYINPUT107), .Z(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n682), .A2(new_n638), .ZN(new_n960));
  XOR2_X1   g0760(.A(KEYINPUT108), .B(KEYINPUT42), .Z(new_n961));
  XOR2_X1   g0761(.A(new_n960), .B(new_n961), .Z(new_n962));
  OAI21_X1  g0762(.A(new_n622), .B1(new_n938), .B2(new_n512), .ZN(new_n963));
  AND2_X1   g0763(.A1(new_n963), .A2(new_n676), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n959), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n965), .A2(new_n966), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n678), .A2(new_n938), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n970), .B(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n958), .A2(new_n796), .ZN(new_n973));
  INV_X1    g0773(.A(G150), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n747), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n765), .A2(G77), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n772), .A2(G137), .ZN(new_n977));
  AOI22_X1  g0777(.A1(G58), .A2(new_n827), .B1(new_n751), .B2(G68), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n976), .A2(new_n326), .A3(new_n977), .A4(new_n978), .ZN(new_n979));
  AOI211_X1 g0779(.A(new_n975), .B(new_n979), .C1(G143), .C2(new_n767), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n980), .B1(new_n217), .B2(new_n740), .C1(new_n742), .C2(new_n756), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n756), .A2(new_n489), .B1(new_n213), .B2(new_n761), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n759), .A2(new_n763), .ZN(new_n983));
  AOI21_X1  g0783(.A(KEYINPUT46), .B1(new_n827), .B2(G116), .ZN(new_n984));
  NOR4_X1   g0784(.A1(new_n982), .A2(new_n326), .A3(new_n983), .A4(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n739), .A2(G283), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n827), .A2(KEYINPUT46), .A3(G116), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT109), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n748), .A2(G303), .B1(G317), .B2(new_n772), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n985), .A2(new_n986), .A3(new_n988), .A4(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n735), .A2(new_n209), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n981), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT47), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n729), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n786), .B1(new_n234), .B2(new_n557), .C1(new_n244), .C2(new_n789), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n994), .A2(new_n781), .A3(new_n995), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n954), .A2(new_n972), .B1(new_n973), .B2(new_n996), .ZN(G387));
  OR2_X1    g0797(.A1(new_n950), .A2(new_n727), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n950), .A2(new_n727), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n998), .A2(new_n686), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n950), .A2(new_n780), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n788), .B1(new_n241), .B2(new_n776), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n688), .A2(new_n234), .A3(new_n326), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NOR3_X1   g0804(.A1(new_n277), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n1005), .A2(G45), .ZN(new_n1006));
  OAI21_X1  g0806(.A(KEYINPUT50), .B1(new_n277), .B2(G50), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n1006), .B(new_n1007), .C1(new_n363), .C2(new_n219), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1004), .B1(new_n688), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n685), .A2(new_n213), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n787), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n759), .A2(new_n742), .B1(new_n219), .B2(new_n754), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n258), .B(new_n1012), .C1(G50), .C2(new_n748), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n991), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n739), .A2(G68), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n741), .A2(new_n974), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n761), .A2(new_n557), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n1016), .B(new_n1017), .C1(new_n276), .C2(new_n755), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .A4(new_n1018), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n755), .A2(G311), .B1(new_n748), .B2(G317), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n767), .A2(G322), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n1020), .B(new_n1021), .C1(new_n517), .C2(new_n740), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT48), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1023), .B1(new_n839), .B2(new_n761), .C1(new_n489), .C2(new_n754), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT49), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n765), .A2(G116), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n772), .A2(G326), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1026), .A2(new_n258), .A3(new_n1027), .A4(new_n1028), .ZN(new_n1029));
  AND2_X1   g0829(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1019), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1011), .B1(new_n1031), .B2(new_n729), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1032), .B(new_n781), .C1(new_n677), .C2(new_n796), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1000), .A2(new_n1001), .A3(new_n1033), .ZN(G393));
  OAI21_X1  g0834(.A(new_n999), .B1(new_n944), .B2(new_n945), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n951), .A2(new_n686), .A3(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n786), .B1(new_n209), .B2(new_n234), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(new_n788), .B2(new_n251), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1038), .B(KEYINPUT110), .Z(new_n1039));
  AND2_X1   g0839(.A1(new_n772), .A2(G322), .ZN(new_n1040));
  INV_X1    g0840(.A(G317), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n763), .A2(new_n747), .B1(new_n759), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT52), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n326), .B(new_n1040), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1044), .B1(new_n525), .B2(new_n761), .C1(new_n839), .C2(new_n754), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n756), .A2(new_n517), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n740), .A2(new_n489), .B1(new_n735), .B2(new_n213), .ZN(new_n1048));
  NOR4_X1   g0848(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n739), .A2(new_n276), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n258), .B1(new_n751), .B2(G77), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n827), .A2(G68), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(G50), .B2(new_n755), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n765), .A2(G87), .B1(G143), .B2(new_n772), .ZN(new_n1055));
  AND2_X1   g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n974), .A2(new_n759), .B1(new_n747), .B2(new_n742), .ZN(new_n1057));
  XOR2_X1   g0857(.A(KEYINPUT111), .B(KEYINPUT51), .Z(new_n1058));
  XNOR2_X1  g0858(.A(new_n1057), .B(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1049), .B1(new_n1056), .B2(new_n1059), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n1060), .B(KEYINPUT112), .Z(new_n1061));
  OAI211_X1 g0861(.A(new_n781), .B(new_n1039), .C1(new_n1061), .C2(new_n730), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(new_n785), .B2(new_n938), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(new_n946), .B2(new_n780), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1036), .A2(new_n1064), .ZN(G390));
  INV_X1    g0865(.A(G128), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n326), .B1(new_n759), .B2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(G132), .B2(new_n748), .ZN(new_n1068));
  XOR2_X1   g0868(.A(KEYINPUT54), .B(G143), .Z(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1068), .B1(new_n217), .B2(new_n735), .C1(new_n740), .C2(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(G125), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n741), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n827), .A2(G150), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT53), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n756), .A2(new_n830), .B1(new_n742), .B2(new_n761), .ZN(new_n1076));
  NOR4_X1   g0876(.A1(new_n1071), .A2(new_n1073), .A3(new_n1075), .A4(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n765), .A2(G68), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n827), .A2(G87), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n739), .A2(G97), .B1(G77), .B2(new_n751), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1078), .A2(new_n258), .A3(new_n1079), .A4(new_n1080), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n741), .A2(new_n489), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n756), .A2(new_n213), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n525), .A2(new_n747), .B1(new_n759), .B2(new_n839), .ZN(new_n1084));
  NOR4_X1   g0884(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .A4(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n729), .B1(new_n1077), .B2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n781), .B1(new_n276), .B2(new_n825), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT120), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1086), .B(new_n1088), .C1(new_n906), .C2(new_n784), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT114), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n888), .A2(new_n889), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n903), .A2(new_n881), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n907), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n858), .A2(KEYINPUT113), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT113), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n856), .A2(new_n1097), .A3(new_n857), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n703), .A2(new_n676), .A3(new_n822), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n851), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1099), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1090), .B1(new_n1095), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1099), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n665), .B(new_n817), .C1(new_n701), .C2(new_n702), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1104), .B1(new_n1105), .B2(new_n851), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n904), .A2(new_n907), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1106), .A2(new_n1107), .A3(KEYINPUT114), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1094), .B1(new_n852), .B2(new_n859), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n1103), .A2(new_n1108), .B1(new_n1109), .B2(new_n905), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n915), .A2(G330), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1110), .A2(KEYINPUT115), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1111), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1109), .A2(new_n905), .ZN(new_n1114));
  NOR3_X1   g0914(.A1(new_n1095), .A2(new_n1102), .A3(new_n1090), .ZN(new_n1115));
  AOI21_X1  g0915(.A(KEYINPUT114), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1114), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT115), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1113), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1112), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n780), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1089), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT119), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n852), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n722), .A2(new_n723), .A3(G330), .A4(new_n822), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n859), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(new_n725), .B2(new_n913), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n915), .A2(G330), .B1(new_n1127), .B2(new_n1099), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n665), .B1(new_n701), .B2(new_n702), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n851), .B1(new_n1131), .B2(new_n822), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n1126), .A2(new_n1129), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT117), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n446), .A2(new_n722), .A3(G330), .A4(new_n723), .ZN(new_n1135));
  AND2_X1   g0935(.A1(new_n1135), .A2(KEYINPUT116), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1135), .A2(KEYINPUT116), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n637), .B(new_n910), .C1(new_n1136), .C2(new_n1137), .ZN(new_n1138));
  NOR3_X1   g0938(.A1(new_n1133), .A2(new_n1134), .A3(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1127), .A2(new_n1099), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1111), .A2(new_n1132), .A3(new_n1140), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n915), .A2(G330), .B1(new_n1127), .B2(new_n859), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1141), .B1(new_n852), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT116), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1135), .B(new_n1144), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1145), .A2(new_n911), .ZN(new_n1146));
  AOI21_X1  g0946(.A(KEYINPUT117), .B1(new_n1143), .B2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(KEYINPUT118), .B1(new_n1139), .B2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1134), .B1(new_n1133), .B2(new_n1138), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT118), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1143), .A2(new_n1146), .A3(KEYINPUT117), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1148), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n1121), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1112), .B(new_n1155), .C1(new_n1119), .C2(new_n1120), .ZN(new_n1156));
  AND4_X1   g0956(.A1(new_n1125), .A2(new_n1154), .A3(new_n686), .A4(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n686), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(new_n1153), .B2(new_n1121), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1125), .B1(new_n1159), .B2(new_n1156), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1124), .B1(new_n1157), .B2(new_n1160), .ZN(G378));
  XNOR2_X1  g0961(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n435), .B(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n663), .B1(new_n418), .B2(new_n423), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1163), .B(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n781), .B1(new_n1165), .B2(new_n784), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(new_n217), .B2(new_n824), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n735), .A2(new_n222), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1168), .B(KEYINPUT121), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n767), .A2(G116), .B1(G68), .B2(new_n751), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n1171), .A2(KEYINPUT122), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1171), .A2(KEYINPUT122), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n1172), .A2(new_n1173), .B1(new_n219), .B2(new_n754), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n286), .B1(new_n756), .B2(new_n209), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n258), .B1(new_n740), .B2(new_n557), .ZN(new_n1176));
  NOR4_X1   g0976(.A1(new_n1170), .A2(new_n1174), .A3(new_n1175), .A4(new_n1176), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n1177), .B1(new_n213), .B2(new_n747), .C1(new_n839), .C2(new_n741), .ZN(new_n1178));
  XOR2_X1   g0978(.A(new_n1178), .B(KEYINPUT123), .Z(new_n1179));
  XNOR2_X1  g0979(.A(new_n1179), .B(KEYINPUT58), .ZN(new_n1180));
  INV_X1    g0980(.A(G124), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n285), .B1(new_n741), .B2(new_n1181), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n1072), .A2(new_n759), .B1(new_n747), .B2(new_n1066), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n755), .A2(G132), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(new_n754), .B2(new_n1070), .ZN(new_n1185));
  AOI211_X1 g0985(.A(new_n1183), .B(new_n1185), .C1(G150), .C2(new_n751), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1186), .B1(new_n830), .B2(new_n740), .ZN(new_n1187));
  AOI211_X1 g0987(.A(G41), .B(new_n1182), .C1(new_n1187), .C2(KEYINPUT59), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n1188), .B1(KEYINPUT59), .B2(new_n1187), .C1(new_n742), .C2(new_n735), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n217), .B1(new_n256), .B2(G41), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n729), .B1(new_n1180), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1167), .A2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1165), .B1(new_n918), .B2(new_n725), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n914), .A2(new_n917), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1165), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1195), .A2(G330), .A3(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1194), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n885), .A2(new_n908), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n909), .A2(new_n1197), .A3(new_n1194), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1193), .B1(new_n1202), .B2(new_n1122), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1156), .A2(new_n1146), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1202), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1205), .A2(KEYINPUT57), .A3(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(new_n686), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1202), .B1(new_n1156), .B2(new_n1146), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1209), .A2(KEYINPUT57), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1204), .B1(new_n1208), .B2(new_n1210), .ZN(G375));
  NAND2_X1  g1011(.A1(new_n1133), .A2(new_n1138), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1153), .A2(new_n953), .A3(new_n1212), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n1104), .A2(new_n784), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n976), .B1(new_n209), .B2(new_n754), .C1(new_n517), .C2(new_n741), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n1017), .B(new_n1215), .C1(G116), .C2(new_n755), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n258), .B1(new_n747), .B2(new_n839), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(G294), .B2(new_n767), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n1216), .B(new_n1218), .C1(new_n213), .C2(new_n740), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1219), .B(KEYINPUT124), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n740), .A2(new_n974), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n767), .A2(G132), .B1(G50), .B2(new_n751), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n742), .B2(new_n754), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n326), .B1(new_n741), .B2(new_n1066), .ZN(new_n1224));
  NOR4_X1   g1024(.A1(new_n1170), .A2(new_n1221), .A3(new_n1223), .A4(new_n1224), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n1225), .B1(new_n830), .B2(new_n747), .C1(new_n756), .C2(new_n1070), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n730), .B1(new_n1220), .B2(new_n1226), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n825), .A2(G68), .ZN(new_n1228));
  NOR4_X1   g1028(.A1(new_n1214), .A2(new_n782), .A3(new_n1227), .A4(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(new_n1143), .B2(new_n780), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1213), .A2(new_n1230), .ZN(G381));
  AOI21_X1  g1031(.A(new_n1158), .B1(new_n1209), .B2(KEYINPUT57), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT57), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1103), .A2(new_n1108), .ZN(new_n1234));
  AND4_X1   g1034(.A1(KEYINPUT115), .A2(new_n1234), .A3(new_n1114), .A4(new_n1111), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1110), .A2(KEYINPUT115), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1111), .B1(new_n1110), .B2(KEYINPUT115), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1235), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1138), .B1(new_n1238), .B2(new_n1155), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1233), .B1(new_n1239), .B2(new_n1202), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1203), .B1(new_n1232), .B2(new_n1240), .ZN(new_n1241));
  OR2_X1    g1041(.A1(new_n1241), .A2(KEYINPUT125), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(KEYINPUT125), .ZN(new_n1243));
  AND3_X1   g1043(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1150), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n686), .B(new_n1156), .C1(new_n1246), .C2(new_n1238), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n1124), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1242), .A2(new_n1243), .A3(new_n1249), .ZN(new_n1250));
  NOR3_X1   g1050(.A1(new_n1250), .A2(G384), .A3(G381), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(G387), .A2(G390), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  NOR3_X1   g1053(.A1(new_n1253), .A2(G396), .A3(G393), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1251), .A2(new_n1254), .ZN(G407));
  OAI211_X1 g1055(.A(G407), .B(G213), .C1(G343), .C2(new_n1250), .ZN(G409));
  XOR2_X1   g1056(.A(G393), .B(G396), .Z(new_n1257));
  NAND2_X1  g1057(.A1(G387), .A2(G390), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1257), .B1(new_n1259), .B2(new_n1252), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1257), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1253), .A2(new_n1261), .A3(new_n1258), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1260), .A2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(G213), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1264), .A2(G343), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1158), .B1(new_n1155), .B2(new_n1212), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1212), .A2(KEYINPUT126), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(KEYINPUT60), .ZN(new_n1268));
  OR2_X1    g1068(.A1(new_n1267), .A2(KEYINPUT60), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1266), .A2(new_n1268), .A3(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1270), .A2(G384), .A3(new_n1230), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(G384), .B1(new_n1270), .B2(new_n1230), .ZN(new_n1273));
  OAI211_X1 g1073(.A(G2897), .B(new_n1265), .C1(new_n1272), .C2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1270), .A2(new_n1230), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(new_n846), .ZN(new_n1276));
  INV_X1    g1076(.A(G2897), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1265), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n1276), .B(new_n1271), .C1(new_n1277), .C2(new_n1278), .ZN(new_n1279));
  AND2_X1   g1079(.A1(new_n1274), .A2(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1203), .B1(new_n1209), .B2(new_n953), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1248), .A2(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1282), .B1(G378), .B2(new_n1241), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1280), .B1(new_n1283), .B2(new_n1265), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  NOR3_X1   g1086(.A1(new_n1283), .A2(new_n1265), .A3(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT62), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1284), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT61), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1247), .A2(KEYINPUT119), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1159), .A2(new_n1125), .A3(new_n1156), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1123), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  OAI22_X1  g1093(.A1(G375), .A2(new_n1293), .B1(new_n1248), .B2(new_n1281), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1294), .A2(new_n1278), .A3(new_n1285), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1290), .B1(new_n1295), .B2(KEYINPUT62), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1263), .B1(new_n1289), .B2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1274), .A2(new_n1279), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1298), .B1(new_n1294), .B2(new_n1278), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1263), .B1(new_n1299), .B2(KEYINPUT127), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT127), .ZN(new_n1301));
  AOI21_X1  g1101(.A(KEYINPUT61), .B1(new_n1284), .B2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT63), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1295), .A2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1287), .A2(KEYINPUT63), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1300), .A2(new_n1302), .A3(new_n1304), .A4(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1297), .A2(new_n1306), .ZN(G405));
  NOR2_X1   g1107(.A1(new_n1241), .A2(new_n1248), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1308), .B1(G378), .B2(new_n1241), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1263), .A2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1263), .A2(new_n1309), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1311), .A2(new_n1285), .A3(new_n1312), .ZN(new_n1313));
  AND2_X1   g1113(.A1(new_n1263), .A2(new_n1309), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1286), .B1(new_n1314), .B2(new_n1310), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1313), .A2(new_n1315), .ZN(G402));
endmodule


