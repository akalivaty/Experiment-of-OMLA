

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  BUF_X1 U557 ( .A(n713), .Z(n714) );
  AND2_X2 U558 ( .A1(n527), .A2(G2104), .ZN(n888) );
  XNOR2_X1 U559 ( .A(KEYINPUT32), .B(KEYINPUT100), .ZN(n669) );
  NOR2_X2 U560 ( .A1(G164), .A2(G1384), .ZN(n692) );
  NAND2_X1 U561 ( .A1(n616), .A2(n615), .ZN(n992) );
  OR2_X1 U562 ( .A1(KEYINPUT33), .A2(n689), .ZN(n522) );
  AND2_X1 U563 ( .A1(n695), .A2(n694), .ZN(n523) );
  NOR2_X4 U564 ( .A1(n552), .A2(n551), .ZN(G160) );
  NOR2_X1 U565 ( .A1(n992), .A2(n623), .ZN(n624) );
  INV_X1 U566 ( .A(KEYINPUT29), .ZN(n642) );
  XNOR2_X1 U567 ( .A(n643), .B(n642), .ZN(n648) );
  XNOR2_X1 U568 ( .A(n670), .B(n669), .ZN(n679) );
  INV_X1 U569 ( .A(n975), .ZN(n694) );
  NOR2_X1 U570 ( .A1(G543), .A2(n537), .ZN(n538) );
  AND2_X1 U571 ( .A1(G2105), .A2(G2104), .ZN(n884) );
  NOR2_X1 U572 ( .A1(G651), .A2(n577), .ZN(n798) );
  NOR2_X1 U573 ( .A1(G2104), .A2(G2105), .ZN(n524) );
  XOR2_X1 U574 ( .A(KEYINPUT17), .B(n524), .Z(n712) );
  NAND2_X1 U575 ( .A1(n712), .A2(G138), .ZN(n531) );
  NAND2_X1 U576 ( .A1(G114), .A2(n884), .ZN(n526) );
  INV_X1 U577 ( .A(G2105), .ZN(n527) );
  NOR2_X1 U578 ( .A1(G2104), .A2(n527), .ZN(n713) );
  NAND2_X1 U579 ( .A1(G126), .A2(n713), .ZN(n525) );
  AND2_X1 U580 ( .A1(n526), .A2(n525), .ZN(n529) );
  NAND2_X1 U581 ( .A1(G102), .A2(n888), .ZN(n528) );
  AND2_X1 U582 ( .A1(n529), .A2(n528), .ZN(n530) );
  AND2_X1 U583 ( .A1(n531), .A2(n530), .ZN(G164) );
  NOR2_X1 U584 ( .A1(G651), .A2(G543), .ZN(n791) );
  NAND2_X1 U585 ( .A1(n791), .A2(G89), .ZN(n532) );
  XNOR2_X1 U586 ( .A(n532), .B(KEYINPUT4), .ZN(n535) );
  XNOR2_X1 U587 ( .A(G543), .B(KEYINPUT0), .ZN(n533) );
  XNOR2_X1 U588 ( .A(n533), .B(KEYINPUT65), .ZN(n577) );
  INV_X1 U589 ( .A(G651), .ZN(n537) );
  NOR2_X2 U590 ( .A1(n577), .A2(n537), .ZN(n794) );
  NAND2_X1 U591 ( .A1(G76), .A2(n794), .ZN(n534) );
  NAND2_X1 U592 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U593 ( .A(n536), .B(KEYINPUT5), .ZN(n543) );
  XOR2_X1 U594 ( .A(KEYINPUT1), .B(n538), .Z(n790) );
  NAND2_X1 U595 ( .A1(G63), .A2(n790), .ZN(n540) );
  NAND2_X1 U596 ( .A1(G51), .A2(n798), .ZN(n539) );
  NAND2_X1 U597 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U598 ( .A(KEYINPUT6), .B(n541), .Z(n542) );
  NAND2_X1 U599 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U600 ( .A(n544), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U601 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U602 ( .A1(G101), .A2(n888), .ZN(n545) );
  XOR2_X1 U603 ( .A(KEYINPUT23), .B(n545), .Z(n548) );
  NAND2_X1 U604 ( .A1(G125), .A2(n713), .ZN(n546) );
  XNOR2_X1 U605 ( .A(n546), .B(KEYINPUT64), .ZN(n547) );
  NAND2_X1 U606 ( .A1(n548), .A2(n547), .ZN(n552) );
  NAND2_X1 U607 ( .A1(G137), .A2(n712), .ZN(n550) );
  NAND2_X1 U608 ( .A1(G113), .A2(n884), .ZN(n549) );
  NAND2_X1 U609 ( .A1(n550), .A2(n549), .ZN(n551) );
  NAND2_X1 U610 ( .A1(G78), .A2(n794), .ZN(n553) );
  XNOR2_X1 U611 ( .A(n553), .B(KEYINPUT70), .ZN(n560) );
  NAND2_X1 U612 ( .A1(G65), .A2(n790), .ZN(n555) );
  NAND2_X1 U613 ( .A1(G53), .A2(n798), .ZN(n554) );
  NAND2_X1 U614 ( .A1(n555), .A2(n554), .ZN(n558) );
  NAND2_X1 U615 ( .A1(G91), .A2(n791), .ZN(n556) );
  XNOR2_X1 U616 ( .A(KEYINPUT69), .B(n556), .ZN(n557) );
  NOR2_X1 U617 ( .A1(n558), .A2(n557), .ZN(n559) );
  NAND2_X1 U618 ( .A1(n560), .A2(n559), .ZN(G299) );
  NAND2_X1 U619 ( .A1(n794), .A2(G77), .ZN(n561) );
  XNOR2_X1 U620 ( .A(n561), .B(KEYINPUT68), .ZN(n563) );
  NAND2_X1 U621 ( .A1(G90), .A2(n791), .ZN(n562) );
  NAND2_X1 U622 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U623 ( .A(n564), .B(KEYINPUT9), .ZN(n566) );
  NAND2_X1 U624 ( .A1(G64), .A2(n790), .ZN(n565) );
  NAND2_X1 U625 ( .A1(n566), .A2(n565), .ZN(n569) );
  NAND2_X1 U626 ( .A1(G52), .A2(n798), .ZN(n567) );
  XNOR2_X1 U627 ( .A(KEYINPUT67), .B(n567), .ZN(n568) );
  NOR2_X1 U628 ( .A1(n569), .A2(n568), .ZN(G171) );
  NAND2_X1 U629 ( .A1(G75), .A2(n794), .ZN(n571) );
  NAND2_X1 U630 ( .A1(G88), .A2(n791), .ZN(n570) );
  NAND2_X1 U631 ( .A1(n571), .A2(n570), .ZN(n574) );
  NAND2_X1 U632 ( .A1(G62), .A2(n790), .ZN(n572) );
  XNOR2_X1 U633 ( .A(KEYINPUT83), .B(n572), .ZN(n573) );
  NOR2_X1 U634 ( .A1(n574), .A2(n573), .ZN(n576) );
  NAND2_X1 U635 ( .A1(n798), .A2(G50), .ZN(n575) );
  NAND2_X1 U636 ( .A1(n576), .A2(n575), .ZN(G303) );
  NAND2_X1 U637 ( .A1(G49), .A2(n798), .ZN(n579) );
  NAND2_X1 U638 ( .A1(G87), .A2(n577), .ZN(n578) );
  NAND2_X1 U639 ( .A1(n579), .A2(n578), .ZN(n580) );
  NOR2_X1 U640 ( .A1(n790), .A2(n580), .ZN(n582) );
  NAND2_X1 U641 ( .A1(G651), .A2(G74), .ZN(n581) );
  NAND2_X1 U642 ( .A1(n582), .A2(n581), .ZN(G288) );
  NAND2_X1 U643 ( .A1(G72), .A2(n794), .ZN(n584) );
  NAND2_X1 U644 ( .A1(G85), .A2(n791), .ZN(n583) );
  NAND2_X1 U645 ( .A1(n584), .A2(n583), .ZN(n587) );
  NAND2_X1 U646 ( .A1(n790), .A2(G60), .ZN(n585) );
  XOR2_X1 U647 ( .A(KEYINPUT66), .B(n585), .Z(n586) );
  NOR2_X1 U648 ( .A1(n587), .A2(n586), .ZN(n589) );
  NAND2_X1 U649 ( .A1(n798), .A2(G47), .ZN(n588) );
  NAND2_X1 U650 ( .A1(n589), .A2(n588), .ZN(G290) );
  NAND2_X1 U651 ( .A1(G86), .A2(n791), .ZN(n591) );
  NAND2_X1 U652 ( .A1(G48), .A2(n798), .ZN(n590) );
  NAND2_X1 U653 ( .A1(n591), .A2(n590), .ZN(n594) );
  NAND2_X1 U654 ( .A1(G73), .A2(n794), .ZN(n592) );
  XOR2_X1 U655 ( .A(KEYINPUT2), .B(n592), .Z(n593) );
  NOR2_X1 U656 ( .A1(n594), .A2(n593), .ZN(n596) );
  NAND2_X1 U657 ( .A1(n790), .A2(G61), .ZN(n595) );
  NAND2_X1 U658 ( .A1(n596), .A2(n595), .ZN(G305) );
  NAND2_X1 U659 ( .A1(G66), .A2(n790), .ZN(n597) );
  XNOR2_X1 U660 ( .A(n597), .B(KEYINPUT74), .ZN(n604) );
  NAND2_X1 U661 ( .A1(G79), .A2(n794), .ZN(n599) );
  NAND2_X1 U662 ( .A1(G54), .A2(n798), .ZN(n598) );
  NAND2_X1 U663 ( .A1(n599), .A2(n598), .ZN(n602) );
  NAND2_X1 U664 ( .A1(G92), .A2(n791), .ZN(n600) );
  XNOR2_X1 U665 ( .A(KEYINPUT75), .B(n600), .ZN(n601) );
  NOR2_X1 U666 ( .A1(n602), .A2(n601), .ZN(n603) );
  NAND2_X1 U667 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X2 U668 ( .A(KEYINPUT15), .B(n605), .ZN(n977) );
  XOR2_X1 U669 ( .A(KEYINPUT72), .B(KEYINPUT14), .Z(n607) );
  NAND2_X1 U670 ( .A1(G56), .A2(n790), .ZN(n606) );
  XNOR2_X1 U671 ( .A(n607), .B(n606), .ZN(n614) );
  NAND2_X1 U672 ( .A1(n794), .A2(G68), .ZN(n608) );
  XNOR2_X1 U673 ( .A(KEYINPUT73), .B(n608), .ZN(n611) );
  NAND2_X1 U674 ( .A1(n791), .A2(G81), .ZN(n609) );
  XOR2_X1 U675 ( .A(KEYINPUT12), .B(n609), .Z(n610) );
  NOR2_X1 U676 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U677 ( .A(n612), .B(KEYINPUT13), .ZN(n613) );
  NOR2_X1 U678 ( .A1(n614), .A2(n613), .ZN(n616) );
  NAND2_X1 U679 ( .A1(n798), .A2(G43), .ZN(n615) );
  AND2_X1 U680 ( .A1(G160), .A2(G40), .ZN(n618) );
  AND2_X2 U681 ( .A1(n618), .A2(n692), .ZN(n644) );
  NAND2_X1 U682 ( .A1(G1996), .A2(n644), .ZN(n617) );
  XNOR2_X1 U683 ( .A(n617), .B(KEYINPUT26), .ZN(n620) );
  NAND2_X1 U684 ( .A1(n692), .A2(n618), .ZN(n658) );
  NAND2_X1 U685 ( .A1(G1341), .A2(n658), .ZN(n619) );
  NAND2_X1 U686 ( .A1(n620), .A2(n619), .ZN(n622) );
  INV_X1 U687 ( .A(KEYINPUT95), .ZN(n621) );
  XNOR2_X1 U688 ( .A(n622), .B(n621), .ZN(n623) );
  OR2_X1 U689 ( .A1(n977), .A2(n624), .ZN(n631) );
  NAND2_X1 U690 ( .A1(n977), .A2(n624), .ZN(n629) );
  NAND2_X1 U691 ( .A1(n658), .A2(G1348), .ZN(n625) );
  XNOR2_X1 U692 ( .A(n625), .B(KEYINPUT96), .ZN(n627) );
  NAND2_X1 U693 ( .A1(n644), .A2(G2067), .ZN(n626) );
  NAND2_X1 U694 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X1 U695 ( .A1(n629), .A2(n628), .ZN(n630) );
  NAND2_X1 U696 ( .A1(n631), .A2(n630), .ZN(n636) );
  NAND2_X1 U697 ( .A1(n644), .A2(G2072), .ZN(n632) );
  XNOR2_X1 U698 ( .A(n632), .B(KEYINPUT27), .ZN(n634) );
  INV_X1 U699 ( .A(G1956), .ZN(n1004) );
  NOR2_X1 U700 ( .A1(n1004), .A2(n644), .ZN(n633) );
  NOR2_X1 U701 ( .A1(n634), .A2(n633), .ZN(n637) );
  INV_X1 U702 ( .A(G299), .ZN(n978) );
  NAND2_X1 U703 ( .A1(n637), .A2(n978), .ZN(n635) );
  NAND2_X1 U704 ( .A1(n636), .A2(n635), .ZN(n641) );
  NOR2_X1 U705 ( .A1(n637), .A2(n978), .ZN(n639) );
  XOR2_X1 U706 ( .A(KEYINPUT94), .B(KEYINPUT28), .Z(n638) );
  XNOR2_X1 U707 ( .A(n639), .B(n638), .ZN(n640) );
  NAND2_X1 U708 ( .A1(n641), .A2(n640), .ZN(n643) );
  XNOR2_X1 U709 ( .A(G1961), .B(KEYINPUT93), .ZN(n1014) );
  NAND2_X1 U710 ( .A1(n658), .A2(n1014), .ZN(n646) );
  XNOR2_X1 U711 ( .A(G2078), .B(KEYINPUT25), .ZN(n961) );
  NAND2_X1 U712 ( .A1(n644), .A2(n961), .ZN(n645) );
  NAND2_X1 U713 ( .A1(n646), .A2(n645), .ZN(n649) );
  NAND2_X1 U714 ( .A1(n649), .A2(G171), .ZN(n647) );
  NAND2_X1 U715 ( .A1(n648), .A2(n647), .ZN(n657) );
  NOR2_X1 U716 ( .A1(G171), .A2(n649), .ZN(n654) );
  NAND2_X1 U717 ( .A1(G8), .A2(n658), .ZN(n703) );
  NOR2_X1 U718 ( .A1(G1966), .A2(n703), .ZN(n675) );
  NOR2_X1 U719 ( .A1(G2084), .A2(n658), .ZN(n671) );
  NOR2_X1 U720 ( .A1(n675), .A2(n671), .ZN(n650) );
  NAND2_X1 U721 ( .A1(G8), .A2(n650), .ZN(n651) );
  XNOR2_X1 U722 ( .A(KEYINPUT30), .B(n651), .ZN(n652) );
  NOR2_X1 U723 ( .A1(G168), .A2(n652), .ZN(n653) );
  NOR2_X1 U724 ( .A1(n654), .A2(n653), .ZN(n655) );
  XOR2_X1 U725 ( .A(KEYINPUT31), .B(n655), .Z(n656) );
  NAND2_X1 U726 ( .A1(n657), .A2(n656), .ZN(n673) );
  NAND2_X1 U727 ( .A1(n673), .A2(G286), .ZN(n665) );
  NOR2_X1 U728 ( .A1(n658), .A2(G2090), .ZN(n659) );
  XNOR2_X1 U729 ( .A(n659), .B(KEYINPUT98), .ZN(n662) );
  NOR2_X1 U730 ( .A1(G1971), .A2(n703), .ZN(n660) );
  XOR2_X1 U731 ( .A(KEYINPUT97), .B(n660), .Z(n661) );
  NOR2_X1 U732 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U733 ( .A1(n663), .A2(G303), .ZN(n664) );
  NAND2_X1 U734 ( .A1(n665), .A2(n664), .ZN(n667) );
  INV_X1 U735 ( .A(KEYINPUT99), .ZN(n666) );
  XNOR2_X1 U736 ( .A(n667), .B(n666), .ZN(n668) );
  NAND2_X1 U737 ( .A1(n668), .A2(G8), .ZN(n670) );
  NAND2_X1 U738 ( .A1(G8), .A2(n671), .ZN(n672) );
  XNOR2_X1 U739 ( .A(KEYINPUT92), .B(n672), .ZN(n677) );
  INV_X1 U740 ( .A(n673), .ZN(n674) );
  NOR2_X1 U741 ( .A1(n675), .A2(n674), .ZN(n676) );
  NAND2_X1 U742 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U743 ( .A1(n679), .A2(n678), .ZN(n681) );
  INV_X1 U744 ( .A(KEYINPUT101), .ZN(n680) );
  XNOR2_X1 U745 ( .A(n681), .B(n680), .ZN(n696) );
  NOR2_X1 U746 ( .A1(G1976), .A2(G288), .ZN(n682) );
  XOR2_X1 U747 ( .A(KEYINPUT102), .B(n682), .Z(n981) );
  NOR2_X1 U748 ( .A1(G1971), .A2(G303), .ZN(n683) );
  XNOR2_X1 U749 ( .A(n683), .B(KEYINPUT103), .ZN(n684) );
  AND2_X1 U750 ( .A1(n981), .A2(n684), .ZN(n685) );
  NAND2_X1 U751 ( .A1(n696), .A2(n685), .ZN(n686) );
  XNOR2_X1 U752 ( .A(n686), .B(KEYINPUT104), .ZN(n687) );
  NAND2_X1 U753 ( .A1(G1976), .A2(G288), .ZN(n982) );
  NAND2_X1 U754 ( .A1(n687), .A2(n982), .ZN(n688) );
  NOR2_X1 U755 ( .A1(n688), .A2(n703), .ZN(n689) );
  NOR2_X1 U756 ( .A1(n703), .A2(n981), .ZN(n690) );
  NAND2_X1 U757 ( .A1(KEYINPUT33), .A2(n690), .ZN(n693) );
  NAND2_X1 U758 ( .A1(G160), .A2(G40), .ZN(n691) );
  NOR2_X1 U759 ( .A1(n692), .A2(n691), .ZN(n759) );
  XNOR2_X1 U760 ( .A(G1986), .B(G290), .ZN(n985) );
  NAND2_X1 U761 ( .A1(n759), .A2(n985), .ZN(n706) );
  AND2_X1 U762 ( .A1(n693), .A2(n706), .ZN(n695) );
  XNOR2_X1 U763 ( .A(G1981), .B(G305), .ZN(n975) );
  NAND2_X1 U764 ( .A1(n522), .A2(n523), .ZN(n710) );
  NOR2_X1 U765 ( .A1(G2090), .A2(G303), .ZN(n697) );
  NAND2_X1 U766 ( .A1(G8), .A2(n697), .ZN(n698) );
  NAND2_X1 U767 ( .A1(n696), .A2(n698), .ZN(n699) );
  NAND2_X1 U768 ( .A1(n703), .A2(n699), .ZN(n700) );
  XNOR2_X1 U769 ( .A(n700), .B(KEYINPUT105), .ZN(n705) );
  NOR2_X1 U770 ( .A1(G1981), .A2(G305), .ZN(n701) );
  XOR2_X1 U771 ( .A(n701), .B(KEYINPUT24), .Z(n702) );
  NOR2_X1 U772 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U773 ( .A1(n705), .A2(n704), .ZN(n708) );
  INV_X1 U774 ( .A(n706), .ZN(n707) );
  OR2_X1 U775 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U776 ( .A1(n710), .A2(n709), .ZN(n745) );
  INV_X1 U777 ( .A(G1996), .ZN(n954) );
  NAND2_X1 U778 ( .A1(G105), .A2(n888), .ZN(n711) );
  XNOR2_X1 U779 ( .A(n711), .B(KEYINPUT38), .ZN(n721) );
  BUF_X1 U780 ( .A(n712), .Z(n887) );
  NAND2_X1 U781 ( .A1(G141), .A2(n887), .ZN(n716) );
  NAND2_X1 U782 ( .A1(G129), .A2(n714), .ZN(n715) );
  NAND2_X1 U783 ( .A1(n716), .A2(n715), .ZN(n719) );
  NAND2_X1 U784 ( .A1(G117), .A2(n884), .ZN(n717) );
  XNOR2_X1 U785 ( .A(KEYINPUT89), .B(n717), .ZN(n718) );
  NOR2_X1 U786 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U787 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U788 ( .A(KEYINPUT90), .B(n722), .ZN(n870) );
  INV_X1 U789 ( .A(n870), .ZN(n723) );
  NOR2_X1 U790 ( .A1(n954), .A2(n723), .ZN(n731) );
  NAND2_X1 U791 ( .A1(G131), .A2(n887), .ZN(n725) );
  NAND2_X1 U792 ( .A1(G95), .A2(n888), .ZN(n724) );
  NAND2_X1 U793 ( .A1(n725), .A2(n724), .ZN(n729) );
  NAND2_X1 U794 ( .A1(G107), .A2(n884), .ZN(n727) );
  NAND2_X1 U795 ( .A1(G119), .A2(n714), .ZN(n726) );
  NAND2_X1 U796 ( .A1(n727), .A2(n726), .ZN(n728) );
  OR2_X1 U797 ( .A1(n729), .A2(n728), .ZN(n874) );
  AND2_X1 U798 ( .A1(G1991), .A2(n874), .ZN(n730) );
  NOR2_X1 U799 ( .A1(n731), .A2(n730), .ZN(n934) );
  XNOR2_X1 U800 ( .A(KEYINPUT91), .B(n759), .ZN(n732) );
  NOR2_X1 U801 ( .A1(n934), .A2(n732), .ZN(n750) );
  INV_X1 U802 ( .A(n750), .ZN(n743) );
  XNOR2_X1 U803 ( .A(KEYINPUT37), .B(G2067), .ZN(n755) );
  NAND2_X1 U804 ( .A1(n884), .A2(G116), .ZN(n733) );
  XNOR2_X1 U805 ( .A(n733), .B(KEYINPUT88), .ZN(n735) );
  NAND2_X1 U806 ( .A1(G128), .A2(n714), .ZN(n734) );
  NAND2_X1 U807 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U808 ( .A(n736), .B(KEYINPUT35), .ZN(n741) );
  NAND2_X1 U809 ( .A1(G140), .A2(n887), .ZN(n738) );
  NAND2_X1 U810 ( .A1(G104), .A2(n888), .ZN(n737) );
  NAND2_X1 U811 ( .A1(n738), .A2(n737), .ZN(n739) );
  XOR2_X1 U812 ( .A(KEYINPUT34), .B(n739), .Z(n740) );
  NAND2_X1 U813 ( .A1(n741), .A2(n740), .ZN(n742) );
  XOR2_X1 U814 ( .A(n742), .B(KEYINPUT36), .Z(n902) );
  NOR2_X1 U815 ( .A1(n755), .A2(n902), .ZN(n936) );
  NAND2_X1 U816 ( .A1(n759), .A2(n936), .ZN(n753) );
  NAND2_X1 U817 ( .A1(n743), .A2(n753), .ZN(n744) );
  NOR2_X1 U818 ( .A1(n745), .A2(n744), .ZN(n762) );
  NOR2_X1 U819 ( .A1(G1996), .A2(n870), .ZN(n927) );
  NOR2_X1 U820 ( .A1(G1991), .A2(n874), .ZN(n746) );
  XOR2_X1 U821 ( .A(KEYINPUT107), .B(n746), .Z(n932) );
  NOR2_X1 U822 ( .A1(G1986), .A2(G290), .ZN(n747) );
  XNOR2_X1 U823 ( .A(KEYINPUT106), .B(n747), .ZN(n748) );
  NOR2_X1 U824 ( .A1(n932), .A2(n748), .ZN(n749) );
  NOR2_X1 U825 ( .A1(n750), .A2(n749), .ZN(n751) );
  NOR2_X1 U826 ( .A1(n927), .A2(n751), .ZN(n752) );
  XNOR2_X1 U827 ( .A(KEYINPUT39), .B(n752), .ZN(n754) );
  NAND2_X1 U828 ( .A1(n754), .A2(n753), .ZN(n757) );
  AND2_X1 U829 ( .A1(n755), .A2(n902), .ZN(n756) );
  XOR2_X1 U830 ( .A(KEYINPUT108), .B(n756), .Z(n943) );
  NAND2_X1 U831 ( .A1(n757), .A2(n943), .ZN(n758) );
  NAND2_X1 U832 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U833 ( .A(n760), .B(KEYINPUT109), .ZN(n761) );
  OR2_X1 U834 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U835 ( .A(n763), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U836 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U837 ( .A1(G135), .A2(n887), .ZN(n765) );
  NAND2_X1 U838 ( .A1(G111), .A2(n884), .ZN(n764) );
  NAND2_X1 U839 ( .A1(n765), .A2(n764), .ZN(n770) );
  XOR2_X1 U840 ( .A(KEYINPUT18), .B(KEYINPUT79), .Z(n767) );
  NAND2_X1 U841 ( .A1(G123), .A2(n714), .ZN(n766) );
  XNOR2_X1 U842 ( .A(n767), .B(n766), .ZN(n768) );
  XOR2_X1 U843 ( .A(KEYINPUT78), .B(n768), .Z(n769) );
  NOR2_X1 U844 ( .A1(n770), .A2(n769), .ZN(n772) );
  NAND2_X1 U845 ( .A1(n888), .A2(G99), .ZN(n771) );
  NAND2_X1 U846 ( .A1(n772), .A2(n771), .ZN(n929) );
  XNOR2_X1 U847 ( .A(G2096), .B(n929), .ZN(n773) );
  OR2_X1 U848 ( .A1(G2100), .A2(n773), .ZN(G156) );
  INV_X1 U849 ( .A(G57), .ZN(G237) );
  INV_X1 U850 ( .A(G132), .ZN(G219) );
  INV_X1 U851 ( .A(G82), .ZN(G220) );
  NAND2_X1 U852 ( .A1(G7), .A2(G661), .ZN(n774) );
  XNOR2_X1 U853 ( .A(n774), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U854 ( .A(G223), .ZN(n834) );
  NAND2_X1 U855 ( .A1(n834), .A2(G567), .ZN(n775) );
  XNOR2_X1 U856 ( .A(n775), .B(KEYINPUT71), .ZN(n776) );
  XNOR2_X1 U857 ( .A(KEYINPUT11), .B(n776), .ZN(G234) );
  INV_X1 U858 ( .A(n992), .ZN(n777) );
  NAND2_X1 U859 ( .A1(n777), .A2(G860), .ZN(G153) );
  INV_X1 U860 ( .A(G171), .ZN(G301) );
  NAND2_X1 U861 ( .A1(G868), .A2(G301), .ZN(n779) );
  OR2_X1 U862 ( .A1(n977), .A2(G868), .ZN(n778) );
  NAND2_X1 U863 ( .A1(n779), .A2(n778), .ZN(G284) );
  INV_X1 U864 ( .A(G868), .ZN(n815) );
  NOR2_X1 U865 ( .A1(G286), .A2(n815), .ZN(n780) );
  XNOR2_X1 U866 ( .A(n780), .B(KEYINPUT76), .ZN(n782) );
  NOR2_X1 U867 ( .A1(G299), .A2(G868), .ZN(n781) );
  NOR2_X1 U868 ( .A1(n782), .A2(n781), .ZN(G297) );
  INV_X1 U869 ( .A(G559), .ZN(n783) );
  NOR2_X1 U870 ( .A1(G860), .A2(n783), .ZN(n784) );
  XNOR2_X1 U871 ( .A(KEYINPUT77), .B(n784), .ZN(n785) );
  NAND2_X1 U872 ( .A1(n785), .A2(n977), .ZN(n786) );
  XNOR2_X1 U873 ( .A(n786), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U874 ( .A1(G868), .A2(n992), .ZN(n789) );
  NAND2_X1 U875 ( .A1(G868), .A2(n977), .ZN(n787) );
  NOR2_X1 U876 ( .A1(G559), .A2(n787), .ZN(n788) );
  NOR2_X1 U877 ( .A1(n789), .A2(n788), .ZN(G282) );
  NAND2_X1 U878 ( .A1(G67), .A2(n790), .ZN(n793) );
  NAND2_X1 U879 ( .A1(G93), .A2(n791), .ZN(n792) );
  NAND2_X1 U880 ( .A1(n793), .A2(n792), .ZN(n797) );
  NAND2_X1 U881 ( .A1(n794), .A2(G80), .ZN(n795) );
  XOR2_X1 U882 ( .A(KEYINPUT82), .B(n795), .Z(n796) );
  NOR2_X1 U883 ( .A1(n797), .A2(n796), .ZN(n800) );
  NAND2_X1 U884 ( .A1(n798), .A2(G55), .ZN(n799) );
  NAND2_X1 U885 ( .A1(n800), .A2(n799), .ZN(n814) );
  NAND2_X1 U886 ( .A1(G559), .A2(n977), .ZN(n801) );
  XNOR2_X1 U887 ( .A(n801), .B(KEYINPUT80), .ZN(n812) );
  XOR2_X1 U888 ( .A(n812), .B(KEYINPUT81), .Z(n802) );
  XNOR2_X1 U889 ( .A(n992), .B(n802), .ZN(n803) );
  NOR2_X1 U890 ( .A1(G860), .A2(n803), .ZN(n804) );
  XOR2_X1 U891 ( .A(n814), .B(n804), .Z(G145) );
  INV_X1 U892 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U893 ( .A(G166), .B(G290), .ZN(n811) );
  XNOR2_X1 U894 ( .A(KEYINPUT19), .B(KEYINPUT84), .ZN(n805) );
  XOR2_X1 U895 ( .A(n805), .B(n814), .Z(n808) );
  XNOR2_X1 U896 ( .A(n978), .B(G305), .ZN(n806) );
  XNOR2_X1 U897 ( .A(n806), .B(n992), .ZN(n807) );
  XNOR2_X1 U898 ( .A(n808), .B(n807), .ZN(n809) );
  XNOR2_X1 U899 ( .A(n809), .B(G288), .ZN(n810) );
  XNOR2_X1 U900 ( .A(n811), .B(n810), .ZN(n905) );
  XNOR2_X1 U901 ( .A(n812), .B(n905), .ZN(n813) );
  NAND2_X1 U902 ( .A1(n813), .A2(G868), .ZN(n817) );
  NAND2_X1 U903 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U904 ( .A1(n817), .A2(n816), .ZN(G295) );
  NAND2_X1 U905 ( .A1(G2084), .A2(G2078), .ZN(n818) );
  XNOR2_X1 U906 ( .A(n818), .B(KEYINPUT85), .ZN(n819) );
  XNOR2_X1 U907 ( .A(KEYINPUT20), .B(n819), .ZN(n820) );
  NAND2_X1 U908 ( .A1(n820), .A2(G2090), .ZN(n821) );
  XNOR2_X1 U909 ( .A(KEYINPUT21), .B(n821), .ZN(n822) );
  NAND2_X1 U910 ( .A1(n822), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U911 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U912 ( .A1(G220), .A2(G219), .ZN(n823) );
  XOR2_X1 U913 ( .A(KEYINPUT22), .B(n823), .Z(n824) );
  NOR2_X1 U914 ( .A1(G218), .A2(n824), .ZN(n825) );
  NAND2_X1 U915 ( .A1(G96), .A2(n825), .ZN(n841) );
  NAND2_X1 U916 ( .A1(G2106), .A2(n841), .ZN(n829) );
  NAND2_X1 U917 ( .A1(G108), .A2(G120), .ZN(n826) );
  NOR2_X1 U918 ( .A1(G237), .A2(n826), .ZN(n827) );
  NAND2_X1 U919 ( .A1(G69), .A2(n827), .ZN(n842) );
  NAND2_X1 U920 ( .A1(G567), .A2(n842), .ZN(n828) );
  NAND2_X1 U921 ( .A1(n829), .A2(n828), .ZN(n830) );
  XOR2_X1 U922 ( .A(KEYINPUT86), .B(n830), .Z(G319) );
  INV_X1 U923 ( .A(G319), .ZN(n833) );
  NAND2_X1 U924 ( .A1(G661), .A2(G483), .ZN(n831) );
  XOR2_X1 U925 ( .A(KEYINPUT87), .B(n831), .Z(n832) );
  NOR2_X1 U926 ( .A1(n833), .A2(n832), .ZN(n840) );
  NAND2_X1 U927 ( .A1(n840), .A2(G36), .ZN(G176) );
  NAND2_X1 U928 ( .A1(G2106), .A2(n834), .ZN(G217) );
  INV_X1 U929 ( .A(G661), .ZN(n836) );
  NAND2_X1 U930 ( .A1(G2), .A2(G15), .ZN(n835) );
  NOR2_X1 U931 ( .A1(n836), .A2(n835), .ZN(n837) );
  XOR2_X1 U932 ( .A(KEYINPUT110), .B(n837), .Z(G259) );
  NAND2_X1 U933 ( .A1(G3), .A2(G1), .ZN(n838) );
  XOR2_X1 U934 ( .A(KEYINPUT111), .B(n838), .Z(n839) );
  NAND2_X1 U935 ( .A1(n840), .A2(n839), .ZN(G188) );
  XOR2_X1 U936 ( .A(G120), .B(KEYINPUT112), .Z(G236) );
  INV_X1 U938 ( .A(G108), .ZN(G238) );
  INV_X1 U939 ( .A(G96), .ZN(G221) );
  NOR2_X1 U940 ( .A1(n842), .A2(n841), .ZN(G325) );
  INV_X1 U941 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U942 ( .A(G1996), .B(KEYINPUT41), .ZN(n852) );
  XOR2_X1 U943 ( .A(G1956), .B(G1961), .Z(n844) );
  XNOR2_X1 U944 ( .A(G1991), .B(G1981), .ZN(n843) );
  XNOR2_X1 U945 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U946 ( .A(G1986), .B(G1966), .Z(n846) );
  XNOR2_X1 U947 ( .A(G1976), .B(G1971), .ZN(n845) );
  XNOR2_X1 U948 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U949 ( .A(n848), .B(n847), .Z(n850) );
  XNOR2_X1 U950 ( .A(KEYINPUT114), .B(G2474), .ZN(n849) );
  XNOR2_X1 U951 ( .A(n850), .B(n849), .ZN(n851) );
  XNOR2_X1 U952 ( .A(n852), .B(n851), .ZN(G229) );
  XOR2_X1 U953 ( .A(G2678), .B(G2084), .Z(n854) );
  XNOR2_X1 U954 ( .A(G2090), .B(G2078), .ZN(n853) );
  XNOR2_X1 U955 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U956 ( .A(n855), .B(G2100), .Z(n857) );
  XNOR2_X1 U957 ( .A(G2067), .B(G2072), .ZN(n856) );
  XNOR2_X1 U958 ( .A(n857), .B(n856), .ZN(n861) );
  XOR2_X1 U959 ( .A(G2096), .B(KEYINPUT113), .Z(n859) );
  XNOR2_X1 U960 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n858) );
  XNOR2_X1 U961 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U962 ( .A(n861), .B(n860), .Z(G227) );
  NAND2_X1 U963 ( .A1(G124), .A2(n714), .ZN(n862) );
  XOR2_X1 U964 ( .A(KEYINPUT115), .B(n862), .Z(n863) );
  XNOR2_X1 U965 ( .A(n863), .B(KEYINPUT44), .ZN(n865) );
  NAND2_X1 U966 ( .A1(G112), .A2(n884), .ZN(n864) );
  NAND2_X1 U967 ( .A1(n865), .A2(n864), .ZN(n869) );
  NAND2_X1 U968 ( .A1(G136), .A2(n887), .ZN(n867) );
  NAND2_X1 U969 ( .A1(G100), .A2(n888), .ZN(n866) );
  NAND2_X1 U970 ( .A1(n867), .A2(n866), .ZN(n868) );
  NOR2_X1 U971 ( .A1(n869), .A2(n868), .ZN(G162) );
  XOR2_X1 U972 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n872) );
  XNOR2_X1 U973 ( .A(n870), .B(KEYINPUT118), .ZN(n871) );
  XNOR2_X1 U974 ( .A(n872), .B(n871), .ZN(n873) );
  XOR2_X1 U975 ( .A(n874), .B(n873), .Z(n900) );
  NAND2_X1 U976 ( .A1(G139), .A2(n887), .ZN(n876) );
  NAND2_X1 U977 ( .A1(G103), .A2(n888), .ZN(n875) );
  NAND2_X1 U978 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U979 ( .A(KEYINPUT117), .B(n877), .Z(n882) );
  NAND2_X1 U980 ( .A1(G115), .A2(n884), .ZN(n879) );
  NAND2_X1 U981 ( .A1(G127), .A2(n714), .ZN(n878) );
  NAND2_X1 U982 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U983 ( .A(KEYINPUT47), .B(n880), .Z(n881) );
  NOR2_X1 U984 ( .A1(n882), .A2(n881), .ZN(n939) );
  XOR2_X1 U985 ( .A(n939), .B(G162), .Z(n883) );
  XNOR2_X1 U986 ( .A(n929), .B(n883), .ZN(n896) );
  NAND2_X1 U987 ( .A1(G118), .A2(n884), .ZN(n886) );
  NAND2_X1 U988 ( .A1(G130), .A2(n714), .ZN(n885) );
  NAND2_X1 U989 ( .A1(n886), .A2(n885), .ZN(n894) );
  NAND2_X1 U990 ( .A1(G142), .A2(n887), .ZN(n890) );
  NAND2_X1 U991 ( .A1(G106), .A2(n888), .ZN(n889) );
  NAND2_X1 U992 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U993 ( .A(KEYINPUT45), .B(n891), .Z(n892) );
  XNOR2_X1 U994 ( .A(KEYINPUT116), .B(n892), .ZN(n893) );
  NOR2_X1 U995 ( .A1(n894), .A2(n893), .ZN(n895) );
  XOR2_X1 U996 ( .A(n896), .B(n895), .Z(n898) );
  XNOR2_X1 U997 ( .A(G164), .B(G160), .ZN(n897) );
  XNOR2_X1 U998 ( .A(n898), .B(n897), .ZN(n899) );
  XNOR2_X1 U999 ( .A(n900), .B(n899), .ZN(n901) );
  XOR2_X1 U1000 ( .A(n902), .B(n901), .Z(n903) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n903), .ZN(n904) );
  XOR2_X1 U1002 ( .A(KEYINPUT119), .B(n904), .Z(G395) );
  XOR2_X1 U1003 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n907) );
  XNOR2_X1 U1004 ( .A(n977), .B(n905), .ZN(n906) );
  XNOR2_X1 U1005 ( .A(n907), .B(n906), .ZN(n909) );
  XOR2_X1 U1006 ( .A(G171), .B(G286), .Z(n908) );
  XNOR2_X1 U1007 ( .A(n909), .B(n908), .ZN(n910) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n910), .ZN(G397) );
  XOR2_X1 U1009 ( .A(G2451), .B(G2430), .Z(n912) );
  XNOR2_X1 U1010 ( .A(G2438), .B(G2443), .ZN(n911) );
  XNOR2_X1 U1011 ( .A(n912), .B(n911), .ZN(n918) );
  XOR2_X1 U1012 ( .A(G2435), .B(G2454), .Z(n914) );
  XNOR2_X1 U1013 ( .A(G1348), .B(G1341), .ZN(n913) );
  XNOR2_X1 U1014 ( .A(n914), .B(n913), .ZN(n916) );
  XOR2_X1 U1015 ( .A(G2446), .B(G2427), .Z(n915) );
  XNOR2_X1 U1016 ( .A(n916), .B(n915), .ZN(n917) );
  XOR2_X1 U1017 ( .A(n918), .B(n917), .Z(n919) );
  NAND2_X1 U1018 ( .A1(G14), .A2(n919), .ZN(n925) );
  NAND2_X1 U1019 ( .A1(n925), .A2(G319), .ZN(n922) );
  NOR2_X1 U1020 ( .A1(G229), .A2(G227), .ZN(n920) );
  XNOR2_X1 U1021 ( .A(KEYINPUT49), .B(n920), .ZN(n921) );
  NOR2_X1 U1022 ( .A1(n922), .A2(n921), .ZN(n924) );
  NOR2_X1 U1023 ( .A1(G395), .A2(G397), .ZN(n923) );
  NAND2_X1 U1024 ( .A1(n924), .A2(n923), .ZN(G225) );
  INV_X1 U1025 ( .A(G225), .ZN(G308) );
  INV_X1 U1026 ( .A(G69), .ZN(G235) );
  INV_X1 U1027 ( .A(n925), .ZN(G401) );
  XOR2_X1 U1028 ( .A(G2090), .B(G162), .Z(n926) );
  NOR2_X1 U1029 ( .A1(n927), .A2(n926), .ZN(n928) );
  XOR2_X1 U1030 ( .A(KEYINPUT51), .B(n928), .Z(n938) );
  XNOR2_X1 U1031 ( .A(G160), .B(G2084), .ZN(n930) );
  NAND2_X1 U1032 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1033 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1034 ( .A1(n934), .A2(n933), .ZN(n935) );
  NOR2_X1 U1035 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1036 ( .A1(n938), .A2(n937), .ZN(n946) );
  XOR2_X1 U1037 ( .A(G2072), .B(n939), .Z(n941) );
  XOR2_X1 U1038 ( .A(G164), .B(G2078), .Z(n940) );
  NOR2_X1 U1039 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1040 ( .A(KEYINPUT50), .B(n942), .ZN(n944) );
  NAND2_X1 U1041 ( .A1(n944), .A2(n943), .ZN(n945) );
  NOR2_X1 U1042 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1043 ( .A(KEYINPUT52), .B(n947), .ZN(n949) );
  INV_X1 U1044 ( .A(KEYINPUT55), .ZN(n948) );
  NAND2_X1 U1045 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1046 ( .A1(n950), .A2(G29), .ZN(n1030) );
  XOR2_X1 U1047 ( .A(G29), .B(KEYINPUT124), .Z(n972) );
  XOR2_X1 U1048 ( .A(G2084), .B(G34), .Z(n951) );
  XNOR2_X1 U1049 ( .A(KEYINPUT54), .B(n951), .ZN(n968) );
  XNOR2_X1 U1050 ( .A(G2090), .B(G35), .ZN(n966) );
  XNOR2_X1 U1051 ( .A(G1991), .B(G25), .ZN(n953) );
  XNOR2_X1 U1052 ( .A(G33), .B(G2072), .ZN(n952) );
  NOR2_X1 U1053 ( .A1(n953), .A2(n952), .ZN(n960) );
  XNOR2_X1 U1054 ( .A(G32), .B(n954), .ZN(n955) );
  NAND2_X1 U1055 ( .A1(n955), .A2(G28), .ZN(n958) );
  XNOR2_X1 U1056 ( .A(KEYINPUT122), .B(G2067), .ZN(n956) );
  XNOR2_X1 U1057 ( .A(G26), .B(n956), .ZN(n957) );
  NOR2_X1 U1058 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1059 ( .A1(n960), .A2(n959), .ZN(n963) );
  XOR2_X1 U1060 ( .A(G27), .B(n961), .Z(n962) );
  NOR2_X1 U1061 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1062 ( .A(KEYINPUT53), .B(n964), .ZN(n965) );
  NOR2_X1 U1063 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1064 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1065 ( .A(n969), .B(KEYINPUT123), .ZN(n970) );
  XNOR2_X1 U1066 ( .A(n970), .B(KEYINPUT55), .ZN(n971) );
  NAND2_X1 U1067 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1068 ( .A1(G11), .A2(n973), .ZN(n1028) );
  XNOR2_X1 U1069 ( .A(G16), .B(KEYINPUT56), .ZN(n998) );
  XOR2_X1 U1070 ( .A(G168), .B(G1966), .Z(n974) );
  NOR2_X1 U1071 ( .A1(n975), .A2(n974), .ZN(n976) );
  XOR2_X1 U1072 ( .A(KEYINPUT57), .B(n976), .Z(n996) );
  XNOR2_X1 U1073 ( .A(G171), .B(G1961), .ZN(n991) );
  XNOR2_X1 U1074 ( .A(G1348), .B(n977), .ZN(n980) );
  XNOR2_X1 U1075 ( .A(n978), .B(G1956), .ZN(n979) );
  NAND2_X1 U1076 ( .A1(n980), .A2(n979), .ZN(n989) );
  NAND2_X1 U1077 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1078 ( .A(n983), .B(KEYINPUT125), .ZN(n987) );
  XNOR2_X1 U1079 ( .A(G1971), .B(G303), .ZN(n984) );
  NOR2_X1 U1080 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1081 ( .A1(n987), .A2(n986), .ZN(n988) );
  NOR2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n994) );
  XNOR2_X1 U1084 ( .A(G1341), .B(n992), .ZN(n993) );
  NOR2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n1026) );
  INV_X1 U1088 ( .A(G16), .ZN(n1024) );
  XOR2_X1 U1089 ( .A(G1986), .B(G24), .Z(n1002) );
  XNOR2_X1 U1090 ( .A(G1976), .B(G23), .ZN(n1000) );
  XNOR2_X1 U1091 ( .A(G1971), .B(G22), .ZN(n999) );
  NOR2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1094 ( .A(KEYINPUT58), .B(n1003), .ZN(n1021) );
  XNOR2_X1 U1095 ( .A(G20), .B(n1004), .ZN(n1008) );
  XNOR2_X1 U1096 ( .A(G1981), .B(G6), .ZN(n1006) );
  XNOR2_X1 U1097 ( .A(G1341), .B(G19), .ZN(n1005) );
  NOR2_X1 U1098 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1099 ( .A1(n1008), .A2(n1007), .ZN(n1011) );
  XOR2_X1 U1100 ( .A(KEYINPUT59), .B(G1348), .Z(n1009) );
  XNOR2_X1 U1101 ( .A(G4), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1102 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1103 ( .A(KEYINPUT126), .B(n1012), .ZN(n1013) );
  XNOR2_X1 U1104 ( .A(n1013), .B(KEYINPUT60), .ZN(n1018) );
  XOR2_X1 U1105 ( .A(n1014), .B(G5), .Z(n1016) );
  XNOR2_X1 U1106 ( .A(G21), .B(G1966), .ZN(n1015) );
  NOR2_X1 U1107 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1108 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1109 ( .A(KEYINPUT127), .B(n1019), .Z(n1020) );
  NOR2_X1 U1110 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1111 ( .A(KEYINPUT61), .B(n1022), .ZN(n1023) );
  NAND2_X1 U1112 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1113 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1114 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1115 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1116 ( .A(KEYINPUT62), .B(n1031), .Z(G311) );
  INV_X1 U1117 ( .A(G311), .ZN(G150) );
endmodule

