

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588;

  XOR2_X1 U322 ( .A(KEYINPUT124), .B(n471), .Z(n584) );
  XNOR2_X1 U323 ( .A(n494), .B(n381), .ZN(n404) );
  INV_X1 U324 ( .A(KEYINPUT27), .ZN(n380) );
  XOR2_X1 U325 ( .A(n377), .B(KEYINPUT93), .Z(n290) );
  AND2_X1 U326 ( .A1(G231GAT), .A2(G233GAT), .ZN(n291) );
  AND2_X1 U327 ( .A1(G226GAT), .A2(G233GAT), .ZN(n292) );
  XNOR2_X1 U328 ( .A(n412), .B(n292), .ZN(n370) );
  XNOR2_X1 U329 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U330 ( .A(n466), .B(KEYINPUT122), .ZN(n467) );
  XOR2_X1 U331 ( .A(G22GAT), .B(G155GAT), .Z(n355) );
  XNOR2_X1 U332 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U333 ( .A(n380), .B(KEYINPUT95), .ZN(n381) );
  XNOR2_X1 U334 ( .A(n332), .B(n291), .ZN(n333) );
  XNOR2_X1 U335 ( .A(n334), .B(n333), .ZN(n338) );
  XNOR2_X1 U336 ( .A(n474), .B(KEYINPUT62), .ZN(n475) );
  XNOR2_X1 U337 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U338 ( .A(n476), .B(n475), .ZN(G1355GAT) );
  XNOR2_X1 U339 ( .A(n453), .B(n452), .ZN(G1330GAT) );
  XNOR2_X1 U340 ( .A(G127GAT), .B(G134GAT), .ZN(n293) );
  XNOR2_X1 U341 ( .A(n293), .B(KEYINPUT0), .ZN(n294) );
  XOR2_X1 U342 ( .A(n294), .B(KEYINPUT80), .Z(n296) );
  XNOR2_X1 U343 ( .A(G113GAT), .B(G120GAT), .ZN(n295) );
  XNOR2_X1 U344 ( .A(n296), .B(n295), .ZN(n392) );
  XOR2_X1 U345 ( .A(KEYINPUT81), .B(KEYINPUT17), .Z(n298) );
  XNOR2_X1 U346 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n297) );
  XNOR2_X1 U347 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U348 ( .A(G169GAT), .B(n299), .Z(n374) );
  XNOR2_X1 U349 ( .A(n392), .B(n374), .ZN(n309) );
  XOR2_X1 U350 ( .A(G176GAT), .B(G183GAT), .Z(n301) );
  XNOR2_X1 U351 ( .A(G43GAT), .B(KEYINPUT20), .ZN(n300) );
  XNOR2_X1 U352 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U353 ( .A(G190GAT), .B(G99GAT), .Z(n303) );
  XNOR2_X1 U354 ( .A(G15GAT), .B(G71GAT), .ZN(n302) );
  XNOR2_X1 U355 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U356 ( .A(n305), .B(n304), .Z(n307) );
  NAND2_X1 U357 ( .A1(G227GAT), .A2(G233GAT), .ZN(n306) );
  XNOR2_X1 U358 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U359 ( .A(n309), .B(n308), .Z(n518) );
  INV_X1 U360 ( .A(n518), .ZN(n560) );
  XOR2_X1 U361 ( .A(KEYINPUT8), .B(KEYINPUT66), .Z(n311) );
  XNOR2_X1 U362 ( .A(G43GAT), .B(G29GAT), .ZN(n310) );
  XNOR2_X1 U363 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U364 ( .A(KEYINPUT7), .B(n312), .Z(n444) );
  XOR2_X1 U365 ( .A(KEYINPUT9), .B(KEYINPUT74), .Z(n314) );
  XNOR2_X1 U366 ( .A(G134GAT), .B(G106GAT), .ZN(n313) );
  XNOR2_X1 U367 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U368 ( .A(n444), .B(n315), .ZN(n327) );
  XOR2_X1 U369 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n317) );
  NAND2_X1 U370 ( .A1(G232GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U371 ( .A(n317), .B(n316), .ZN(n319) );
  XNOR2_X1 U372 ( .A(G36GAT), .B(G190GAT), .ZN(n318) );
  XNOR2_X1 U373 ( .A(n318), .B(KEYINPUT75), .ZN(n378) );
  XOR2_X1 U374 ( .A(n319), .B(n378), .Z(n325) );
  XOR2_X1 U375 ( .A(G162GAT), .B(KEYINPUT73), .Z(n321) );
  XNOR2_X1 U376 ( .A(G50GAT), .B(G218GAT), .ZN(n320) );
  XNOR2_X1 U377 ( .A(n321), .B(n320), .ZN(n359) );
  XOR2_X1 U378 ( .A(G92GAT), .B(KEYINPUT69), .Z(n323) );
  XNOR2_X1 U379 ( .A(G99GAT), .B(G85GAT), .ZN(n322) );
  XNOR2_X1 U380 ( .A(n323), .B(n322), .ZN(n422) );
  XNOR2_X1 U381 ( .A(n359), .B(n422), .ZN(n324) );
  XNOR2_X1 U382 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U383 ( .A(n327), .B(n326), .Z(n555) );
  INV_X1 U384 ( .A(n555), .ZN(n571) );
  XOR2_X1 U385 ( .A(KEYINPUT36), .B(n571), .Z(n472) );
  XOR2_X1 U386 ( .A(n355), .B(G78GAT), .Z(n329) );
  XOR2_X1 U387 ( .A(G15GAT), .B(G1GAT), .Z(n434) );
  XNOR2_X1 U388 ( .A(n434), .B(G127GAT), .ZN(n328) );
  XNOR2_X1 U389 ( .A(n329), .B(n328), .ZN(n334) );
  XOR2_X1 U390 ( .A(KEYINPUT79), .B(KEYINPUT78), .Z(n331) );
  XNOR2_X1 U391 ( .A(G64GAT), .B(KEYINPUT77), .ZN(n330) );
  XNOR2_X1 U392 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U393 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n336) );
  XNOR2_X1 U394 ( .A(G211GAT), .B(KEYINPUT15), .ZN(n335) );
  XNOR2_X1 U395 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U396 ( .A(n338), .B(n337), .Z(n342) );
  XNOR2_X1 U397 ( .A(G71GAT), .B(G57GAT), .ZN(n339) );
  XNOR2_X1 U398 ( .A(n339), .B(KEYINPUT13), .ZN(n413) );
  XNOR2_X1 U399 ( .A(G8GAT), .B(G183GAT), .ZN(n340) );
  XNOR2_X1 U400 ( .A(n340), .B(KEYINPUT76), .ZN(n369) );
  XNOR2_X1 U401 ( .A(n413), .B(n369), .ZN(n341) );
  XOR2_X1 U402 ( .A(n342), .B(n341), .Z(n551) );
  INV_X1 U403 ( .A(n551), .ZN(n585) );
  NOR2_X1 U404 ( .A1(n472), .A2(n585), .ZN(n410) );
  XOR2_X1 U405 ( .A(KEYINPUT87), .B(KEYINPUT2), .Z(n344) );
  XNOR2_X1 U406 ( .A(KEYINPUT3), .B(KEYINPUT88), .ZN(n343) );
  XNOR2_X1 U407 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U408 ( .A(G141GAT), .B(n345), .Z(n391) );
  XOR2_X1 U409 ( .A(G148GAT), .B(G106GAT), .Z(n347) );
  XNOR2_X1 U410 ( .A(G204GAT), .B(G78GAT), .ZN(n346) );
  XNOR2_X1 U411 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U412 ( .A(KEYINPUT68), .B(n348), .ZN(n429) );
  XOR2_X1 U413 ( .A(KEYINPUT86), .B(KEYINPUT85), .Z(n350) );
  XNOR2_X1 U414 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n349) );
  XNOR2_X1 U415 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U416 ( .A(G197GAT), .B(n351), .Z(n373) );
  XOR2_X1 U417 ( .A(n429), .B(n373), .Z(n363) );
  XOR2_X1 U418 ( .A(KEYINPUT82), .B(KEYINPUT84), .Z(n353) );
  XNOR2_X1 U419 ( .A(KEYINPUT22), .B(KEYINPUT83), .ZN(n352) );
  XNOR2_X1 U420 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U421 ( .A(n355), .B(n354), .Z(n357) );
  NAND2_X1 U422 ( .A1(G228GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U423 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U424 ( .A(n358), .B(KEYINPUT24), .Z(n361) );
  XNOR2_X1 U425 ( .A(n359), .B(KEYINPUT23), .ZN(n360) );
  XNOR2_X1 U426 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U427 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U428 ( .A(n391), .B(n364), .ZN(n557) );
  NOR2_X1 U429 ( .A1(n560), .A2(n557), .ZN(n366) );
  XNOR2_X1 U430 ( .A(KEYINPUT26), .B(KEYINPUT98), .ZN(n365) );
  XNOR2_X1 U431 ( .A(n366), .B(n365), .ZN(n470) );
  XOR2_X1 U432 ( .A(KEYINPUT92), .B(G92GAT), .Z(n368) );
  XNOR2_X1 U433 ( .A(G204GAT), .B(G218GAT), .ZN(n367) );
  XNOR2_X1 U434 ( .A(n368), .B(n367), .ZN(n372) );
  XOR2_X1 U435 ( .A(G176GAT), .B(G64GAT), .Z(n412) );
  XOR2_X1 U436 ( .A(n372), .B(n371), .Z(n376) );
  XNOR2_X1 U437 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U438 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U439 ( .A(n378), .B(KEYINPUT94), .ZN(n379) );
  XOR2_X1 U440 ( .A(n290), .B(n379), .Z(n494) );
  NAND2_X1 U441 ( .A1(n470), .A2(n404), .ZN(n540) );
  NAND2_X1 U442 ( .A1(n560), .A2(n494), .ZN(n382) );
  NAND2_X1 U443 ( .A1(n557), .A2(n382), .ZN(n383) );
  XOR2_X1 U444 ( .A(KEYINPUT25), .B(n383), .Z(n384) );
  NAND2_X1 U445 ( .A1(n540), .A2(n384), .ZN(n403) );
  XOR2_X1 U446 ( .A(KEYINPUT6), .B(KEYINPUT91), .Z(n386) );
  XNOR2_X1 U447 ( .A(G1GAT), .B(KEYINPUT90), .ZN(n385) );
  XNOR2_X1 U448 ( .A(n386), .B(n385), .ZN(n390) );
  XOR2_X1 U449 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n388) );
  XNOR2_X1 U450 ( .A(KEYINPUT89), .B(KEYINPUT1), .ZN(n387) );
  XNOR2_X1 U451 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U452 ( .A(n390), .B(n389), .Z(n394) );
  XNOR2_X1 U453 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U454 ( .A(n394), .B(n393), .ZN(n402) );
  NAND2_X1 U455 ( .A1(G225GAT), .A2(G233GAT), .ZN(n400) );
  XOR2_X1 U456 ( .A(G57GAT), .B(G155GAT), .Z(n396) );
  XNOR2_X1 U457 ( .A(G29GAT), .B(G148GAT), .ZN(n395) );
  XNOR2_X1 U458 ( .A(n396), .B(n395), .ZN(n398) );
  XOR2_X1 U459 ( .A(G162GAT), .B(G85GAT), .Z(n397) );
  XNOR2_X1 U460 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U461 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U462 ( .A(n402), .B(n401), .ZN(n514) );
  NAND2_X1 U463 ( .A1(n403), .A2(n514), .ZN(n409) );
  XNOR2_X1 U464 ( .A(KEYINPUT28), .B(n557), .ZN(n521) );
  AND2_X1 U465 ( .A1(n404), .A2(n521), .ZN(n405) );
  INV_X1 U466 ( .A(n514), .ZN(n542) );
  NAND2_X1 U467 ( .A1(n405), .A2(n542), .ZN(n525) );
  XNOR2_X1 U468 ( .A(KEYINPUT96), .B(n525), .ZN(n406) );
  NOR2_X1 U469 ( .A1(n560), .A2(n406), .ZN(n407) );
  XNOR2_X1 U470 ( .A(KEYINPUT97), .B(n407), .ZN(n408) );
  NAND2_X1 U471 ( .A1(n409), .A2(n408), .ZN(n479) );
  NAND2_X1 U472 ( .A1(n410), .A2(n479), .ZN(n411) );
  XNOR2_X1 U473 ( .A(n411), .B(KEYINPUT37), .ZN(n513) );
  XNOR2_X1 U474 ( .A(n413), .B(n412), .ZN(n417) );
  INV_X1 U475 ( .A(n417), .ZN(n415) );
  AND2_X1 U476 ( .A1(G230GAT), .A2(G233GAT), .ZN(n416) );
  INV_X1 U477 ( .A(n416), .ZN(n414) );
  NAND2_X1 U478 ( .A1(n415), .A2(n414), .ZN(n419) );
  NAND2_X1 U479 ( .A1(n417), .A2(n416), .ZN(n418) );
  NAND2_X1 U480 ( .A1(n419), .A2(n418), .ZN(n421) );
  INV_X1 U481 ( .A(KEYINPUT70), .ZN(n420) );
  XNOR2_X1 U482 ( .A(n421), .B(n420), .ZN(n424) );
  XNOR2_X1 U483 ( .A(n422), .B(KEYINPUT71), .ZN(n423) );
  XNOR2_X1 U484 ( .A(n424), .B(n423), .ZN(n428) );
  XOR2_X1 U485 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n426) );
  XNOR2_X1 U486 ( .A(G120GAT), .B(KEYINPUT33), .ZN(n425) );
  XNOR2_X1 U487 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U488 ( .A(n428), .B(n427), .ZN(n430) );
  XNOR2_X1 U489 ( .A(n430), .B(n429), .ZN(n580) );
  XOR2_X1 U490 ( .A(G113GAT), .B(G36GAT), .Z(n432) );
  XNOR2_X1 U491 ( .A(G169GAT), .B(G50GAT), .ZN(n431) );
  XNOR2_X1 U492 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U493 ( .A(n434), .B(n433), .Z(n436) );
  NAND2_X1 U494 ( .A1(G229GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U495 ( .A(n436), .B(n435), .ZN(n440) );
  XOR2_X1 U496 ( .A(KEYINPUT30), .B(KEYINPUT65), .Z(n438) );
  XNOR2_X1 U497 ( .A(KEYINPUT29), .B(KEYINPUT67), .ZN(n437) );
  XNOR2_X1 U498 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U499 ( .A(n440), .B(n439), .Z(n446) );
  XOR2_X1 U500 ( .A(G8GAT), .B(G141GAT), .Z(n442) );
  XNOR2_X1 U501 ( .A(G197GAT), .B(G22GAT), .ZN(n441) );
  XNOR2_X1 U502 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U503 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U504 ( .A(n446), .B(n445), .Z(n576) );
  INV_X1 U505 ( .A(n576), .ZN(n562) );
  NOR2_X1 U506 ( .A1(n580), .A2(n562), .ZN(n447) );
  XNOR2_X1 U507 ( .A(n447), .B(KEYINPUT72), .ZN(n480) );
  NAND2_X1 U508 ( .A1(n513), .A2(n480), .ZN(n448) );
  XNOR2_X1 U509 ( .A(n448), .B(KEYINPUT38), .ZN(n449) );
  XNOR2_X1 U510 ( .A(KEYINPUT103), .B(n449), .ZN(n498) );
  NAND2_X1 U511 ( .A1(n560), .A2(n498), .ZN(n453) );
  XOR2_X1 U512 ( .A(KEYINPUT40), .B(KEYINPUT106), .Z(n451) );
  XNOR2_X1 U513 ( .A(G43GAT), .B(KEYINPUT105), .ZN(n450) );
  INV_X1 U514 ( .A(n494), .ZN(n516) );
  XNOR2_X1 U515 ( .A(KEYINPUT41), .B(n580), .ZN(n564) );
  NOR2_X1 U516 ( .A1(n562), .A2(n564), .ZN(n454) );
  XNOR2_X1 U517 ( .A(n454), .B(KEYINPUT46), .ZN(n455) );
  XOR2_X1 U518 ( .A(n551), .B(KEYINPUT112), .Z(n569) );
  NOR2_X1 U519 ( .A1(n455), .A2(n569), .ZN(n456) );
  XNOR2_X1 U520 ( .A(n456), .B(KEYINPUT113), .ZN(n457) );
  NOR2_X1 U521 ( .A1(n457), .A2(n571), .ZN(n458) );
  XNOR2_X1 U522 ( .A(n458), .B(KEYINPUT47), .ZN(n463) );
  NOR2_X1 U523 ( .A1(n472), .A2(n551), .ZN(n459) );
  XOR2_X1 U524 ( .A(KEYINPUT45), .B(n459), .Z(n460) );
  NOR2_X1 U525 ( .A1(n580), .A2(n460), .ZN(n461) );
  NAND2_X1 U526 ( .A1(n461), .A2(n562), .ZN(n462) );
  AND2_X1 U527 ( .A1(n463), .A2(n462), .ZN(n465) );
  XNOR2_X1 U528 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n464) );
  XNOR2_X1 U529 ( .A(n465), .B(n464), .ZN(n541) );
  NOR2_X1 U530 ( .A1(n516), .A2(n541), .ZN(n468) );
  INV_X1 U531 ( .A(KEYINPUT54), .ZN(n466) );
  NOR2_X1 U532 ( .A1(n469), .A2(n542), .ZN(n558) );
  NAND2_X1 U533 ( .A1(n470), .A2(n558), .ZN(n471) );
  INV_X1 U534 ( .A(n584), .ZN(n473) );
  NOR2_X1 U535 ( .A1(n473), .A2(n472), .ZN(n476) );
  INV_X1 U536 ( .A(G218GAT), .ZN(n474) );
  NAND2_X1 U537 ( .A1(n585), .A2(n555), .ZN(n477) );
  XOR2_X1 U538 ( .A(KEYINPUT16), .B(n477), .Z(n478) );
  AND2_X1 U539 ( .A1(n479), .A2(n478), .ZN(n501) );
  NAND2_X1 U540 ( .A1(n501), .A2(n480), .ZN(n489) );
  NOR2_X1 U541 ( .A1(n514), .A2(n489), .ZN(n481) );
  XOR2_X1 U542 ( .A(KEYINPUT34), .B(n481), .Z(n482) );
  XNOR2_X1 U543 ( .A(G1GAT), .B(n482), .ZN(G1324GAT) );
  NOR2_X1 U544 ( .A1(n516), .A2(n489), .ZN(n483) );
  XOR2_X1 U545 ( .A(G8GAT), .B(n483), .Z(G1325GAT) );
  XOR2_X1 U546 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n485) );
  XNOR2_X1 U547 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n484) );
  XNOR2_X1 U548 ( .A(n485), .B(n484), .ZN(n487) );
  NOR2_X1 U549 ( .A1(n518), .A2(n489), .ZN(n486) );
  XOR2_X1 U550 ( .A(n487), .B(n486), .Z(n488) );
  XNOR2_X1 U551 ( .A(KEYINPUT99), .B(n488), .ZN(G1326GAT) );
  NOR2_X1 U552 ( .A1(n521), .A2(n489), .ZN(n490) );
  XOR2_X1 U553 ( .A(KEYINPUT102), .B(n490), .Z(n491) );
  XNOR2_X1 U554 ( .A(G22GAT), .B(n491), .ZN(G1327GAT) );
  XOR2_X1 U555 ( .A(G29GAT), .B(KEYINPUT39), .Z(n493) );
  NAND2_X1 U556 ( .A1(n498), .A2(n542), .ZN(n492) );
  XNOR2_X1 U557 ( .A(n493), .B(n492), .ZN(G1328GAT) );
  NAND2_X1 U558 ( .A1(n498), .A2(n494), .ZN(n495) );
  XNOR2_X1 U559 ( .A(n495), .B(KEYINPUT104), .ZN(n496) );
  XNOR2_X1 U560 ( .A(G36GAT), .B(n496), .ZN(G1329GAT) );
  INV_X1 U561 ( .A(n521), .ZN(n497) );
  NAND2_X1 U562 ( .A1(n498), .A2(n497), .ZN(n499) );
  XNOR2_X1 U563 ( .A(n499), .B(G50GAT), .ZN(G1331GAT) );
  NOR2_X1 U564 ( .A1(n576), .A2(n564), .ZN(n500) );
  XNOR2_X1 U565 ( .A(n500), .B(KEYINPUT108), .ZN(n512) );
  NAND2_X1 U566 ( .A1(n501), .A2(n512), .ZN(n508) );
  NOR2_X1 U567 ( .A1(n508), .A2(n514), .ZN(n505) );
  XOR2_X1 U568 ( .A(KEYINPUT107), .B(KEYINPUT42), .Z(n503) );
  XNOR2_X1 U569 ( .A(G57GAT), .B(KEYINPUT109), .ZN(n502) );
  XNOR2_X1 U570 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U571 ( .A(n505), .B(n504), .ZN(G1332GAT) );
  NOR2_X1 U572 ( .A1(n516), .A2(n508), .ZN(n506) );
  XOR2_X1 U573 ( .A(G64GAT), .B(n506), .Z(G1333GAT) );
  NOR2_X1 U574 ( .A1(n518), .A2(n508), .ZN(n507) );
  XOR2_X1 U575 ( .A(G71GAT), .B(n507), .Z(G1334GAT) );
  NOR2_X1 U576 ( .A1(n521), .A2(n508), .ZN(n510) );
  XNOR2_X1 U577 ( .A(KEYINPUT110), .B(KEYINPUT43), .ZN(n509) );
  XNOR2_X1 U578 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U579 ( .A(G78GAT), .B(n511), .ZN(G1335GAT) );
  NAND2_X1 U580 ( .A1(n513), .A2(n512), .ZN(n520) );
  NOR2_X1 U581 ( .A1(n514), .A2(n520), .ZN(n515) );
  XOR2_X1 U582 ( .A(G85GAT), .B(n515), .Z(G1336GAT) );
  NOR2_X1 U583 ( .A1(n516), .A2(n520), .ZN(n517) );
  XOR2_X1 U584 ( .A(G92GAT), .B(n517), .Z(G1337GAT) );
  NOR2_X1 U585 ( .A1(n518), .A2(n520), .ZN(n519) );
  XOR2_X1 U586 ( .A(G99GAT), .B(n519), .Z(G1338GAT) );
  NOR2_X1 U587 ( .A1(n521), .A2(n520), .ZN(n523) );
  XNOR2_X1 U588 ( .A(KEYINPUT44), .B(KEYINPUT111), .ZN(n522) );
  XNOR2_X1 U589 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U590 ( .A(G106GAT), .B(n524), .ZN(G1339GAT) );
  NOR2_X1 U591 ( .A1(n541), .A2(n525), .ZN(n526) );
  NAND2_X1 U592 ( .A1(n526), .A2(n560), .ZN(n527) );
  XOR2_X1 U593 ( .A(n527), .B(KEYINPUT114), .Z(n537) );
  INV_X1 U594 ( .A(n537), .ZN(n529) );
  NOR2_X1 U595 ( .A1(n562), .A2(n529), .ZN(n528) );
  XOR2_X1 U596 ( .A(G113GAT), .B(n528), .Z(G1340GAT) );
  NOR2_X1 U597 ( .A1(n529), .A2(n564), .ZN(n533) );
  XOR2_X1 U598 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n531) );
  XNOR2_X1 U599 ( .A(G120GAT), .B(KEYINPUT116), .ZN(n530) );
  XNOR2_X1 U600 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U601 ( .A(n533), .B(n532), .ZN(G1341GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n535) );
  NAND2_X1 U603 ( .A1(n537), .A2(n569), .ZN(n534) );
  XNOR2_X1 U604 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U605 ( .A(G127GAT), .B(n536), .ZN(G1342GAT) );
  XOR2_X1 U606 ( .A(G134GAT), .B(KEYINPUT51), .Z(n539) );
  NAND2_X1 U607 ( .A1(n571), .A2(n537), .ZN(n538) );
  XNOR2_X1 U608 ( .A(n539), .B(n538), .ZN(G1343GAT) );
  NOR2_X1 U609 ( .A1(n541), .A2(n540), .ZN(n543) );
  NAND2_X1 U610 ( .A1(n543), .A2(n542), .ZN(n554) );
  NOR2_X1 U611 ( .A1(n562), .A2(n554), .ZN(n544) );
  XOR2_X1 U612 ( .A(KEYINPUT118), .B(n544), .Z(n545) );
  XNOR2_X1 U613 ( .A(G141GAT), .B(n545), .ZN(G1344GAT) );
  NOR2_X1 U614 ( .A1(n564), .A2(n554), .ZN(n550) );
  XOR2_X1 U615 ( .A(KEYINPUT53), .B(KEYINPUT120), .Z(n547) );
  XNOR2_X1 U616 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n546) );
  XNOR2_X1 U617 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U618 ( .A(KEYINPUT119), .B(n548), .ZN(n549) );
  XNOR2_X1 U619 ( .A(n550), .B(n549), .ZN(G1345GAT) );
  NOR2_X1 U620 ( .A1(n551), .A2(n554), .ZN(n553) );
  XNOR2_X1 U621 ( .A(G155GAT), .B(KEYINPUT121), .ZN(n552) );
  XNOR2_X1 U622 ( .A(n553), .B(n552), .ZN(G1346GAT) );
  NOR2_X1 U623 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U624 ( .A(G162GAT), .B(n556), .Z(G1347GAT) );
  NAND2_X1 U625 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n559), .B(KEYINPUT55), .ZN(n561) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n568) );
  NOR2_X1 U628 ( .A1(n568), .A2(n562), .ZN(n563) );
  XOR2_X1 U629 ( .A(G169GAT), .B(n563), .Z(G1348GAT) );
  NOR2_X1 U630 ( .A1(n564), .A2(n568), .ZN(n566) );
  XNOR2_X1 U631 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n567), .B(G176GAT), .ZN(G1349GAT) );
  INV_X1 U634 ( .A(n568), .ZN(n572) );
  NAND2_X1 U635 ( .A1(n569), .A2(n572), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n570), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n574) );
  NAND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(G190GAT), .ZN(G1351GAT) );
  XNOR2_X1 U641 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n578) );
  AND2_X1 U642 ( .A1(n576), .A2(n584), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n579), .B(G197GAT), .ZN(G1352GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n582) );
  NAND2_X1 U646 ( .A1(n584), .A2(n580), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(n583) );
  XOR2_X1 U648 ( .A(G204GAT), .B(n583), .Z(G1353GAT) );
  XOR2_X1 U649 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n587) );
  NAND2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U652 ( .A(G211GAT), .B(n588), .ZN(G1354GAT) );
endmodule

