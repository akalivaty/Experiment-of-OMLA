

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588;

  XNOR2_X1 U322 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U323 ( .A(n446), .B(n445), .ZN(n447) );
  INV_X1 U324 ( .A(G113GAT), .ZN(n352) );
  XNOR2_X1 U325 ( .A(n353), .B(n352), .ZN(n354) );
  INV_X1 U326 ( .A(KEYINPUT54), .ZN(n469) );
  XNOR2_X1 U327 ( .A(n465), .B(KEYINPUT48), .ZN(n466) );
  XNOR2_X1 U328 ( .A(n469), .B(KEYINPUT119), .ZN(n470) );
  XNOR2_X1 U329 ( .A(n467), .B(n466), .ZN(n534) );
  NOR2_X1 U330 ( .A1(n409), .A2(n408), .ZN(n490) );
  XNOR2_X1 U331 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U332 ( .A(KEYINPUT37), .B(KEYINPUT104), .ZN(n411) );
  XNOR2_X1 U333 ( .A(n448), .B(n447), .ZN(n453) );
  XNOR2_X1 U334 ( .A(n412), .B(n411), .ZN(n523) );
  XNOR2_X1 U335 ( .A(n364), .B(n378), .ZN(n535) );
  XNOR2_X1 U336 ( .A(n476), .B(G190GAT), .ZN(n477) );
  XNOR2_X1 U337 ( .A(n450), .B(G43GAT), .ZN(n451) );
  XNOR2_X1 U338 ( .A(n478), .B(n477), .ZN(G1351GAT) );
  XNOR2_X1 U339 ( .A(n452), .B(n451), .ZN(G1330GAT) );
  XOR2_X1 U340 ( .A(KEYINPUT15), .B(G64GAT), .Z(n291) );
  XNOR2_X1 U341 ( .A(G183GAT), .B(G71GAT), .ZN(n290) );
  XNOR2_X1 U342 ( .A(n291), .B(n290), .ZN(n295) );
  XOR2_X1 U343 ( .A(KEYINPUT80), .B(KEYINPUT12), .Z(n293) );
  XNOR2_X1 U344 ( .A(G1GAT), .B(KEYINPUT14), .ZN(n292) );
  XNOR2_X1 U345 ( .A(n293), .B(n292), .ZN(n294) );
  XNOR2_X1 U346 ( .A(n295), .B(n294), .ZN(n305) );
  XOR2_X1 U347 ( .A(G15GAT), .B(G127GAT), .Z(n348) );
  XNOR2_X1 U348 ( .A(G57GAT), .B(KEYINPUT72), .ZN(n296) );
  XNOR2_X1 U349 ( .A(n296), .B(KEYINPUT13), .ZN(n441) );
  XOR2_X1 U350 ( .A(n441), .B(KEYINPUT79), .Z(n298) );
  NAND2_X1 U351 ( .A1(G231GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U352 ( .A(n298), .B(n297), .ZN(n299) );
  XNOR2_X1 U353 ( .A(n348), .B(n299), .ZN(n303) );
  XOR2_X1 U354 ( .A(G8GAT), .B(KEYINPUT78), .Z(n365) );
  XOR2_X1 U355 ( .A(G22GAT), .B(G155GAT), .Z(n382) );
  XOR2_X1 U356 ( .A(n365), .B(n382), .Z(n301) );
  XNOR2_X1 U357 ( .A(G211GAT), .B(G78GAT), .ZN(n300) );
  XNOR2_X1 U358 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U359 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U360 ( .A(n305), .B(n304), .Z(n557) );
  INV_X1 U361 ( .A(n557), .ZN(n581) );
  XOR2_X1 U362 ( .A(KEYINPUT67), .B(KEYINPUT75), .Z(n307) );
  XNOR2_X1 U363 ( .A(G92GAT), .B(KEYINPUT10), .ZN(n306) );
  XNOR2_X1 U364 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U365 ( .A(G50GAT), .B(G162GAT), .Z(n381) );
  XOR2_X1 U366 ( .A(n308), .B(n381), .Z(n310) );
  XNOR2_X1 U367 ( .A(G218GAT), .B(G106GAT), .ZN(n309) );
  XNOR2_X1 U368 ( .A(n310), .B(n309), .ZN(n315) );
  XNOR2_X1 U369 ( .A(G36GAT), .B(G190GAT), .ZN(n311) );
  XNOR2_X1 U370 ( .A(n311), .B(KEYINPUT77), .ZN(n368) );
  XNOR2_X1 U371 ( .A(G99GAT), .B(G85GAT), .ZN(n445) );
  XNOR2_X1 U372 ( .A(n368), .B(n445), .ZN(n313) );
  NAND2_X1 U373 ( .A1(G232GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U374 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U375 ( .A(n315), .B(n314), .Z(n323) );
  XOR2_X1 U376 ( .A(KEYINPUT71), .B(KEYINPUT7), .Z(n317) );
  XNOR2_X1 U377 ( .A(G43GAT), .B(G29GAT), .ZN(n316) );
  XNOR2_X1 U378 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U379 ( .A(KEYINPUT8), .B(n318), .Z(n426) );
  XOR2_X1 U380 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n320) );
  XNOR2_X1 U381 ( .A(G134GAT), .B(KEYINPUT76), .ZN(n319) );
  XNOR2_X1 U382 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U383 ( .A(n426), .B(n321), .ZN(n322) );
  XOR2_X1 U384 ( .A(n323), .B(n322), .Z(n561) );
  XOR2_X1 U385 ( .A(KEYINPUT36), .B(n561), .Z(n586) );
  XOR2_X1 U386 ( .A(KEYINPUT90), .B(KEYINPUT1), .Z(n325) );
  XNOR2_X1 U387 ( .A(G120GAT), .B(G57GAT), .ZN(n324) );
  XNOR2_X1 U388 ( .A(n325), .B(n324), .ZN(n329) );
  XOR2_X1 U389 ( .A(KEYINPUT6), .B(KEYINPUT93), .Z(n327) );
  XNOR2_X1 U390 ( .A(KEYINPUT91), .B(KEYINPUT92), .ZN(n326) );
  XNOR2_X1 U391 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U392 ( .A(n329), .B(n328), .Z(n334) );
  XOR2_X1 U393 ( .A(KEYINPUT89), .B(KEYINPUT4), .Z(n331) );
  NAND2_X1 U394 ( .A1(G225GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U395 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U396 ( .A(KEYINPUT5), .B(n332), .ZN(n333) );
  XNOR2_X1 U397 ( .A(n334), .B(n333), .ZN(n341) );
  XOR2_X1 U398 ( .A(G85GAT), .B(G155GAT), .Z(n336) );
  XNOR2_X1 U399 ( .A(G127GAT), .B(G162GAT), .ZN(n335) );
  XNOR2_X1 U400 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U401 ( .A(n337), .B(G148GAT), .Z(n339) );
  XOR2_X1 U402 ( .A(G113GAT), .B(G1GAT), .Z(n416) );
  XNOR2_X1 U403 ( .A(G29GAT), .B(n416), .ZN(n338) );
  XNOR2_X1 U404 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U405 ( .A(n341), .B(n340), .Z(n345) );
  XNOR2_X1 U406 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n342) );
  XNOR2_X1 U407 ( .A(n342), .B(KEYINPUT83), .ZN(n355) );
  XNOR2_X1 U408 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n343) );
  XNOR2_X1 U409 ( .A(n343), .B(KEYINPUT2), .ZN(n380) );
  XNOR2_X1 U410 ( .A(n355), .B(n380), .ZN(n344) );
  XNOR2_X1 U411 ( .A(n345), .B(n344), .ZN(n548) );
  XOR2_X1 U412 ( .A(KEYINPUT66), .B(KEYINPUT20), .Z(n347) );
  XNOR2_X1 U413 ( .A(G176GAT), .B(KEYINPUT85), .ZN(n346) );
  XNOR2_X1 U414 ( .A(n347), .B(n346), .ZN(n360) );
  XOR2_X1 U415 ( .A(G99GAT), .B(G190GAT), .Z(n350) );
  XOR2_X1 U416 ( .A(G120GAT), .B(G71GAT), .Z(n446) );
  XNOR2_X1 U417 ( .A(n348), .B(n446), .ZN(n349) );
  XNOR2_X1 U418 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U419 ( .A(n351), .B(KEYINPUT84), .Z(n358) );
  NAND2_X1 U420 ( .A1(G227GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U421 ( .A(G43GAT), .B(n356), .ZN(n357) );
  XNOR2_X1 U422 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U423 ( .A(n360), .B(n359), .ZN(n364) );
  XOR2_X1 U424 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n362) );
  XNOR2_X1 U425 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n361) );
  XNOR2_X1 U426 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U427 ( .A(G169GAT), .B(n363), .ZN(n378) );
  XOR2_X1 U428 ( .A(KEYINPUT94), .B(n365), .Z(n367) );
  NAND2_X1 U429 ( .A1(G226GAT), .A2(G233GAT), .ZN(n366) );
  XNOR2_X1 U430 ( .A(n367), .B(n366), .ZN(n369) );
  XOR2_X1 U431 ( .A(n369), .B(n368), .Z(n377) );
  XNOR2_X1 U432 ( .A(G211GAT), .B(KEYINPUT88), .ZN(n370) );
  XNOR2_X1 U433 ( .A(n370), .B(KEYINPUT21), .ZN(n371) );
  XOR2_X1 U434 ( .A(n371), .B(KEYINPUT87), .Z(n373) );
  XNOR2_X1 U435 ( .A(G197GAT), .B(G218GAT), .ZN(n372) );
  XNOR2_X1 U436 ( .A(n373), .B(n372), .ZN(n392) );
  XOR2_X1 U437 ( .A(G64GAT), .B(G92GAT), .Z(n375) );
  XNOR2_X1 U438 ( .A(G176GAT), .B(G204GAT), .ZN(n374) );
  XNOR2_X1 U439 ( .A(n375), .B(n374), .ZN(n442) );
  XNOR2_X1 U440 ( .A(n392), .B(n442), .ZN(n376) );
  XNOR2_X1 U441 ( .A(n377), .B(n376), .ZN(n379) );
  XNOR2_X1 U442 ( .A(n379), .B(n378), .ZN(n526) );
  NAND2_X1 U443 ( .A1(n535), .A2(n526), .ZN(n395) );
  XNOR2_X1 U444 ( .A(n381), .B(n380), .ZN(n383) );
  XNOR2_X1 U445 ( .A(n383), .B(n382), .ZN(n388) );
  XNOR2_X1 U446 ( .A(G106GAT), .B(G78GAT), .ZN(n384) );
  XNOR2_X1 U447 ( .A(n384), .B(G148GAT), .ZN(n431) );
  XOR2_X1 U448 ( .A(n431), .B(KEYINPUT86), .Z(n386) );
  NAND2_X1 U449 ( .A1(G228GAT), .A2(G233GAT), .ZN(n385) );
  XNOR2_X1 U450 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U451 ( .A(n388), .B(n387), .Z(n394) );
  XOR2_X1 U452 ( .A(KEYINPUT23), .B(G204GAT), .Z(n390) );
  XNOR2_X1 U453 ( .A(KEYINPUT24), .B(KEYINPUT22), .ZN(n389) );
  XNOR2_X1 U454 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U455 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U456 ( .A(n394), .B(n393), .ZN(n473) );
  NAND2_X1 U457 ( .A1(n395), .A2(n473), .ZN(n396) );
  XNOR2_X1 U458 ( .A(n396), .B(KEYINPUT98), .ZN(n398) );
  XOR2_X1 U459 ( .A(KEYINPUT97), .B(KEYINPUT25), .Z(n397) );
  XNOR2_X1 U460 ( .A(n398), .B(n397), .ZN(n402) );
  NOR2_X1 U461 ( .A1(n473), .A2(n535), .ZN(n399) );
  XOR2_X1 U462 ( .A(KEYINPUT26), .B(n399), .Z(n400) );
  XNOR2_X1 U463 ( .A(KEYINPUT95), .B(n400), .ZN(n569) );
  XNOR2_X1 U464 ( .A(n526), .B(KEYINPUT27), .ZN(n404) );
  NAND2_X1 U465 ( .A1(n569), .A2(n404), .ZN(n550) );
  XOR2_X1 U466 ( .A(KEYINPUT96), .B(n550), .Z(n401) );
  NOR2_X1 U467 ( .A1(n402), .A2(n401), .ZN(n403) );
  NOR2_X1 U468 ( .A1(n548), .A2(n403), .ZN(n409) );
  INV_X1 U469 ( .A(n404), .ZN(n406) );
  XOR2_X1 U470 ( .A(n473), .B(KEYINPUT68), .Z(n405) );
  XNOR2_X1 U471 ( .A(KEYINPUT28), .B(n405), .ZN(n529) );
  NOR2_X1 U472 ( .A1(n406), .A2(n529), .ZN(n407) );
  NAND2_X1 U473 ( .A1(n548), .A2(n407), .ZN(n537) );
  NOR2_X1 U474 ( .A1(n537), .A2(n535), .ZN(n408) );
  NOR2_X1 U475 ( .A1(n586), .A2(n490), .ZN(n410) );
  NAND2_X1 U476 ( .A1(n581), .A2(n410), .ZN(n412) );
  XOR2_X1 U477 ( .A(G22GAT), .B(G141GAT), .Z(n414) );
  XNOR2_X1 U478 ( .A(G36GAT), .B(G50GAT), .ZN(n413) );
  XNOR2_X1 U479 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U480 ( .A(n416), .B(n415), .Z(n418) );
  NAND2_X1 U481 ( .A1(G229GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U482 ( .A(n418), .B(n417), .ZN(n422) );
  XOR2_X1 U483 ( .A(KEYINPUT30), .B(KEYINPUT69), .Z(n420) );
  XNOR2_X1 U484 ( .A(KEYINPUT29), .B(KEYINPUT70), .ZN(n419) );
  XNOR2_X1 U485 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U486 ( .A(n422), .B(n421), .Z(n428) );
  XOR2_X1 U487 ( .A(G8GAT), .B(G15GAT), .Z(n424) );
  XNOR2_X1 U488 ( .A(G169GAT), .B(G197GAT), .ZN(n423) );
  XNOR2_X1 U489 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U490 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U491 ( .A(n428), .B(n427), .Z(n551) );
  INV_X1 U492 ( .A(n551), .ZN(n571) );
  XNOR2_X1 U493 ( .A(n431), .B(KEYINPUT33), .ZN(n429) );
  AND2_X1 U494 ( .A1(G230GAT), .A2(G233GAT), .ZN(n432) );
  NAND2_X1 U495 ( .A1(n429), .A2(n432), .ZN(n436) );
  INV_X1 U496 ( .A(KEYINPUT33), .ZN(n430) );
  XNOR2_X1 U497 ( .A(n431), .B(n430), .ZN(n434) );
  INV_X1 U498 ( .A(n432), .ZN(n433) );
  NAND2_X1 U499 ( .A1(n434), .A2(n433), .ZN(n435) );
  NAND2_X1 U500 ( .A1(n436), .A2(n435), .ZN(n440) );
  XOR2_X1 U501 ( .A(KEYINPUT32), .B(KEYINPUT74), .Z(n438) );
  XNOR2_X1 U502 ( .A(KEYINPUT73), .B(KEYINPUT31), .ZN(n437) );
  XNOR2_X1 U503 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U504 ( .A(n440), .B(n439), .ZN(n444) );
  XOR2_X1 U505 ( .A(n442), .B(n441), .Z(n443) );
  XNOR2_X1 U506 ( .A(n444), .B(n443), .ZN(n448) );
  NOR2_X1 U507 ( .A1(n571), .A2(n453), .ZN(n491) );
  NAND2_X1 U508 ( .A1(n523), .A2(n491), .ZN(n449) );
  XOR2_X1 U509 ( .A(KEYINPUT38), .B(n449), .Z(n507) );
  NAND2_X1 U510 ( .A1(n507), .A2(n535), .ZN(n452) );
  XOR2_X1 U511 ( .A(KEYINPUT40), .B(KEYINPUT105), .Z(n450) );
  INV_X1 U512 ( .A(n561), .ZN(n485) );
  XNOR2_X1 U513 ( .A(KEYINPUT118), .B(n526), .ZN(n468) );
  XNOR2_X1 U514 ( .A(KEYINPUT41), .B(KEYINPUT65), .ZN(n454) );
  XOR2_X1 U515 ( .A(n454), .B(n453), .Z(n564) );
  INV_X1 U516 ( .A(n564), .ZN(n539) );
  NAND2_X1 U517 ( .A1(n551), .A2(n539), .ZN(n455) );
  XNOR2_X1 U518 ( .A(n455), .B(KEYINPUT46), .ZN(n456) );
  NAND2_X1 U519 ( .A1(n456), .A2(n581), .ZN(n457) );
  XNOR2_X1 U520 ( .A(n457), .B(KEYINPUT113), .ZN(n458) );
  NAND2_X1 U521 ( .A1(n458), .A2(n485), .ZN(n459) );
  XNOR2_X1 U522 ( .A(n459), .B(KEYINPUT47), .ZN(n464) );
  NOR2_X1 U523 ( .A1(n581), .A2(n586), .ZN(n460) );
  XNOR2_X1 U524 ( .A(KEYINPUT45), .B(n460), .ZN(n461) );
  NAND2_X1 U525 ( .A1(n461), .A2(n571), .ZN(n462) );
  NOR2_X1 U526 ( .A1(n453), .A2(n462), .ZN(n463) );
  NOR2_X1 U527 ( .A1(n464), .A2(n463), .ZN(n467) );
  XOR2_X1 U528 ( .A(KEYINPUT64), .B(KEYINPUT114), .Z(n465) );
  NAND2_X1 U529 ( .A1(n468), .A2(n534), .ZN(n471) );
  NOR2_X1 U530 ( .A1(n548), .A2(n472), .ZN(n570) );
  NAND2_X1 U531 ( .A1(n473), .A2(n570), .ZN(n474) );
  XNOR2_X1 U532 ( .A(n474), .B(KEYINPUT55), .ZN(n475) );
  NAND2_X1 U533 ( .A1(n475), .A2(n535), .ZN(n563) );
  NOR2_X1 U534 ( .A1(n485), .A2(n563), .ZN(n478) );
  INV_X1 U535 ( .A(KEYINPUT58), .ZN(n476) );
  NOR2_X1 U536 ( .A1(n581), .A2(n563), .ZN(n481) );
  INV_X1 U537 ( .A(G183GAT), .ZN(n479) );
  XNOR2_X1 U538 ( .A(n479), .B(KEYINPUT122), .ZN(n480) );
  XNOR2_X1 U539 ( .A(n481), .B(n480), .ZN(G1350GAT) );
  INV_X1 U540 ( .A(G169GAT), .ZN(n484) );
  NOR2_X1 U541 ( .A1(n571), .A2(n563), .ZN(n482) );
  XNOR2_X1 U542 ( .A(n482), .B(KEYINPUT120), .ZN(n483) );
  XNOR2_X1 U543 ( .A(n484), .B(n483), .ZN(G1348GAT) );
  XOR2_X1 U544 ( .A(KEYINPUT16), .B(KEYINPUT82), .Z(n487) );
  NAND2_X1 U545 ( .A1(n485), .A2(n557), .ZN(n486) );
  XNOR2_X1 U546 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U547 ( .A(n488), .B(KEYINPUT81), .ZN(n489) );
  NOR2_X1 U548 ( .A1(n490), .A2(n489), .ZN(n511) );
  NAND2_X1 U549 ( .A1(n491), .A2(n511), .ZN(n492) );
  XNOR2_X1 U550 ( .A(KEYINPUT99), .B(n492), .ZN(n501) );
  NAND2_X1 U551 ( .A1(n501), .A2(n548), .ZN(n496) );
  XOR2_X1 U552 ( .A(KEYINPUT34), .B(KEYINPUT101), .Z(n494) );
  XNOR2_X1 U553 ( .A(G1GAT), .B(KEYINPUT100), .ZN(n493) );
  XNOR2_X1 U554 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U555 ( .A(n496), .B(n495), .ZN(G1324GAT) );
  NAND2_X1 U556 ( .A1(n501), .A2(n526), .ZN(n497) );
  XNOR2_X1 U557 ( .A(n497), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U558 ( .A(KEYINPUT102), .B(KEYINPUT35), .Z(n499) );
  NAND2_X1 U559 ( .A1(n501), .A2(n535), .ZN(n498) );
  XNOR2_X1 U560 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U561 ( .A(G15GAT), .B(n500), .ZN(G1326GAT) );
  XOR2_X1 U562 ( .A(G22GAT), .B(KEYINPUT103), .Z(n503) );
  NAND2_X1 U563 ( .A1(n501), .A2(n529), .ZN(n502) );
  XNOR2_X1 U564 ( .A(n503), .B(n502), .ZN(G1327GAT) );
  XOR2_X1 U565 ( .A(G29GAT), .B(KEYINPUT39), .Z(n505) );
  NAND2_X1 U566 ( .A1(n548), .A2(n507), .ZN(n504) );
  XNOR2_X1 U567 ( .A(n505), .B(n504), .ZN(G1328GAT) );
  NAND2_X1 U568 ( .A1(n507), .A2(n526), .ZN(n506) );
  XNOR2_X1 U569 ( .A(n506), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U570 ( .A1(n507), .A2(n529), .ZN(n508) );
  XNOR2_X1 U571 ( .A(n508), .B(KEYINPUT106), .ZN(n509) );
  XNOR2_X1 U572 ( .A(G50GAT), .B(n509), .ZN(G1331GAT) );
  NOR2_X1 U573 ( .A1(n551), .A2(n564), .ZN(n510) );
  XNOR2_X1 U574 ( .A(n510), .B(KEYINPUT108), .ZN(n522) );
  NAND2_X1 U575 ( .A1(n522), .A2(n511), .ZN(n512) );
  XNOR2_X1 U576 ( .A(n512), .B(KEYINPUT109), .ZN(n519) );
  NAND2_X1 U577 ( .A1(n519), .A2(n548), .ZN(n515) );
  XOR2_X1 U578 ( .A(G57GAT), .B(KEYINPUT107), .Z(n513) );
  XNOR2_X1 U579 ( .A(KEYINPUT42), .B(n513), .ZN(n514) );
  XNOR2_X1 U580 ( .A(n515), .B(n514), .ZN(G1332GAT) );
  NAND2_X1 U581 ( .A1(n519), .A2(n526), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n516), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U583 ( .A1(n535), .A2(n519), .ZN(n517) );
  XNOR2_X1 U584 ( .A(n517), .B(KEYINPUT110), .ZN(n518) );
  XNOR2_X1 U585 ( .A(G71GAT), .B(n518), .ZN(G1334GAT) );
  XOR2_X1 U586 ( .A(G78GAT), .B(KEYINPUT43), .Z(n521) );
  NAND2_X1 U587 ( .A1(n519), .A2(n529), .ZN(n520) );
  XNOR2_X1 U588 ( .A(n521), .B(n520), .ZN(G1335GAT) );
  AND2_X1 U589 ( .A1(n523), .A2(n522), .ZN(n530) );
  NAND2_X1 U590 ( .A1(n548), .A2(n530), .ZN(n524) );
  XOR2_X1 U591 ( .A(KEYINPUT111), .B(n524), .Z(n525) );
  XNOR2_X1 U592 ( .A(G85GAT), .B(n525), .ZN(G1336GAT) );
  NAND2_X1 U593 ( .A1(n530), .A2(n526), .ZN(n527) );
  XNOR2_X1 U594 ( .A(n527), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U595 ( .A1(n535), .A2(n530), .ZN(n528) );
  XNOR2_X1 U596 ( .A(n528), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT112), .B(KEYINPUT44), .Z(n532) );
  NAND2_X1 U598 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U599 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U600 ( .A(G106GAT), .B(n533), .Z(G1339GAT) );
  NAND2_X1 U601 ( .A1(n534), .A2(n535), .ZN(n536) );
  NOR2_X1 U602 ( .A1(n537), .A2(n536), .ZN(n545) );
  NAND2_X1 U603 ( .A1(n551), .A2(n545), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n538), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n541) );
  NAND2_X1 U606 ( .A1(n545), .A2(n539), .ZN(n540) );
  XNOR2_X1 U607 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U608 ( .A(G120GAT), .B(n542), .Z(G1341GAT) );
  NAND2_X1 U609 ( .A1(n557), .A2(n545), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n543), .B(KEYINPUT50), .ZN(n544) );
  XNOR2_X1 U611 ( .A(G127GAT), .B(n544), .ZN(G1342GAT) );
  XOR2_X1 U612 ( .A(G134GAT), .B(KEYINPUT51), .Z(n547) );
  NAND2_X1 U613 ( .A1(n545), .A2(n561), .ZN(n546) );
  XNOR2_X1 U614 ( .A(n547), .B(n546), .ZN(G1343GAT) );
  NAND2_X1 U615 ( .A1(n534), .A2(n548), .ZN(n549) );
  NOR2_X1 U616 ( .A1(n550), .A2(n549), .ZN(n560) );
  NAND2_X1 U617 ( .A1(n551), .A2(n560), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n552), .B(G141GAT), .ZN(G1344GAT) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(KEYINPUT116), .ZN(n556) );
  XOR2_X1 U620 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n554) );
  NAND2_X1 U621 ( .A1(n560), .A2(n539), .ZN(n553) );
  XNOR2_X1 U622 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(G1345GAT) );
  XOR2_X1 U624 ( .A(G155GAT), .B(KEYINPUT117), .Z(n559) );
  NAND2_X1 U625 ( .A1(n560), .A2(n557), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(G1346GAT) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U629 ( .A1(n563), .A2(n564), .ZN(n568) );
  XOR2_X1 U630 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n566) );
  XNOR2_X1 U631 ( .A(G176GAT), .B(KEYINPUT121), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(G1349GAT) );
  NAND2_X1 U634 ( .A1(n570), .A2(n569), .ZN(n585) );
  NOR2_X1 U635 ( .A1(n571), .A2(n585), .ZN(n576) );
  XOR2_X1 U636 ( .A(KEYINPUT60), .B(KEYINPUT124), .Z(n573) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(KEYINPUT123), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(KEYINPUT59), .B(n574), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n576), .B(n575), .ZN(G1352GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n579) );
  INV_X1 U642 ( .A(n585), .ZN(n577) );
  NAND2_X1 U643 ( .A1(n577), .A2(n453), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XOR2_X1 U645 ( .A(G204GAT), .B(n580), .Z(G1353GAT) );
  NOR2_X1 U646 ( .A1(n581), .A2(n585), .ZN(n582) );
  XOR2_X1 U647 ( .A(G211GAT), .B(n582), .Z(G1354GAT) );
  XOR2_X1 U648 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n584) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n584), .B(n583), .ZN(n588) );
  NOR2_X1 U651 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U652 ( .A(n588), .B(n587), .Z(G1355GAT) );
endmodule

