

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589;

  XOR2_X2 U325 ( .A(n446), .B(n410), .Z(n433) );
  XNOR2_X1 U326 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U327 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U328 ( .A(KEYINPUT45), .B(n437), .Z(n293) );
  INV_X1 U329 ( .A(KEYINPUT106), .ZN(n434) );
  XNOR2_X1 U330 ( .A(n459), .B(KEYINPUT122), .ZN(n460) );
  XNOR2_X1 U331 ( .A(n434), .B(KEYINPUT36), .ZN(n435) );
  XNOR2_X1 U332 ( .A(n568), .B(n435), .ZN(n586) );
  XNOR2_X1 U333 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U334 ( .A(n417), .B(n393), .Z(n564) );
  XNOR2_X1 U335 ( .A(n467), .B(G176GAT), .ZN(n468) );
  XNOR2_X1 U336 ( .A(n469), .B(n468), .ZN(G1349GAT) );
  XOR2_X1 U337 ( .A(KEYINPUT84), .B(KEYINPUT85), .Z(n295) );
  XNOR2_X1 U338 ( .A(G176GAT), .B(KEYINPUT83), .ZN(n294) );
  XNOR2_X1 U339 ( .A(n295), .B(n294), .ZN(n307) );
  XOR2_X1 U340 ( .A(KEYINPUT20), .B(G190GAT), .Z(n297) );
  XOR2_X1 U341 ( .A(G120GAT), .B(G71GAT), .Z(n407) );
  XOR2_X1 U342 ( .A(G15GAT), .B(G127GAT), .Z(n367) );
  XNOR2_X1 U343 ( .A(n407), .B(n367), .ZN(n296) );
  XNOR2_X1 U344 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U345 ( .A(n298), .B(G99GAT), .Z(n305) );
  XOR2_X1 U346 ( .A(KEYINPUT0), .B(KEYINPUT82), .Z(n300) );
  XNOR2_X1 U347 ( .A(G113GAT), .B(G134GAT), .ZN(n299) );
  XNOR2_X1 U348 ( .A(n300), .B(n299), .ZN(n339) );
  XOR2_X1 U349 ( .A(n339), .B(G183GAT), .Z(n302) );
  NAND2_X1 U350 ( .A1(G227GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U351 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U352 ( .A(G43GAT), .B(n303), .ZN(n304) );
  XNOR2_X1 U353 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U354 ( .A(n307), .B(n306), .ZN(n311) );
  XOR2_X1 U355 ( .A(KEYINPUT86), .B(KEYINPUT19), .Z(n309) );
  XNOR2_X1 U356 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n308) );
  XNOR2_X1 U357 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U358 ( .A(G169GAT), .B(n310), .Z(n445) );
  XOR2_X1 U359 ( .A(n311), .B(n445), .Z(n477) );
  XOR2_X1 U360 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n313) );
  XNOR2_X1 U361 ( .A(G204GAT), .B(KEYINPUT91), .ZN(n312) );
  XNOR2_X1 U362 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U363 ( .A(n314), .B(KEYINPUT90), .Z(n316) );
  XOR2_X1 U364 ( .A(G22GAT), .B(G155GAT), .Z(n366) );
  XNOR2_X1 U365 ( .A(n366), .B(KEYINPUT22), .ZN(n315) );
  XNOR2_X1 U366 ( .A(n316), .B(n315), .ZN(n321) );
  XNOR2_X1 U367 ( .A(G106GAT), .B(G78GAT), .ZN(n317) );
  XNOR2_X1 U368 ( .A(n317), .B(G148GAT), .ZN(n402) );
  XOR2_X1 U369 ( .A(G50GAT), .B(G162GAT), .Z(n423) );
  XOR2_X1 U370 ( .A(n402), .B(n423), .Z(n319) );
  NAND2_X1 U371 ( .A1(G228GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U372 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U373 ( .A(n321), .B(n320), .Z(n329) );
  XOR2_X1 U374 ( .A(KEYINPUT89), .B(KEYINPUT88), .Z(n323) );
  XNOR2_X1 U375 ( .A(KEYINPUT3), .B(KEYINPUT2), .ZN(n322) );
  XNOR2_X1 U376 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U377 ( .A(G141GAT), .B(n324), .Z(n352) );
  XOR2_X1 U378 ( .A(KEYINPUT87), .B(G218GAT), .Z(n326) );
  XNOR2_X1 U379 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n325) );
  XNOR2_X1 U380 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U381 ( .A(G197GAT), .B(n327), .Z(n447) );
  XNOR2_X1 U382 ( .A(n352), .B(n447), .ZN(n328) );
  XOR2_X1 U383 ( .A(n329), .B(n328), .Z(n475) );
  INV_X1 U384 ( .A(n475), .ZN(n478) );
  XOR2_X1 U385 ( .A(KEYINPUT95), .B(G148GAT), .Z(n331) );
  XNOR2_X1 U386 ( .A(G120GAT), .B(G127GAT), .ZN(n330) );
  XNOR2_X1 U387 ( .A(n331), .B(n330), .ZN(n335) );
  XOR2_X1 U388 ( .A(KEYINPUT5), .B(KEYINPUT96), .Z(n333) );
  XNOR2_X1 U389 ( .A(G1GAT), .B(KEYINPUT94), .ZN(n332) );
  XNOR2_X1 U390 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U391 ( .A(n335), .B(n334), .Z(n341) );
  XOR2_X1 U392 ( .A(G85GAT), .B(G155GAT), .Z(n337) );
  XNOR2_X1 U393 ( .A(G29GAT), .B(G162GAT), .ZN(n336) );
  XNOR2_X1 U394 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U395 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U396 ( .A(n341), .B(n340), .ZN(n348) );
  XOR2_X1 U397 ( .A(G57GAT), .B(KEYINPUT92), .Z(n343) );
  XNOR2_X1 U398 ( .A(KEYINPUT6), .B(KEYINPUT93), .ZN(n342) );
  XNOR2_X1 U399 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U400 ( .A(KEYINPUT97), .B(n344), .Z(n346) );
  NAND2_X1 U401 ( .A1(G225GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U402 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U403 ( .A(n348), .B(n347), .Z(n350) );
  XNOR2_X1 U404 ( .A(KEYINPUT4), .B(KEYINPUT1), .ZN(n349) );
  XNOR2_X1 U405 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U406 ( .A(n352), .B(n351), .ZN(n524) );
  XNOR2_X1 U407 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n444) );
  XOR2_X1 U408 ( .A(KEYINPUT47), .B(KEYINPUT115), .Z(n432) );
  XOR2_X1 U409 ( .A(KEYINPUT14), .B(KEYINPUT77), .Z(n354) );
  NAND2_X1 U410 ( .A1(G231GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U411 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U412 ( .A(KEYINPUT15), .B(n355), .ZN(n371) );
  XOR2_X1 U413 ( .A(G8GAT), .B(G183GAT), .Z(n448) );
  XOR2_X1 U414 ( .A(n448), .B(G78GAT), .Z(n357) );
  XOR2_X1 U415 ( .A(G1GAT), .B(KEYINPUT72), .Z(n386) );
  XNOR2_X1 U416 ( .A(n386), .B(G211GAT), .ZN(n356) );
  XNOR2_X1 U417 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U418 ( .A(n358), .B(G64GAT), .Z(n363) );
  XOR2_X1 U419 ( .A(KEYINPUT80), .B(KEYINPUT78), .Z(n360) );
  XNOR2_X1 U420 ( .A(KEYINPUT12), .B(KEYINPUT79), .ZN(n359) );
  XNOR2_X1 U421 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U422 ( .A(G71GAT), .B(n361), .ZN(n362) );
  XNOR2_X1 U423 ( .A(n363), .B(n362), .ZN(n365) );
  XNOR2_X1 U424 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n364) );
  XNOR2_X1 U425 ( .A(n364), .B(KEYINPUT74), .ZN(n397) );
  XNOR2_X1 U426 ( .A(n365), .B(n397), .ZN(n369) );
  XOR2_X1 U427 ( .A(n367), .B(n366), .Z(n368) );
  XOR2_X1 U428 ( .A(n369), .B(n368), .Z(n370) );
  XNOR2_X1 U429 ( .A(n371), .B(n370), .ZN(n583) );
  INV_X1 U430 ( .A(n583), .ZN(n566) );
  XOR2_X1 U431 ( .A(KEYINPUT71), .B(KEYINPUT7), .Z(n373) );
  XNOR2_X1 U432 ( .A(G43GAT), .B(G29GAT), .ZN(n372) );
  XNOR2_X1 U433 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U434 ( .A(KEYINPUT8), .B(n374), .ZN(n417) );
  XOR2_X1 U435 ( .A(G113GAT), .B(G15GAT), .Z(n376) );
  XNOR2_X1 U436 ( .A(G169GAT), .B(G22GAT), .ZN(n375) );
  XNOR2_X1 U437 ( .A(n376), .B(n375), .ZN(n380) );
  XOR2_X1 U438 ( .A(G8GAT), .B(KEYINPUT68), .Z(n378) );
  XNOR2_X1 U439 ( .A(KEYINPUT67), .B(KEYINPUT29), .ZN(n377) );
  XNOR2_X1 U440 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U441 ( .A(n380), .B(n379), .Z(n392) );
  XOR2_X1 U442 ( .A(KEYINPUT73), .B(KEYINPUT70), .Z(n382) );
  XNOR2_X1 U443 ( .A(KEYINPUT69), .B(KEYINPUT30), .ZN(n381) );
  XNOR2_X1 U444 ( .A(n382), .B(n381), .ZN(n390) );
  XOR2_X1 U445 ( .A(G197GAT), .B(G141GAT), .Z(n384) );
  XNOR2_X1 U446 ( .A(G36GAT), .B(G50GAT), .ZN(n383) );
  XNOR2_X1 U447 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U448 ( .A(n386), .B(n385), .Z(n388) );
  NAND2_X1 U449 ( .A1(G229GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U450 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U451 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U452 ( .A(n392), .B(n391), .ZN(n393) );
  INV_X1 U453 ( .A(n564), .ZN(n574) );
  INV_X1 U454 ( .A(KEYINPUT41), .ZN(n411) );
  XOR2_X1 U455 ( .A(KEYINPUT75), .B(G64GAT), .Z(n395) );
  XNOR2_X1 U456 ( .A(G204GAT), .B(G92GAT), .ZN(n394) );
  XNOR2_X1 U457 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U458 ( .A(G176GAT), .B(n396), .Z(n446) );
  XOR2_X1 U459 ( .A(G99GAT), .B(G85GAT), .Z(n418) );
  XOR2_X1 U460 ( .A(n418), .B(n397), .Z(n399) );
  NAND2_X1 U461 ( .A1(G230GAT), .A2(G233GAT), .ZN(n398) );
  XNOR2_X1 U462 ( .A(n399), .B(n398), .ZN(n401) );
  INV_X1 U463 ( .A(KEYINPUT31), .ZN(n400) );
  XNOR2_X1 U464 ( .A(n401), .B(n400), .ZN(n404) );
  XNOR2_X1 U465 ( .A(n402), .B(KEYINPUT33), .ZN(n403) );
  XNOR2_X1 U466 ( .A(n404), .B(n403), .ZN(n406) );
  INV_X1 U467 ( .A(KEYINPUT32), .ZN(n405) );
  XNOR2_X1 U468 ( .A(n406), .B(n405), .ZN(n409) );
  XNOR2_X1 U469 ( .A(n407), .B(KEYINPUT76), .ZN(n408) );
  XNOR2_X1 U470 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U471 ( .A(n411), .B(n433), .ZN(n466) );
  NOR2_X1 U472 ( .A1(n574), .A2(n466), .ZN(n412) );
  XNOR2_X1 U473 ( .A(n412), .B(KEYINPUT46), .ZN(n413) );
  NOR2_X1 U474 ( .A1(n566), .A2(n413), .ZN(n430) );
  XOR2_X1 U475 ( .A(KEYINPUT11), .B(KEYINPUT66), .Z(n415) );
  XNOR2_X1 U476 ( .A(G92GAT), .B(KEYINPUT10), .ZN(n414) );
  XNOR2_X1 U477 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U478 ( .A(n417), .B(n416), .Z(n429) );
  XOR2_X1 U479 ( .A(G36GAT), .B(G190GAT), .Z(n452) );
  XNOR2_X1 U480 ( .A(n452), .B(n418), .ZN(n420) );
  XOR2_X1 U481 ( .A(G134GAT), .B(G218GAT), .Z(n419) );
  XNOR2_X1 U482 ( .A(n420), .B(n419), .ZN(n427) );
  XOR2_X1 U483 ( .A(KEYINPUT9), .B(KEYINPUT65), .Z(n422) );
  NAND2_X1 U484 ( .A1(G232GAT), .A2(G233GAT), .ZN(n421) );
  XOR2_X1 U485 ( .A(n422), .B(n421), .Z(n425) );
  XNOR2_X1 U486 ( .A(n423), .B(G106GAT), .ZN(n424) );
  XOR2_X1 U487 ( .A(n429), .B(n428), .Z(n568) );
  INV_X1 U488 ( .A(n568), .ZN(n562) );
  NAND2_X1 U489 ( .A1(n430), .A2(n562), .ZN(n431) );
  XNOR2_X1 U490 ( .A(n432), .B(n431), .ZN(n442) );
  INV_X1 U491 ( .A(n433), .ZN(n438) );
  NOR2_X1 U492 ( .A1(n583), .A2(n586), .ZN(n436) );
  XNOR2_X1 U493 ( .A(n436), .B(KEYINPUT116), .ZN(n437) );
  NOR2_X1 U494 ( .A1(n438), .A2(n293), .ZN(n439) );
  XNOR2_X1 U495 ( .A(n439), .B(KEYINPUT117), .ZN(n440) );
  NOR2_X1 U496 ( .A1(n440), .A2(n564), .ZN(n441) );
  NOR2_X1 U497 ( .A1(n442), .A2(n441), .ZN(n443) );
  XNOR2_X1 U498 ( .A(n444), .B(n443), .ZN(n537) );
  INV_X1 U499 ( .A(n445), .ZN(n458) );
  XNOR2_X1 U500 ( .A(n447), .B(n446), .ZN(n456) );
  XOR2_X1 U501 ( .A(n448), .B(KEYINPUT100), .Z(n450) );
  NAND2_X1 U502 ( .A1(G226GAT), .A2(G233GAT), .ZN(n449) );
  XNOR2_X1 U503 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U504 ( .A(n451), .B(KEYINPUT99), .Z(n454) );
  XNOR2_X1 U505 ( .A(n452), .B(KEYINPUT98), .ZN(n453) );
  XNOR2_X1 U506 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U507 ( .A(n456), .B(n455), .ZN(n457) );
  XOR2_X1 U508 ( .A(n458), .B(n457), .Z(n473) );
  NOR2_X1 U509 ( .A1(n537), .A2(n473), .ZN(n461) );
  XNOR2_X1 U510 ( .A(KEYINPUT123), .B(KEYINPUT54), .ZN(n459) );
  NOR2_X1 U511 ( .A1(n524), .A2(n462), .ZN(n573) );
  NAND2_X1 U512 ( .A1(n478), .A2(n573), .ZN(n464) );
  INV_X1 U513 ( .A(KEYINPUT55), .ZN(n463) );
  XNOR2_X1 U514 ( .A(n464), .B(n463), .ZN(n465) );
  NOR2_X2 U515 ( .A1(n477), .A2(n465), .ZN(n569) );
  INV_X1 U516 ( .A(n466), .ZN(n542) );
  NAND2_X1 U517 ( .A1(n569), .A2(n542), .ZN(n469) );
  XOR2_X1 U518 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n467) );
  XOR2_X1 U519 ( .A(KEYINPUT34), .B(KEYINPUT105), .Z(n491) );
  XNOR2_X1 U520 ( .A(KEYINPUT27), .B(KEYINPUT101), .ZN(n470) );
  INV_X1 U521 ( .A(n473), .ZN(n527) );
  XOR2_X1 U522 ( .A(n470), .B(n527), .Z(n480) );
  NAND2_X1 U523 ( .A1(n480), .A2(n524), .ZN(n471) );
  XNOR2_X1 U524 ( .A(n471), .B(KEYINPUT102), .ZN(n552) );
  XNOR2_X1 U525 ( .A(n475), .B(KEYINPUT28), .ZN(n531) );
  NOR2_X1 U526 ( .A1(n552), .A2(n531), .ZN(n538) );
  NAND2_X1 U527 ( .A1(n538), .A2(n477), .ZN(n472) );
  XNOR2_X1 U528 ( .A(n472), .B(KEYINPUT103), .ZN(n485) );
  NOR2_X1 U529 ( .A1(n477), .A2(n473), .ZN(n474) );
  NOR2_X1 U530 ( .A1(n475), .A2(n474), .ZN(n476) );
  XOR2_X1 U531 ( .A(KEYINPUT25), .B(n476), .Z(n482) );
  INV_X1 U532 ( .A(n477), .ZN(n539) );
  NOR2_X1 U533 ( .A1(n539), .A2(n478), .ZN(n479) );
  XNOR2_X1 U534 ( .A(KEYINPUT26), .B(n479), .ZN(n572) );
  AND2_X1 U535 ( .A1(n572), .A2(n480), .ZN(n481) );
  NOR2_X1 U536 ( .A1(n482), .A2(n481), .ZN(n483) );
  NOR2_X1 U537 ( .A1(n524), .A2(n483), .ZN(n484) );
  NOR2_X1 U538 ( .A1(n485), .A2(n484), .ZN(n498) );
  XOR2_X1 U539 ( .A(KEYINPUT16), .B(KEYINPUT81), .Z(n487) );
  NAND2_X1 U540 ( .A1(n566), .A2(n562), .ZN(n486) );
  XNOR2_X1 U541 ( .A(n487), .B(n486), .ZN(n488) );
  NOR2_X1 U542 ( .A1(n498), .A2(n488), .ZN(n489) );
  XOR2_X1 U543 ( .A(KEYINPUT104), .B(n489), .Z(n511) );
  NAND2_X1 U544 ( .A1(n564), .A2(n433), .ZN(n501) );
  NOR2_X1 U545 ( .A1(n511), .A2(n501), .ZN(n496) );
  NAND2_X1 U546 ( .A1(n496), .A2(n524), .ZN(n490) );
  XNOR2_X1 U547 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U548 ( .A(G1GAT), .B(n492), .ZN(G1324GAT) );
  NAND2_X1 U549 ( .A1(n496), .A2(n527), .ZN(n493) );
  XNOR2_X1 U550 ( .A(n493), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U551 ( .A(G15GAT), .B(KEYINPUT35), .Z(n495) );
  NAND2_X1 U552 ( .A1(n496), .A2(n539), .ZN(n494) );
  XNOR2_X1 U553 ( .A(n495), .B(n494), .ZN(G1326GAT) );
  NAND2_X1 U554 ( .A1(n496), .A2(n531), .ZN(n497) );
  XNOR2_X1 U555 ( .A(n497), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U556 ( .A(G29GAT), .B(KEYINPUT39), .Z(n504) );
  NOR2_X1 U557 ( .A1(n586), .A2(n498), .ZN(n499) );
  NAND2_X1 U558 ( .A1(n583), .A2(n499), .ZN(n500) );
  XOR2_X1 U559 ( .A(n500), .B(KEYINPUT37), .Z(n523) );
  OR2_X1 U560 ( .A1(n523), .A2(n501), .ZN(n502) );
  XOR2_X1 U561 ( .A(KEYINPUT38), .B(n502), .Z(n509) );
  NAND2_X1 U562 ( .A1(n509), .A2(n524), .ZN(n503) );
  XNOR2_X1 U563 ( .A(n504), .B(n503), .ZN(G1328GAT) );
  NAND2_X1 U564 ( .A1(n527), .A2(n509), .ZN(n505) );
  XNOR2_X1 U565 ( .A(G36GAT), .B(n505), .ZN(G1329GAT) );
  XOR2_X1 U566 ( .A(KEYINPUT40), .B(KEYINPUT107), .Z(n507) );
  NAND2_X1 U567 ( .A1(n539), .A2(n509), .ZN(n506) );
  XNOR2_X1 U568 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U569 ( .A(G43GAT), .B(n508), .ZN(G1330GAT) );
  NAND2_X1 U570 ( .A1(n509), .A2(n531), .ZN(n510) );
  XNOR2_X1 U571 ( .A(n510), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U572 ( .A(KEYINPUT108), .B(KEYINPUT42), .Z(n513) );
  NAND2_X1 U573 ( .A1(n574), .A2(n542), .ZN(n522) );
  NOR2_X1 U574 ( .A1(n511), .A2(n522), .ZN(n518) );
  NAND2_X1 U575 ( .A1(n518), .A2(n524), .ZN(n512) );
  XNOR2_X1 U576 ( .A(n513), .B(n512), .ZN(n514) );
  XOR2_X1 U577 ( .A(G57GAT), .B(n514), .Z(G1332GAT) );
  XOR2_X1 U578 ( .A(G64GAT), .B(KEYINPUT109), .Z(n516) );
  NAND2_X1 U579 ( .A1(n518), .A2(n527), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n516), .B(n515), .ZN(G1333GAT) );
  NAND2_X1 U581 ( .A1(n518), .A2(n539), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n517), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U583 ( .A(KEYINPUT110), .B(KEYINPUT43), .Z(n520) );
  NAND2_X1 U584 ( .A1(n518), .A2(n531), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U586 ( .A(G78GAT), .B(n521), .ZN(G1335GAT) );
  XOR2_X1 U587 ( .A(G85GAT), .B(KEYINPUT111), .Z(n526) );
  NOR2_X1 U588 ( .A1(n523), .A2(n522), .ZN(n532) );
  NAND2_X1 U589 ( .A1(n532), .A2(n524), .ZN(n525) );
  XNOR2_X1 U590 ( .A(n526), .B(n525), .ZN(G1336GAT) );
  NAND2_X1 U591 ( .A1(n532), .A2(n527), .ZN(n528) );
  XNOR2_X1 U592 ( .A(n528), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U593 ( .A1(n532), .A2(n539), .ZN(n529) );
  XNOR2_X1 U594 ( .A(n529), .B(KEYINPUT112), .ZN(n530) );
  XNOR2_X1 U595 ( .A(G99GAT), .B(n530), .ZN(G1338GAT) );
  XNOR2_X1 U596 ( .A(G106GAT), .B(KEYINPUT113), .ZN(n536) );
  XOR2_X1 U597 ( .A(KEYINPUT44), .B(KEYINPUT114), .Z(n534) );
  NAND2_X1 U598 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U599 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U600 ( .A(n536), .B(n535), .ZN(G1339GAT) );
  NAND2_X1 U601 ( .A1(n539), .A2(n538), .ZN(n540) );
  NOR2_X1 U602 ( .A1(n537), .A2(n540), .ZN(n548) );
  NAND2_X1 U603 ( .A1(n564), .A2(n548), .ZN(n541) );
  XNOR2_X1 U604 ( .A(n541), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT49), .B(KEYINPUT118), .Z(n544) );
  NAND2_X1 U606 ( .A1(n548), .A2(n542), .ZN(n543) );
  XNOR2_X1 U607 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U608 ( .A(G120GAT), .B(n545), .ZN(G1341GAT) );
  NAND2_X1 U609 ( .A1(n548), .A2(n566), .ZN(n546) );
  XNOR2_X1 U610 ( .A(n546), .B(KEYINPUT50), .ZN(n547) );
  XNOR2_X1 U611 ( .A(G127GAT), .B(n547), .ZN(G1342GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT51), .B(KEYINPUT119), .Z(n550) );
  NAND2_X1 U613 ( .A1(n548), .A2(n568), .ZN(n549) );
  XNOR2_X1 U614 ( .A(n550), .B(n549), .ZN(n551) );
  XOR2_X1 U615 ( .A(G134GAT), .B(n551), .Z(G1343GAT) );
  NOR2_X1 U616 ( .A1(n537), .A2(n552), .ZN(n553) );
  NAND2_X1 U617 ( .A1(n553), .A2(n572), .ZN(n561) );
  NOR2_X1 U618 ( .A1(n574), .A2(n561), .ZN(n554) );
  XOR2_X1 U619 ( .A(G141GAT), .B(n554), .Z(G1344GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT53), .B(KEYINPUT120), .Z(n556) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(n558) );
  NOR2_X1 U623 ( .A1(n466), .A2(n561), .ZN(n557) );
  XOR2_X1 U624 ( .A(n558), .B(n557), .Z(G1345GAT) );
  NOR2_X1 U625 ( .A1(n583), .A2(n561), .ZN(n560) );
  XNOR2_X1 U626 ( .A(G155GAT), .B(KEYINPUT121), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(G1346GAT) );
  NOR2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U629 ( .A(G162GAT), .B(n563), .Z(G1347GAT) );
  NAND2_X1 U630 ( .A1(n564), .A2(n569), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U632 ( .A1(n569), .A2(n566), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n567), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U634 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n571) );
  NAND2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1351GAT) );
  NAND2_X1 U637 ( .A1(n573), .A2(n572), .ZN(n585) );
  NOR2_X1 U638 ( .A1(n574), .A2(n585), .ZN(n578) );
  XNOR2_X1 U639 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(KEYINPUT60), .ZN(n576) );
  XNOR2_X1 U641 ( .A(KEYINPUT124), .B(n576), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n578), .B(n577), .ZN(G1352GAT) );
  NOR2_X1 U643 ( .A1(n585), .A2(n433), .ZN(n582) );
  XOR2_X1 U644 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n580) );
  XNOR2_X1 U645 ( .A(G204GAT), .B(KEYINPUT126), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1353GAT) );
  NOR2_X1 U648 ( .A1(n583), .A2(n585), .ZN(n584) );
  XOR2_X1 U649 ( .A(G211GAT), .B(n584), .Z(G1354GAT) );
  NOR2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n588) );
  XNOR2_X1 U651 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n588), .B(n587), .ZN(n589) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(n589), .ZN(G1355GAT) );
endmodule

