

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587;

  XNOR2_X1 U327 ( .A(KEYINPUT26), .B(n465), .ZN(n570) );
  XNOR2_X1 U328 ( .A(n437), .B(n436), .ZN(n471) );
  XOR2_X1 U329 ( .A(n332), .B(n352), .Z(n580) );
  XOR2_X1 U330 ( .A(G148GAT), .B(KEYINPUT2), .Z(n295) );
  INV_X1 U331 ( .A(G78GAT), .ZN(n427) );
  XNOR2_X1 U332 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U333 ( .A(n430), .B(n429), .ZN(n433) );
  XNOR2_X1 U334 ( .A(n323), .B(n322), .ZN(n324) );
  NAND2_X1 U335 ( .A1(n478), .A2(n477), .ZN(n479) );
  XNOR2_X1 U336 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U337 ( .A(n479), .B(KEYINPUT102), .ZN(n492) );
  NOR2_X1 U338 ( .A1(n518), .A2(n496), .ZN(n497) );
  XOR2_X1 U339 ( .A(KEYINPUT28), .B(n471), .Z(n534) );
  XNOR2_X1 U340 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U341 ( .A(n463), .B(n462), .ZN(G1351GAT) );
  XOR2_X1 U342 ( .A(G29GAT), .B(KEYINPUT7), .Z(n297) );
  XNOR2_X1 U343 ( .A(KEYINPUT8), .B(G43GAT), .ZN(n296) );
  XNOR2_X1 U344 ( .A(n297), .B(n296), .ZN(n299) );
  XOR2_X1 U345 ( .A(KEYINPUT68), .B(KEYINPUT67), .Z(n298) );
  XOR2_X1 U346 ( .A(n299), .B(n298), .Z(n342) );
  INV_X1 U347 ( .A(n342), .ZN(n315) );
  XOR2_X1 U348 ( .A(KEYINPUT9), .B(KEYINPUT77), .Z(n301) );
  XOR2_X1 U349 ( .A(G134GAT), .B(KEYINPUT76), .Z(n405) );
  XOR2_X1 U350 ( .A(G36GAT), .B(G190GAT), .Z(n380) );
  XNOR2_X1 U351 ( .A(n405), .B(n380), .ZN(n300) );
  XNOR2_X1 U352 ( .A(n301), .B(n300), .ZN(n311) );
  XOR2_X1 U353 ( .A(KEYINPUT10), .B(G92GAT), .Z(n303) );
  NAND2_X1 U354 ( .A1(G232GAT), .A2(G233GAT), .ZN(n302) );
  XOR2_X1 U355 ( .A(n303), .B(n302), .Z(n304) );
  XNOR2_X1 U356 ( .A(n304), .B(KEYINPUT11), .ZN(n309) );
  XNOR2_X1 U357 ( .A(G50GAT), .B(KEYINPUT75), .ZN(n305) );
  XNOR2_X1 U358 ( .A(n305), .B(G162GAT), .ZN(n431) );
  XOR2_X1 U359 ( .A(KEYINPUT72), .B(G85GAT), .Z(n307) );
  XNOR2_X1 U360 ( .A(G99GAT), .B(G106GAT), .ZN(n306) );
  XNOR2_X1 U361 ( .A(n307), .B(n306), .ZN(n358) );
  XNOR2_X1 U362 ( .A(n431), .B(n358), .ZN(n308) );
  XNOR2_X1 U363 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U364 ( .A(n311), .B(n310), .Z(n313) );
  XNOR2_X1 U365 ( .A(G218GAT), .B(KEYINPUT65), .ZN(n312) );
  XNOR2_X1 U366 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U367 ( .A(n315), .B(n314), .Z(n480) );
  INV_X1 U368 ( .A(n480), .ZN(n557) );
  XOR2_X1 U369 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n317) );
  XNOR2_X1 U370 ( .A(KEYINPUT14), .B(KEYINPUT79), .ZN(n316) );
  XNOR2_X1 U371 ( .A(n317), .B(n316), .ZN(n327) );
  XOR2_X1 U372 ( .A(KEYINPUT78), .B(G211GAT), .Z(n319) );
  XNOR2_X1 U373 ( .A(G8GAT), .B(G183GAT), .ZN(n318) );
  XNOR2_X1 U374 ( .A(n319), .B(n318), .ZN(n383) );
  XOR2_X1 U375 ( .A(G15GAT), .B(G127GAT), .Z(n448) );
  XOR2_X1 U376 ( .A(n383), .B(n448), .Z(n321) );
  NAND2_X1 U377 ( .A1(G231GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U378 ( .A(n321), .B(n320), .ZN(n325) );
  XOR2_X1 U379 ( .A(G22GAT), .B(G155GAT), .Z(n426) );
  XNOR2_X1 U380 ( .A(G1GAT), .B(n426), .ZN(n323) );
  INV_X1 U381 ( .A(G64GAT), .ZN(n322) );
  XNOR2_X1 U382 ( .A(n327), .B(n326), .ZN(n332) );
  XOR2_X1 U383 ( .A(KEYINPUT70), .B(KEYINPUT13), .Z(n329) );
  XNOR2_X1 U384 ( .A(G57GAT), .B(KEYINPUT71), .ZN(n328) );
  XNOR2_X1 U385 ( .A(n329), .B(n328), .ZN(n331) );
  XOR2_X1 U386 ( .A(G71GAT), .B(G78GAT), .Z(n330) );
  XOR2_X1 U387 ( .A(n331), .B(n330), .Z(n352) );
  XNOR2_X1 U388 ( .A(KEYINPUT112), .B(n580), .ZN(n567) );
  XOR2_X1 U389 ( .A(KEYINPUT66), .B(G8GAT), .Z(n334) );
  XNOR2_X1 U390 ( .A(G197GAT), .B(G22GAT), .ZN(n333) );
  XNOR2_X1 U391 ( .A(n334), .B(n333), .ZN(n348) );
  NAND2_X1 U392 ( .A1(G229GAT), .A2(G233GAT), .ZN(n340) );
  XOR2_X1 U393 ( .A(G141GAT), .B(G113GAT), .Z(n336) );
  XNOR2_X1 U394 ( .A(G169GAT), .B(G15GAT), .ZN(n335) );
  XNOR2_X1 U395 ( .A(n336), .B(n335), .ZN(n338) );
  XOR2_X1 U396 ( .A(G50GAT), .B(G36GAT), .Z(n337) );
  XNOR2_X1 U397 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U398 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U399 ( .A(n342), .B(n341), .Z(n346) );
  XOR2_X1 U400 ( .A(KEYINPUT29), .B(G1GAT), .Z(n344) );
  XNOR2_X1 U401 ( .A(KEYINPUT30), .B(KEYINPUT69), .ZN(n343) );
  XNOR2_X1 U402 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U403 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U404 ( .A(n348), .B(n347), .Z(n535) );
  INV_X1 U405 ( .A(n535), .ZN(n572) );
  XOR2_X1 U406 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n350) );
  XNOR2_X1 U407 ( .A(G120GAT), .B(G148GAT), .ZN(n349) );
  XNOR2_X1 U408 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U409 ( .A(n352), .B(n351), .ZN(n362) );
  XOR2_X1 U410 ( .A(KEYINPUT74), .B(KEYINPUT73), .Z(n354) );
  NAND2_X1 U411 ( .A1(G230GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U412 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U413 ( .A(n355), .B(KEYINPUT31), .Z(n360) );
  XOR2_X1 U414 ( .A(G64GAT), .B(G92GAT), .Z(n357) );
  XNOR2_X1 U415 ( .A(G176GAT), .B(G204GAT), .ZN(n356) );
  XNOR2_X1 U416 ( .A(n357), .B(n356), .ZN(n389) );
  XNOR2_X1 U417 ( .A(n358), .B(n389), .ZN(n359) );
  XNOR2_X1 U418 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U419 ( .A(n362), .B(n361), .Z(n576) );
  XOR2_X1 U420 ( .A(KEYINPUT41), .B(n576), .Z(n564) );
  NOR2_X1 U421 ( .A1(n572), .A2(n564), .ZN(n364) );
  XNOR2_X1 U422 ( .A(KEYINPUT46), .B(KEYINPUT113), .ZN(n363) );
  XNOR2_X1 U423 ( .A(n364), .B(n363), .ZN(n365) );
  NAND2_X1 U424 ( .A1(n567), .A2(n365), .ZN(n366) );
  NOR2_X1 U425 ( .A1(n480), .A2(n366), .ZN(n367) );
  XOR2_X1 U426 ( .A(KEYINPUT47), .B(n367), .Z(n375) );
  XNOR2_X1 U427 ( .A(KEYINPUT36), .B(KEYINPUT105), .ZN(n368) );
  XOR2_X1 U428 ( .A(n368), .B(n557), .Z(n584) );
  NOR2_X1 U429 ( .A1(n580), .A2(n584), .ZN(n369) );
  XNOR2_X1 U430 ( .A(n369), .B(KEYINPUT45), .ZN(n372) );
  INV_X1 U431 ( .A(n576), .ZN(n370) );
  NOR2_X1 U432 ( .A1(n535), .A2(n370), .ZN(n371) );
  AND2_X1 U433 ( .A1(n372), .A2(n371), .ZN(n373) );
  XNOR2_X1 U434 ( .A(n373), .B(KEYINPUT114), .ZN(n374) );
  NOR2_X1 U435 ( .A1(n375), .A2(n374), .ZN(n376) );
  XNOR2_X1 U436 ( .A(KEYINPUT48), .B(n376), .ZN(n531) );
  XOR2_X1 U437 ( .A(KEYINPUT92), .B(G218GAT), .Z(n378) );
  XNOR2_X1 U438 ( .A(KEYINPUT93), .B(KEYINPUT21), .ZN(n377) );
  XNOR2_X1 U439 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U440 ( .A(G197GAT), .B(n379), .Z(n437) );
  XOR2_X1 U441 ( .A(n380), .B(n437), .Z(n382) );
  NAND2_X1 U442 ( .A1(G226GAT), .A2(G233GAT), .ZN(n381) );
  XNOR2_X1 U443 ( .A(n382), .B(n381), .ZN(n384) );
  XOR2_X1 U444 ( .A(n384), .B(n383), .Z(n391) );
  XNOR2_X1 U445 ( .A(KEYINPUT86), .B(KEYINPUT17), .ZN(n385) );
  XNOR2_X1 U446 ( .A(n385), .B(KEYINPUT87), .ZN(n386) );
  XOR2_X1 U447 ( .A(n386), .B(KEYINPUT19), .Z(n388) );
  XNOR2_X1 U448 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n387) );
  XNOR2_X1 U449 ( .A(n388), .B(n387), .ZN(n458) );
  XNOR2_X1 U450 ( .A(n458), .B(n389), .ZN(n390) );
  XNOR2_X1 U451 ( .A(n391), .B(n390), .ZN(n522) );
  XOR2_X1 U452 ( .A(KEYINPUT120), .B(n522), .Z(n392) );
  NOR2_X1 U453 ( .A1(n531), .A2(n392), .ZN(n393) );
  XNOR2_X1 U454 ( .A(KEYINPUT54), .B(n393), .ZN(n417) );
  XOR2_X1 U455 ( .A(KEYINPUT1), .B(G57GAT), .Z(n395) );
  XNOR2_X1 U456 ( .A(G1GAT), .B(G155GAT), .ZN(n394) );
  XNOR2_X1 U457 ( .A(n395), .B(n394), .ZN(n399) );
  XOR2_X1 U458 ( .A(KEYINPUT97), .B(KEYINPUT95), .Z(n397) );
  XNOR2_X1 U459 ( .A(KEYINPUT98), .B(KEYINPUT96), .ZN(n396) );
  XNOR2_X1 U460 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U461 ( .A(n399), .B(n398), .Z(n411) );
  XOR2_X1 U462 ( .A(KEYINPUT99), .B(KEYINPUT4), .Z(n401) );
  XNOR2_X1 U463 ( .A(KEYINPUT6), .B(KEYINPUT5), .ZN(n400) );
  XNOR2_X1 U464 ( .A(n401), .B(n400), .ZN(n409) );
  XOR2_X1 U465 ( .A(G85GAT), .B(G162GAT), .Z(n403) );
  XNOR2_X1 U466 ( .A(G29GAT), .B(G127GAT), .ZN(n402) );
  XNOR2_X1 U467 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U468 ( .A(n405), .B(n404), .Z(n407) );
  NAND2_X1 U469 ( .A1(G225GAT), .A2(G233GAT), .ZN(n406) );
  XNOR2_X1 U470 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U471 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U472 ( .A(n411), .B(n410), .ZN(n416) );
  XOR2_X1 U473 ( .A(G120GAT), .B(KEYINPUT81), .Z(n413) );
  XNOR2_X1 U474 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n412) );
  XNOR2_X1 U475 ( .A(n413), .B(n412), .ZN(n452) );
  XNOR2_X1 U476 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n414) );
  XNOR2_X1 U477 ( .A(n295), .B(n414), .ZN(n425) );
  XOR2_X1 U478 ( .A(n452), .B(n425), .Z(n415) );
  XOR2_X1 U479 ( .A(n416), .B(n415), .Z(n472) );
  AND2_X1 U480 ( .A1(n417), .A2(n472), .ZN(n418) );
  XNOR2_X1 U481 ( .A(n418), .B(KEYINPUT64), .ZN(n571) );
  XOR2_X1 U482 ( .A(G204GAT), .B(KEYINPUT22), .Z(n420) );
  XNOR2_X1 U483 ( .A(KEYINPUT91), .B(KEYINPUT24), .ZN(n419) );
  XNOR2_X1 U484 ( .A(n420), .B(n419), .ZN(n424) );
  XOR2_X1 U485 ( .A(KEYINPUT90), .B(KEYINPUT23), .Z(n422) );
  XNOR2_X1 U486 ( .A(G106GAT), .B(KEYINPUT94), .ZN(n421) );
  XNOR2_X1 U487 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U488 ( .A(n424), .B(n423), .ZN(n435) );
  XOR2_X1 U489 ( .A(n426), .B(n425), .Z(n430) );
  NAND2_X1 U490 ( .A1(G228GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U491 ( .A(n431), .B(G211GAT), .ZN(n432) );
  XNOR2_X1 U492 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U493 ( .A(n435), .B(n434), .ZN(n436) );
  NAND2_X1 U494 ( .A1(n571), .A2(n471), .ZN(n438) );
  XNOR2_X1 U495 ( .A(n438), .B(KEYINPUT55), .ZN(n459) );
  XOR2_X1 U496 ( .A(KEYINPUT20), .B(G176GAT), .Z(n440) );
  XNOR2_X1 U497 ( .A(KEYINPUT89), .B(KEYINPUT83), .ZN(n439) );
  XNOR2_X1 U498 ( .A(n440), .B(n439), .ZN(n444) );
  XOR2_X1 U499 ( .A(KEYINPUT85), .B(KEYINPUT88), .Z(n442) );
  XNOR2_X1 U500 ( .A(KEYINPUT82), .B(G71GAT), .ZN(n441) );
  XNOR2_X1 U501 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U502 ( .A(n444), .B(n443), .ZN(n456) );
  XOR2_X1 U503 ( .A(G99GAT), .B(G190GAT), .Z(n446) );
  XNOR2_X1 U504 ( .A(G43GAT), .B(G134GAT), .ZN(n445) );
  XNOR2_X1 U505 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U506 ( .A(n448), .B(n447), .Z(n450) );
  NAND2_X1 U507 ( .A1(G227GAT), .A2(G233GAT), .ZN(n449) );
  XNOR2_X1 U508 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U509 ( .A(n451), .B(G183GAT), .Z(n454) );
  XNOR2_X1 U510 ( .A(n452), .B(KEYINPUT84), .ZN(n453) );
  XNOR2_X1 U511 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U512 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X2 U513 ( .A(n458), .B(n457), .ZN(n532) );
  NAND2_X1 U514 ( .A1(n459), .A2(n532), .ZN(n559) );
  NOR2_X1 U515 ( .A1(n557), .A2(n559), .ZN(n463) );
  XNOR2_X1 U516 ( .A(KEYINPUT124), .B(KEYINPUT58), .ZN(n461) );
  INV_X1 U517 ( .A(G190GAT), .ZN(n460) );
  XNOR2_X1 U518 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n485) );
  NAND2_X1 U519 ( .A1(n535), .A2(n576), .ZN(n496) );
  XNOR2_X1 U520 ( .A(n522), .B(KEYINPUT27), .ZN(n473) );
  NOR2_X1 U521 ( .A1(n532), .A2(n471), .ZN(n464) );
  XOR2_X1 U522 ( .A(KEYINPUT101), .B(n464), .Z(n465) );
  NAND2_X1 U523 ( .A1(n473), .A2(n570), .ZN(n469) );
  NAND2_X1 U524 ( .A1(n522), .A2(n532), .ZN(n466) );
  NAND2_X1 U525 ( .A1(n471), .A2(n466), .ZN(n467) );
  XOR2_X1 U526 ( .A(KEYINPUT25), .B(n467), .Z(n468) );
  NAND2_X1 U527 ( .A1(n469), .A2(n468), .ZN(n470) );
  NAND2_X1 U528 ( .A1(n470), .A2(n472), .ZN(n478) );
  INV_X1 U529 ( .A(n534), .ZN(n475) );
  INV_X1 U530 ( .A(n472), .ZN(n519) );
  NAND2_X1 U531 ( .A1(n519), .A2(n473), .ZN(n530) );
  NOR2_X1 U532 ( .A1(n532), .A2(n530), .ZN(n474) );
  NAND2_X1 U533 ( .A1(n475), .A2(n474), .ZN(n476) );
  XNOR2_X1 U534 ( .A(n476), .B(KEYINPUT100), .ZN(n477) );
  NOR2_X1 U535 ( .A1(n480), .A2(n580), .ZN(n482) );
  XNOR2_X1 U536 ( .A(KEYINPUT80), .B(KEYINPUT16), .ZN(n481) );
  XNOR2_X1 U537 ( .A(n482), .B(n481), .ZN(n483) );
  NAND2_X1 U538 ( .A1(n492), .A2(n483), .ZN(n508) );
  NOR2_X1 U539 ( .A1(n496), .A2(n508), .ZN(n490) );
  NAND2_X1 U540 ( .A1(n490), .A2(n519), .ZN(n484) );
  XNOR2_X1 U541 ( .A(n485), .B(n484), .ZN(G1324GAT) );
  NAND2_X1 U542 ( .A1(n490), .A2(n522), .ZN(n486) );
  XNOR2_X1 U543 ( .A(n486), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U544 ( .A(KEYINPUT103), .B(KEYINPUT35), .Z(n488) );
  NAND2_X1 U545 ( .A1(n490), .A2(n532), .ZN(n487) );
  XNOR2_X1 U546 ( .A(n488), .B(n487), .ZN(n489) );
  XOR2_X1 U547 ( .A(G15GAT), .B(n489), .Z(G1326GAT) );
  NAND2_X1 U548 ( .A1(n534), .A2(n490), .ZN(n491) );
  XNOR2_X1 U549 ( .A(n491), .B(G22GAT), .ZN(G1327GAT) );
  INV_X1 U550 ( .A(n492), .ZN(n493) );
  NOR2_X1 U551 ( .A1(n584), .A2(n493), .ZN(n494) );
  NAND2_X1 U552 ( .A1(n580), .A2(n494), .ZN(n495) );
  XOR2_X1 U553 ( .A(KEYINPUT37), .B(n495), .Z(n518) );
  XNOR2_X1 U554 ( .A(KEYINPUT38), .B(n497), .ZN(n504) );
  NAND2_X1 U555 ( .A1(n504), .A2(n519), .ZN(n499) );
  XOR2_X1 U556 ( .A(G29GAT), .B(KEYINPUT39), .Z(n498) );
  XNOR2_X1 U557 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U558 ( .A(KEYINPUT104), .B(n500), .ZN(G1328GAT) );
  NAND2_X1 U559 ( .A1(n504), .A2(n522), .ZN(n501) );
  XNOR2_X1 U560 ( .A(n501), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U561 ( .A1(n504), .A2(n532), .ZN(n502) );
  XNOR2_X1 U562 ( .A(n502), .B(KEYINPUT40), .ZN(n503) );
  XNOR2_X1 U563 ( .A(G43GAT), .B(n503), .ZN(G1330GAT) );
  XNOR2_X1 U564 ( .A(G50GAT), .B(KEYINPUT106), .ZN(n506) );
  NAND2_X1 U565 ( .A1(n534), .A2(n504), .ZN(n505) );
  XNOR2_X1 U566 ( .A(n506), .B(n505), .ZN(G1331GAT) );
  XNOR2_X1 U567 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n510) );
  NOR2_X1 U568 ( .A1(n564), .A2(n535), .ZN(n507) );
  XNOR2_X1 U569 ( .A(n507), .B(KEYINPUT107), .ZN(n517) );
  NOR2_X1 U570 ( .A1(n517), .A2(n508), .ZN(n513) );
  NAND2_X1 U571 ( .A1(n513), .A2(n519), .ZN(n509) );
  XNOR2_X1 U572 ( .A(n510), .B(n509), .ZN(G1332GAT) );
  NAND2_X1 U573 ( .A1(n513), .A2(n522), .ZN(n511) );
  XNOR2_X1 U574 ( .A(n511), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U575 ( .A1(n532), .A2(n513), .ZN(n512) );
  XNOR2_X1 U576 ( .A(n512), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U577 ( .A(KEYINPUT108), .B(KEYINPUT43), .Z(n515) );
  NAND2_X1 U578 ( .A1(n513), .A2(n534), .ZN(n514) );
  XNOR2_X1 U579 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U580 ( .A(G78GAT), .B(n516), .ZN(G1335GAT) );
  XOR2_X1 U581 ( .A(G85GAT), .B(KEYINPUT109), .Z(n521) );
  NOR2_X1 U582 ( .A1(n518), .A2(n517), .ZN(n526) );
  NAND2_X1 U583 ( .A1(n526), .A2(n519), .ZN(n520) );
  XNOR2_X1 U584 ( .A(n521), .B(n520), .ZN(G1336GAT) );
  NAND2_X1 U585 ( .A1(n526), .A2(n522), .ZN(n523) );
  XNOR2_X1 U586 ( .A(n523), .B(KEYINPUT110), .ZN(n524) );
  XNOR2_X1 U587 ( .A(G92GAT), .B(n524), .ZN(G1337GAT) );
  NAND2_X1 U588 ( .A1(n532), .A2(n526), .ZN(n525) );
  XNOR2_X1 U589 ( .A(n525), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U590 ( .A(KEYINPUT44), .B(KEYINPUT111), .Z(n528) );
  NAND2_X1 U591 ( .A1(n526), .A2(n534), .ZN(n527) );
  XNOR2_X1 U592 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U593 ( .A(G106GAT), .B(n529), .ZN(G1339GAT) );
  NOR2_X1 U594 ( .A1(n531), .A2(n530), .ZN(n548) );
  NAND2_X1 U595 ( .A1(n548), .A2(n532), .ZN(n533) );
  NOR2_X1 U596 ( .A1(n534), .A2(n533), .ZN(n537) );
  NAND2_X1 U597 ( .A1(n537), .A2(n535), .ZN(n536) );
  XNOR2_X1 U598 ( .A(n536), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U599 ( .A(G120GAT), .B(KEYINPUT49), .Z(n539) );
  INV_X1 U600 ( .A(n537), .ZN(n543) );
  OR2_X1 U601 ( .A1(n543), .A2(n564), .ZN(n538) );
  XNOR2_X1 U602 ( .A(n539), .B(n538), .ZN(G1341GAT) );
  NOR2_X1 U603 ( .A1(n567), .A2(n543), .ZN(n541) );
  XNOR2_X1 U604 ( .A(KEYINPUT50), .B(KEYINPUT115), .ZN(n540) );
  XNOR2_X1 U605 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U606 ( .A(G127GAT), .B(n542), .ZN(G1342GAT) );
  NOR2_X1 U607 ( .A1(n543), .A2(n557), .ZN(n547) );
  XOR2_X1 U608 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n545) );
  XNOR2_X1 U609 ( .A(G134GAT), .B(KEYINPUT116), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U611 ( .A(n547), .B(n546), .ZN(G1343GAT) );
  NAND2_X1 U612 ( .A1(n570), .A2(n548), .ZN(n549) );
  XNOR2_X1 U613 ( .A(n549), .B(KEYINPUT118), .ZN(n556) );
  NOR2_X1 U614 ( .A1(n556), .A2(n572), .ZN(n551) );
  XNOR2_X1 U615 ( .A(G141GAT), .B(KEYINPUT119), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n551), .B(n550), .ZN(G1344GAT) );
  NOR2_X1 U617 ( .A1(n556), .A2(n564), .ZN(n553) );
  XNOR2_X1 U618 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U620 ( .A(G148GAT), .B(n554), .ZN(G1345GAT) );
  NOR2_X1 U621 ( .A1(n556), .A2(n580), .ZN(n555) );
  XOR2_X1 U622 ( .A(G155GAT), .B(n555), .Z(G1346GAT) );
  NOR2_X1 U623 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U624 ( .A(G162GAT), .B(n558), .Z(G1347GAT) );
  NOR2_X1 U625 ( .A1(n572), .A2(n559), .ZN(n561) );
  XNOR2_X1 U626 ( .A(G169GAT), .B(KEYINPUT121), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(G1348GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT122), .B(KEYINPUT56), .Z(n563) );
  XNOR2_X1 U629 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(n566) );
  NOR2_X1 U631 ( .A1(n564), .A2(n559), .ZN(n565) );
  XOR2_X1 U632 ( .A(n566), .B(n565), .Z(G1349GAT) );
  NOR2_X1 U633 ( .A1(n567), .A2(n559), .ZN(n569) );
  XNOR2_X1 U634 ( .A(G183GAT), .B(KEYINPUT123), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(G1350GAT) );
  NAND2_X1 U636 ( .A1(n571), .A2(n570), .ZN(n583) );
  NOR2_X1 U637 ( .A1(n572), .A2(n583), .ZN(n574) );
  XNOR2_X1 U638 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(n575), .ZN(G1352GAT) );
  NOR2_X1 U641 ( .A1(n576), .A2(n583), .ZN(n578) );
  XNOR2_X1 U642 ( .A(KEYINPUT125), .B(KEYINPUT61), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(n579) );
  XOR2_X1 U644 ( .A(G204GAT), .B(n579), .Z(G1353GAT) );
  NOR2_X1 U645 ( .A1(n580), .A2(n583), .ZN(n581) );
  XOR2_X1 U646 ( .A(KEYINPUT126), .B(n581), .Z(n582) );
  XNOR2_X1 U647 ( .A(G211GAT), .B(n582), .ZN(G1354GAT) );
  NOR2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n586) );
  XNOR2_X1 U649 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(n587) );
  XNOR2_X1 U651 ( .A(G218GAT), .B(n587), .ZN(G1355GAT) );
endmodule

