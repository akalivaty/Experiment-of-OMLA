

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587;

  XNOR2_X1 U325 ( .A(n305), .B(n304), .ZN(n307) );
  XNOR2_X1 U326 ( .A(n420), .B(n303), .ZN(n304) );
  XNOR2_X1 U327 ( .A(n395), .B(n394), .ZN(n465) );
  XNOR2_X1 U328 ( .A(n455), .B(KEYINPUT45), .ZN(n456) );
  XNOR2_X1 U329 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U330 ( .A(n467), .B(KEYINPUT47), .ZN(n468) );
  XNOR2_X1 U331 ( .A(n344), .B(n316), .ZN(n299) );
  INV_X1 U332 ( .A(KEYINPUT32), .ZN(n424) );
  XNOR2_X1 U333 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U334 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U335 ( .A(n449), .B(n393), .ZN(n394) );
  INV_X1 U336 ( .A(G169GAT), .ZN(n295) );
  XNOR2_X1 U337 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U338 ( .A(n296), .B(n295), .ZN(n344) );
  XOR2_X1 U339 ( .A(n449), .B(n448), .Z(n571) );
  INV_X1 U340 ( .A(G36GAT), .ZN(n452) );
  XNOR2_X1 U341 ( .A(n486), .B(KEYINPUT58), .ZN(n487) );
  XNOR2_X1 U342 ( .A(n452), .B(KEYINPUT102), .ZN(n453) );
  XNOR2_X1 U343 ( .A(n488), .B(n487), .ZN(G1351GAT) );
  XNOR2_X1 U344 ( .A(n454), .B(n453), .ZN(G1329GAT) );
  XOR2_X1 U345 ( .A(G36GAT), .B(G190GAT), .Z(n377) );
  XOR2_X1 U346 ( .A(KEYINPUT95), .B(G204GAT), .Z(n300) );
  XOR2_X1 U347 ( .A(KEYINPUT85), .B(KEYINPUT17), .Z(n294) );
  XNOR2_X1 U348 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n293) );
  XNOR2_X1 U349 ( .A(n294), .B(n293), .ZN(n296) );
  XOR2_X1 U350 ( .A(KEYINPUT88), .B(KEYINPUT21), .Z(n298) );
  XNOR2_X1 U351 ( .A(G197GAT), .B(G218GAT), .ZN(n297) );
  XNOR2_X1 U352 ( .A(n298), .B(n297), .ZN(n316) );
  XNOR2_X1 U353 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U354 ( .A(n377), .B(n301), .Z(n305) );
  XNOR2_X1 U355 ( .A(G176GAT), .B(G92GAT), .ZN(n302) );
  XNOR2_X1 U356 ( .A(n302), .B(G64GAT), .ZN(n420) );
  NAND2_X1 U357 ( .A1(G226GAT), .A2(G233GAT), .ZN(n303) );
  XOR2_X1 U358 ( .A(G8GAT), .B(G183GAT), .Z(n306) );
  XOR2_X1 U359 ( .A(G211GAT), .B(n306), .Z(n406) );
  XOR2_X1 U360 ( .A(n307), .B(n406), .Z(n308) );
  INV_X1 U361 ( .A(n308), .ZN(n346) );
  XNOR2_X1 U362 ( .A(KEYINPUT27), .B(n346), .ZN(n373) );
  XOR2_X1 U363 ( .A(G211GAT), .B(KEYINPUT22), .Z(n310) );
  XNOR2_X1 U364 ( .A(KEYINPUT90), .B(KEYINPUT24), .ZN(n309) );
  XNOR2_X1 U365 ( .A(n310), .B(n309), .ZN(n312) );
  XOR2_X1 U366 ( .A(G50GAT), .B(G22GAT), .Z(n311) );
  XNOR2_X1 U367 ( .A(n312), .B(n311), .ZN(n320) );
  XNOR2_X1 U368 ( .A(KEYINPUT87), .B(G155GAT), .ZN(n313) );
  XNOR2_X1 U369 ( .A(n313), .B(G148GAT), .ZN(n314) );
  XOR2_X1 U370 ( .A(n314), .B(KEYINPUT23), .Z(n318) );
  XNOR2_X1 U371 ( .A(G106GAT), .B(G78GAT), .ZN(n315) );
  XNOR2_X1 U372 ( .A(n315), .B(G204GAT), .ZN(n415) );
  XNOR2_X1 U373 ( .A(n316), .B(n415), .ZN(n317) );
  XNOR2_X1 U374 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U375 ( .A(n320), .B(n319), .ZN(n322) );
  NAND2_X1 U376 ( .A1(G228GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U377 ( .A(n322), .B(n321), .ZN(n326) );
  XOR2_X1 U378 ( .A(KEYINPUT2), .B(G162GAT), .Z(n324) );
  XNOR2_X1 U379 ( .A(KEYINPUT89), .B(KEYINPUT3), .ZN(n323) );
  XNOR2_X1 U380 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U381 ( .A(G141GAT), .B(n325), .Z(n357) );
  XOR2_X1 U382 ( .A(n326), .B(n357), .Z(n476) );
  XOR2_X1 U383 ( .A(G71GAT), .B(G127GAT), .Z(n328) );
  XNOR2_X1 U384 ( .A(G15GAT), .B(G176GAT), .ZN(n327) );
  XNOR2_X1 U385 ( .A(n328), .B(n327), .ZN(n342) );
  XOR2_X1 U386 ( .A(G120GAT), .B(KEYINPUT66), .Z(n330) );
  XNOR2_X1 U387 ( .A(G43GAT), .B(G190GAT), .ZN(n329) );
  XNOR2_X1 U388 ( .A(n330), .B(n329), .ZN(n334) );
  XOR2_X1 U389 ( .A(G183GAT), .B(KEYINPUT84), .Z(n332) );
  XNOR2_X1 U390 ( .A(KEYINPUT20), .B(KEYINPUT86), .ZN(n331) );
  XNOR2_X1 U391 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U392 ( .A(n334), .B(n333), .Z(n340) );
  XNOR2_X1 U393 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n335) );
  XNOR2_X1 U394 ( .A(n335), .B(KEYINPUT83), .ZN(n358) );
  XOR2_X1 U395 ( .A(G134GAT), .B(n358), .Z(n337) );
  NAND2_X1 U396 ( .A1(G227GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U397 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U398 ( .A(G99GAT), .B(n338), .ZN(n339) );
  XNOR2_X1 U399 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U400 ( .A(n342), .B(n341), .Z(n343) );
  XOR2_X1 U401 ( .A(n344), .B(n343), .Z(n536) );
  NOR2_X1 U402 ( .A1(n476), .A2(n536), .ZN(n345) );
  XNOR2_X1 U403 ( .A(n345), .B(KEYINPUT26), .ZN(n569) );
  NAND2_X1 U404 ( .A1(n373), .A2(n569), .ZN(n549) );
  XNOR2_X1 U405 ( .A(n549), .B(KEYINPUT96), .ZN(n350) );
  NAND2_X1 U406 ( .A1(n536), .A2(n346), .ZN(n347) );
  NAND2_X1 U407 ( .A1(n476), .A2(n347), .ZN(n348) );
  XOR2_X1 U408 ( .A(KEYINPUT25), .B(n348), .Z(n349) );
  NAND2_X1 U409 ( .A1(n350), .A2(n349), .ZN(n369) );
  XOR2_X1 U410 ( .A(KEYINPUT5), .B(KEYINPUT92), .Z(n352) );
  XNOR2_X1 U411 ( .A(G85GAT), .B(KEYINPUT6), .ZN(n351) );
  XNOR2_X1 U412 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U413 ( .A(KEYINPUT4), .B(KEYINPUT91), .Z(n354) );
  XNOR2_X1 U414 ( .A(KEYINPUT1), .B(G57GAT), .ZN(n353) );
  XNOR2_X1 U415 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U416 ( .A(n356), .B(n355), .Z(n364) );
  INV_X1 U417 ( .A(n357), .ZN(n362) );
  XOR2_X1 U418 ( .A(KEYINPUT93), .B(n358), .Z(n360) );
  NAND2_X1 U419 ( .A1(G225GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U420 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U421 ( .A(n362), .B(n361), .Z(n363) );
  XNOR2_X1 U422 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U423 ( .A(G120GAT), .B(G148GAT), .Z(n423) );
  XOR2_X1 U424 ( .A(n365), .B(n423), .Z(n368) );
  XOR2_X1 U425 ( .A(G29GAT), .B(G134GAT), .Z(n378) );
  XNOR2_X1 U426 ( .A(G1GAT), .B(G127GAT), .ZN(n366) );
  XNOR2_X1 U427 ( .A(n366), .B(G155GAT), .ZN(n407) );
  XNOR2_X1 U428 ( .A(n378), .B(n407), .ZN(n367) );
  XNOR2_X1 U429 ( .A(n368), .B(n367), .ZN(n372) );
  NAND2_X1 U430 ( .A1(n369), .A2(n372), .ZN(n370) );
  XNOR2_X1 U431 ( .A(n370), .B(KEYINPUT97), .ZN(n376) );
  XNOR2_X1 U432 ( .A(n476), .B(KEYINPUT67), .ZN(n371) );
  XOR2_X1 U433 ( .A(n371), .B(KEYINPUT28), .Z(n531) );
  XOR2_X1 U434 ( .A(KEYINPUT94), .B(n372), .Z(n552) );
  AND2_X1 U435 ( .A1(n531), .A2(n552), .ZN(n374) );
  NAND2_X1 U436 ( .A1(n374), .A2(n373), .ZN(n534) );
  NOR2_X1 U437 ( .A1(n534), .A2(n536), .ZN(n375) );
  NOR2_X1 U438 ( .A1(n376), .A2(n375), .ZN(n491) );
  XOR2_X1 U439 ( .A(KEYINPUT78), .B(n377), .Z(n380) );
  XNOR2_X1 U440 ( .A(G218GAT), .B(n378), .ZN(n379) );
  XNOR2_X1 U441 ( .A(n380), .B(n379), .ZN(n385) );
  XNOR2_X1 U442 ( .A(G99GAT), .B(G85GAT), .ZN(n381) );
  XNOR2_X1 U443 ( .A(n381), .B(KEYINPUT75), .ZN(n414) );
  XOR2_X1 U444 ( .A(n414), .B(KEYINPUT11), .Z(n383) );
  NAND2_X1 U445 ( .A1(G232GAT), .A2(G233GAT), .ZN(n382) );
  XNOR2_X1 U446 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U447 ( .A(n385), .B(n384), .ZN(n387) );
  XOR2_X1 U448 ( .A(G162GAT), .B(G106GAT), .Z(n386) );
  XNOR2_X1 U449 ( .A(n387), .B(n386), .ZN(n395) );
  XOR2_X1 U450 ( .A(KEYINPUT73), .B(KEYINPUT7), .Z(n389) );
  XNOR2_X1 U451 ( .A(G50GAT), .B(G43GAT), .ZN(n388) );
  XNOR2_X1 U452 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U453 ( .A(KEYINPUT8), .B(n390), .ZN(n449) );
  XOR2_X1 U454 ( .A(KEYINPUT79), .B(KEYINPUT9), .Z(n392) );
  XNOR2_X1 U455 ( .A(G92GAT), .B(KEYINPUT10), .ZN(n391) );
  XNOR2_X1 U456 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U457 ( .A(KEYINPUT36), .B(KEYINPUT99), .ZN(n396) );
  XNOR2_X1 U458 ( .A(n465), .B(n396), .ZN(n584) );
  NOR2_X1 U459 ( .A1(n491), .A2(n584), .ZN(n412) );
  XOR2_X1 U460 ( .A(KEYINPUT82), .B(KEYINPUT80), .Z(n398) );
  XNOR2_X1 U461 ( .A(G78GAT), .B(G64GAT), .ZN(n397) );
  XNOR2_X1 U462 ( .A(n398), .B(n397), .ZN(n411) );
  XNOR2_X1 U463 ( .A(G71GAT), .B(G57GAT), .ZN(n399) );
  XNOR2_X1 U464 ( .A(n399), .B(KEYINPUT13), .ZN(n419) );
  XOR2_X1 U465 ( .A(G15GAT), .B(G22GAT), .Z(n441) );
  XOR2_X1 U466 ( .A(n419), .B(n441), .Z(n401) );
  NAND2_X1 U467 ( .A1(G231GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U468 ( .A(n401), .B(n400), .ZN(n405) );
  XOR2_X1 U469 ( .A(KEYINPUT15), .B(KEYINPUT81), .Z(n403) );
  XNOR2_X1 U470 ( .A(KEYINPUT12), .B(KEYINPUT14), .ZN(n402) );
  XNOR2_X1 U471 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U472 ( .A(n405), .B(n404), .Z(n409) );
  XNOR2_X1 U473 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U474 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U475 ( .A(n411), .B(n410), .ZN(n580) );
  NAND2_X1 U476 ( .A1(n412), .A2(n580), .ZN(n413) );
  XNOR2_X1 U477 ( .A(KEYINPUT37), .B(n413), .ZN(n522) );
  XNOR2_X1 U478 ( .A(n415), .B(n414), .ZN(n429) );
  XOR2_X1 U479 ( .A(KEYINPUT76), .B(KEYINPUT33), .Z(n417) );
  NAND2_X1 U480 ( .A1(G230GAT), .A2(G233GAT), .ZN(n416) );
  XNOR2_X1 U481 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U482 ( .A(n418), .B(KEYINPUT31), .Z(n422) );
  XNOR2_X1 U483 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U484 ( .A(n422), .B(n421), .ZN(n427) );
  XNOR2_X1 U485 ( .A(n423), .B(KEYINPUT77), .ZN(n425) );
  XNOR2_X1 U486 ( .A(n429), .B(n428), .ZN(n462) );
  XOR2_X1 U487 ( .A(G8GAT), .B(G1GAT), .Z(n431) );
  XNOR2_X1 U488 ( .A(G141GAT), .B(G197GAT), .ZN(n430) );
  XNOR2_X1 U489 ( .A(n431), .B(n430), .ZN(n435) );
  XOR2_X1 U490 ( .A(KEYINPUT68), .B(KEYINPUT29), .Z(n433) );
  XNOR2_X1 U491 ( .A(KEYINPUT69), .B(KEYINPUT30), .ZN(n432) );
  XNOR2_X1 U492 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U493 ( .A(n435), .B(n434), .Z(n447) );
  XOR2_X1 U494 ( .A(KEYINPUT72), .B(KEYINPUT71), .Z(n437) );
  XNOR2_X1 U495 ( .A(KEYINPUT70), .B(KEYINPUT74), .ZN(n436) );
  XNOR2_X1 U496 ( .A(n437), .B(n436), .ZN(n445) );
  XOR2_X1 U497 ( .A(G113GAT), .B(G36GAT), .Z(n439) );
  XNOR2_X1 U498 ( .A(G169GAT), .B(G29GAT), .ZN(n438) );
  XNOR2_X1 U499 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U500 ( .A(n441), .B(n440), .Z(n443) );
  NAND2_X1 U501 ( .A1(G229GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U502 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U503 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U504 ( .A(n447), .B(n446), .ZN(n448) );
  NOR2_X1 U505 ( .A1(n462), .A2(n571), .ZN(n492) );
  NAND2_X1 U506 ( .A1(n522), .A2(n492), .ZN(n451) );
  XNOR2_X1 U507 ( .A(KEYINPUT100), .B(KEYINPUT38), .ZN(n450) );
  XNOR2_X1 U508 ( .A(n451), .B(n450), .ZN(n507) );
  NOR2_X1 U509 ( .A1(n507), .A2(n308), .ZN(n454) );
  INV_X1 U510 ( .A(n571), .ZN(n509) );
  NOR2_X1 U511 ( .A1(n584), .A2(n580), .ZN(n457) );
  INV_X1 U512 ( .A(KEYINPUT112), .ZN(n455) );
  NOR2_X1 U513 ( .A1(n462), .A2(n458), .ZN(n459) );
  XNOR2_X1 U514 ( .A(n459), .B(KEYINPUT113), .ZN(n460) );
  NOR2_X1 U515 ( .A1(n509), .A2(n460), .ZN(n471) );
  XNOR2_X1 U516 ( .A(KEYINPUT109), .B(n580), .ZN(n565) );
  XNOR2_X1 U517 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n461) );
  XNOR2_X1 U518 ( .A(n462), .B(n461), .ZN(n557) );
  NOR2_X1 U519 ( .A1(n557), .A2(n571), .ZN(n463) );
  XNOR2_X1 U520 ( .A(n463), .B(KEYINPUT46), .ZN(n464) );
  NOR2_X1 U521 ( .A1(n565), .A2(n464), .ZN(n466) );
  INV_X1 U522 ( .A(n465), .ZN(n562) );
  NAND2_X1 U523 ( .A1(n466), .A2(n562), .ZN(n469) );
  XOR2_X1 U524 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n467) );
  NOR2_X1 U525 ( .A1(n471), .A2(n470), .ZN(n472) );
  XNOR2_X1 U526 ( .A(KEYINPUT48), .B(n472), .ZN(n550) );
  NOR2_X1 U527 ( .A1(n308), .A2(n550), .ZN(n473) );
  XNOR2_X1 U528 ( .A(n473), .B(KEYINPUT54), .ZN(n474) );
  INV_X1 U529 ( .A(n552), .ZN(n523) );
  NAND2_X1 U530 ( .A1(n474), .A2(n523), .ZN(n475) );
  XNOR2_X1 U531 ( .A(n475), .B(KEYINPUT65), .ZN(n570) );
  NAND2_X1 U532 ( .A1(n570), .A2(n476), .ZN(n478) );
  XOR2_X1 U533 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n477) );
  XNOR2_X1 U534 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U535 ( .A(n479), .B(KEYINPUT55), .ZN(n480) );
  NAND2_X1 U536 ( .A1(n480), .A2(n536), .ZN(n564) );
  NOR2_X1 U537 ( .A1(n571), .A2(n564), .ZN(n482) );
  XNOR2_X1 U538 ( .A(G169GAT), .B(KEYINPUT121), .ZN(n481) );
  XNOR2_X1 U539 ( .A(n482), .B(n481), .ZN(G1348GAT) );
  NOR2_X1 U540 ( .A1(n557), .A2(n564), .ZN(n485) );
  XNOR2_X1 U541 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n483) );
  XNOR2_X1 U542 ( .A(n483), .B(G176GAT), .ZN(n484) );
  XNOR2_X1 U543 ( .A(n485), .B(n484), .ZN(G1349GAT) );
  NOR2_X1 U544 ( .A1(n562), .A2(n564), .ZN(n488) );
  INV_X1 U545 ( .A(G190GAT), .ZN(n486) );
  NOR2_X1 U546 ( .A1(n465), .A2(n580), .ZN(n489) );
  XOR2_X1 U547 ( .A(KEYINPUT16), .B(n489), .Z(n490) );
  NOR2_X1 U548 ( .A1(n491), .A2(n490), .ZN(n510) );
  NAND2_X1 U549 ( .A1(n492), .A2(n510), .ZN(n499) );
  NOR2_X1 U550 ( .A1(n523), .A2(n499), .ZN(n493) );
  XOR2_X1 U551 ( .A(G1GAT), .B(n493), .Z(n494) );
  XNOR2_X1 U552 ( .A(KEYINPUT34), .B(n494), .ZN(G1324GAT) );
  NOR2_X1 U553 ( .A1(n308), .A2(n499), .ZN(n495) );
  XOR2_X1 U554 ( .A(G8GAT), .B(n495), .Z(G1325GAT) );
  INV_X1 U555 ( .A(n536), .ZN(n528) );
  NOR2_X1 U556 ( .A1(n528), .A2(n499), .ZN(n497) );
  XNOR2_X1 U557 ( .A(KEYINPUT35), .B(KEYINPUT98), .ZN(n496) );
  XNOR2_X1 U558 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U559 ( .A(G15GAT), .B(n498), .ZN(G1326GAT) );
  NOR2_X1 U560 ( .A1(n531), .A2(n499), .ZN(n500) );
  XOR2_X1 U561 ( .A(G22GAT), .B(n500), .Z(G1327GAT) );
  NOR2_X1 U562 ( .A1(n523), .A2(n507), .ZN(n502) );
  XNOR2_X1 U563 ( .A(KEYINPUT39), .B(KEYINPUT101), .ZN(n501) );
  XNOR2_X1 U564 ( .A(n502), .B(n501), .ZN(n503) );
  XOR2_X1 U565 ( .A(G29GAT), .B(n503), .Z(G1328GAT) );
  NOR2_X1 U566 ( .A1(n528), .A2(n507), .ZN(n505) );
  XNOR2_X1 U567 ( .A(KEYINPUT40), .B(KEYINPUT103), .ZN(n504) );
  XNOR2_X1 U568 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U569 ( .A(G43GAT), .B(n506), .ZN(G1330GAT) );
  NOR2_X1 U570 ( .A1(n531), .A2(n507), .ZN(n508) );
  XOR2_X1 U571 ( .A(G50GAT), .B(n508), .Z(G1331GAT) );
  NOR2_X1 U572 ( .A1(n509), .A2(n557), .ZN(n521) );
  NAND2_X1 U573 ( .A1(n510), .A2(n521), .ZN(n511) );
  XNOR2_X1 U574 ( .A(n511), .B(KEYINPUT104), .ZN(n517) );
  NOR2_X1 U575 ( .A1(n517), .A2(n523), .ZN(n512) );
  XOR2_X1 U576 ( .A(KEYINPUT42), .B(n512), .Z(n513) );
  XNOR2_X1 U577 ( .A(G57GAT), .B(n513), .ZN(G1332GAT) );
  NOR2_X1 U578 ( .A1(n517), .A2(n308), .ZN(n515) );
  XNOR2_X1 U579 ( .A(G64GAT), .B(KEYINPUT105), .ZN(n514) );
  XNOR2_X1 U580 ( .A(n515), .B(n514), .ZN(G1333GAT) );
  NOR2_X1 U581 ( .A1(n517), .A2(n528), .ZN(n516) );
  XOR2_X1 U582 ( .A(G71GAT), .B(n516), .Z(G1334GAT) );
  NOR2_X1 U583 ( .A1(n517), .A2(n531), .ZN(n519) );
  XNOR2_X1 U584 ( .A(KEYINPUT106), .B(KEYINPUT43), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U586 ( .A(G78GAT), .B(n520), .ZN(G1335GAT) );
  NAND2_X1 U587 ( .A1(n522), .A2(n521), .ZN(n530) );
  NOR2_X1 U588 ( .A1(n523), .A2(n530), .ZN(n525) );
  XNOR2_X1 U589 ( .A(KEYINPUT107), .B(KEYINPUT108), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U591 ( .A(G85GAT), .B(n526), .ZN(G1336GAT) );
  NOR2_X1 U592 ( .A1(n308), .A2(n530), .ZN(n527) );
  XOR2_X1 U593 ( .A(G92GAT), .B(n527), .Z(G1337GAT) );
  NOR2_X1 U594 ( .A1(n528), .A2(n530), .ZN(n529) );
  XOR2_X1 U595 ( .A(G99GAT), .B(n529), .Z(G1338GAT) );
  NOR2_X1 U596 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U597 ( .A(KEYINPUT44), .B(n532), .Z(n533) );
  XNOR2_X1 U598 ( .A(G106GAT), .B(n533), .ZN(G1339GAT) );
  NOR2_X1 U599 ( .A1(n550), .A2(n534), .ZN(n535) );
  NAND2_X1 U600 ( .A1(n536), .A2(n535), .ZN(n541) );
  NOR2_X1 U601 ( .A1(n571), .A2(n541), .ZN(n537) );
  XOR2_X1 U602 ( .A(G113GAT), .B(n537), .Z(G1340GAT) );
  NOR2_X1 U603 ( .A1(n557), .A2(n541), .ZN(n539) );
  XNOR2_X1 U604 ( .A(KEYINPUT114), .B(KEYINPUT49), .ZN(n538) );
  XNOR2_X1 U605 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U606 ( .A(G120GAT), .B(n540), .ZN(G1341GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n543) );
  INV_X1 U608 ( .A(n541), .ZN(n545) );
  NAND2_X1 U609 ( .A1(n545), .A2(n565), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U611 ( .A(G127GAT), .B(n544), .ZN(G1342GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT51), .B(KEYINPUT116), .Z(n547) );
  NAND2_X1 U613 ( .A1(n545), .A2(n465), .ZN(n546) );
  XNOR2_X1 U614 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U615 ( .A(G134GAT), .B(n548), .ZN(G1343GAT) );
  NOR2_X1 U616 ( .A1(n550), .A2(n549), .ZN(n551) );
  NAND2_X1 U617 ( .A1(n552), .A2(n551), .ZN(n561) );
  NOR2_X1 U618 ( .A1(n571), .A2(n561), .ZN(n554) );
  XNOR2_X1 U619 ( .A(G141GAT), .B(KEYINPUT117), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n554), .B(n553), .ZN(G1344GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT118), .B(KEYINPUT52), .Z(n556) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(n559) );
  NOR2_X1 U624 ( .A1(n557), .A2(n561), .ZN(n558) );
  XOR2_X1 U625 ( .A(n559), .B(n558), .Z(G1345GAT) );
  NOR2_X1 U626 ( .A1(n580), .A2(n561), .ZN(n560) );
  XOR2_X1 U627 ( .A(G155GAT), .B(n560), .Z(G1346GAT) );
  NOR2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U629 ( .A(G162GAT), .B(n563), .Z(G1347GAT) );
  INV_X1 U630 ( .A(n564), .ZN(n566) );
  NAND2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U632 ( .A(n567), .B(KEYINPUT122), .ZN(n568) );
  XNOR2_X1 U633 ( .A(G183GAT), .B(n568), .ZN(G1350GAT) );
  NAND2_X1 U634 ( .A1(n570), .A2(n569), .ZN(n583) );
  NOR2_X1 U635 ( .A1(n571), .A2(n583), .ZN(n575) );
  XOR2_X1 U636 ( .A(KEYINPUT59), .B(KEYINPUT123), .Z(n573) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n575), .B(n574), .ZN(G1352GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT61), .B(KEYINPUT124), .Z(n578) );
  INV_X1 U641 ( .A(n583), .ZN(n576) );
  NAND2_X1 U642 ( .A1(n576), .A2(n462), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(G204GAT), .B(n579), .ZN(G1353GAT) );
  NOR2_X1 U645 ( .A1(n580), .A2(n583), .ZN(n582) );
  XNOR2_X1 U646 ( .A(G211GAT), .B(KEYINPUT125), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1354GAT) );
  NOR2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n586) );
  XNOR2_X1 U649 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(n587) );
  XOR2_X1 U651 ( .A(G218GAT), .B(n587), .Z(G1355GAT) );
endmodule

