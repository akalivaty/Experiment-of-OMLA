//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 1 1 0 1 1 1 0 0 1 0 1 1 0 1 1 0 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 0 0 0 1 1 0 1 0 0 0 1 0 0 1 1 0 0 1 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:19 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1243;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT0), .Z(new_n212));
  NAND2_X1  g0012(.A1(G107), .A2(G264), .ZN(new_n213));
  INV_X1    g0013(.A(G77), .ZN(new_n214));
  INV_X1    g0014(.A(G244), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT64), .Z(new_n218));
  AOI211_X1 g0018(.A(new_n216), .B(new_n218), .C1(G68), .C2(G238), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G87), .A2(G250), .ZN(new_n220));
  INV_X1    g0020(.A(G232), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n219), .B(new_n220), .C1(new_n201), .C2(new_n221), .ZN(new_n222));
  AND2_X1   g0022(.A1(G97), .A2(G257), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n209), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT1), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n203), .A2(G50), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n212), .B(new_n225), .C1(new_n228), .C2(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G250), .B(G257), .Z(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(new_n205), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT65), .B(G87), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G68), .B(G77), .Z(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  NAND3_X1  g0047(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(new_n226), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(KEYINPUT8), .B(G58), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n252), .A2(G20), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G150), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G20), .A2(G33), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  OAI22_X1  g0057(.A1(new_n251), .A2(new_n254), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  XNOR2_X1  g0058(.A(new_n258), .B(KEYINPUT67), .ZN(new_n259));
  OAI21_X1  g0059(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n250), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G50), .ZN(new_n262));
  INV_X1    g0062(.A(G1), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n263), .A2(G13), .A3(G20), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n261), .B1(new_n262), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n263), .A2(G20), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n250), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n266), .B1(new_n262), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT9), .ZN(new_n270));
  OR2_X1    g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n226), .B1(G33), .B2(G41), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G1698), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT66), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT66), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G1698), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  AOI22_X1  g0078(.A1(new_n278), .A2(G222), .B1(G223), .B2(G1698), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT3), .B(G33), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n273), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n281), .B1(G77), .B2(new_n280), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n263), .B1(G41), .B2(G45), .ZN(new_n283));
  INV_X1    g0083(.A(G274), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n273), .A2(new_n283), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G226), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n282), .A2(new_n286), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G200), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n269), .A2(new_n270), .ZN(new_n292));
  INV_X1    g0092(.A(G190), .ZN(new_n293));
  OR2_X1    g0093(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  NAND4_X1  g0094(.A1(new_n271), .A2(new_n291), .A3(new_n292), .A4(new_n294), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n295), .B(KEYINPUT10), .ZN(new_n296));
  INV_X1    g0096(.A(G169), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n290), .A2(new_n297), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n269), .B(new_n298), .C1(G179), .C2(new_n290), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(G33), .A2(G97), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT68), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(KEYINPUT68), .A2(G33), .A3(G97), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  AOI22_X1  g0106(.A1(new_n278), .A2(G226), .B1(G232), .B2(G1698), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT3), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G33), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n306), .B1(new_n307), .B2(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n285), .B1(new_n312), .B2(new_n272), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n288), .A2(G238), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT13), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT13), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n313), .A2(new_n317), .A3(new_n314), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n319), .A2(new_n293), .ZN(new_n320));
  INV_X1    g0120(.A(G200), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n321), .B1(new_n316), .B2(new_n318), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n253), .A2(G77), .B1(G20), .B2(new_n202), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n323), .B1(new_n262), .B2(new_n257), .ZN(new_n324));
  AOI21_X1  g0124(.A(KEYINPUT11), .B1(new_n324), .B2(new_n249), .ZN(new_n325));
  INV_X1    g0125(.A(new_n268), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n325), .B1(G68), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n324), .A2(KEYINPUT11), .A3(new_n249), .ZN(new_n328));
  OAI21_X1  g0128(.A(KEYINPUT69), .B1(new_n264), .B2(G68), .ZN(new_n329));
  XOR2_X1   g0129(.A(new_n329), .B(KEYINPUT12), .Z(new_n330));
  NAND3_X1  g0130(.A1(new_n327), .A2(new_n328), .A3(new_n330), .ZN(new_n331));
  NOR3_X1   g0131(.A1(new_n320), .A2(new_n322), .A3(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n318), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n317), .B1(new_n313), .B2(new_n314), .ZN(new_n334));
  OAI21_X1  g0134(.A(G169), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(KEYINPUT14), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT14), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n319), .A2(new_n337), .A3(G169), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n316), .A2(G179), .A3(new_n318), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n336), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n332), .B1(new_n340), .B2(new_n331), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n278), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n343));
  INV_X1    g0143(.A(G87), .ZN(new_n344));
  OAI22_X1  g0144(.A1(new_n343), .A2(new_n311), .B1(new_n252), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(new_n272), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n288), .A2(G232), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n346), .A2(new_n286), .A3(new_n347), .ZN(new_n348));
  OR2_X1    g0148(.A1(new_n348), .A2(new_n293), .ZN(new_n349));
  NAND2_X1  g0149(.A1(G58), .A2(G68), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n227), .B1(new_n203), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT7), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n352), .B1(new_n280), .B2(G20), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n311), .A2(KEYINPUT7), .A3(new_n227), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n351), .B1(new_n355), .B2(G68), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n256), .A2(G159), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT16), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n356), .A2(KEYINPUT16), .A3(new_n357), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n360), .A2(new_n249), .A3(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n251), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n267), .ZN(new_n364));
  XOR2_X1   g0164(.A(new_n364), .B(KEYINPUT70), .Z(new_n365));
  NOR2_X1   g0165(.A1(new_n265), .A2(new_n249), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n365), .A2(new_n366), .B1(new_n265), .B2(new_n251), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n348), .A2(G200), .ZN(new_n368));
  AND4_X1   g0168(.A1(new_n349), .A2(new_n362), .A3(new_n367), .A4(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT72), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT17), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n349), .A2(new_n362), .A3(new_n367), .A4(new_n368), .ZN(new_n373));
  OAI21_X1  g0173(.A(KEYINPUT17), .B1(new_n373), .B2(KEYINPUT72), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n348), .A2(G169), .ZN(new_n376));
  INV_X1    g0176(.A(G179), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n376), .B1(new_n377), .B2(new_n348), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT71), .ZN(new_n379));
  AND3_X1   g0179(.A1(new_n362), .A2(new_n379), .A3(new_n367), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n379), .B1(new_n362), .B2(new_n367), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n378), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(KEYINPUT18), .ZN(new_n383));
  INV_X1    g0183(.A(G238), .ZN(new_n384));
  XNOR2_X1  g0184(.A(KEYINPUT66), .B(G1698), .ZN(new_n385));
  OAI221_X1 g0185(.A(new_n280), .B1(new_n384), .B2(new_n274), .C1(new_n385), .C2(new_n221), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n386), .B(new_n272), .C1(G107), .C2(new_n280), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n387), .B(new_n286), .C1(new_n215), .C2(new_n287), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(G200), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(new_n293), .B2(new_n388), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n363), .A2(new_n256), .B1(G20), .B2(G77), .ZN(new_n391));
  XOR2_X1   g0191(.A(KEYINPUT15), .B(G87), .Z(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n391), .B1(new_n254), .B2(new_n393), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n394), .A2(new_n249), .B1(new_n214), .B2(new_n265), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(new_n214), .B2(new_n268), .ZN(new_n396));
  OR2_X1    g0196(.A1(new_n390), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n388), .A2(new_n297), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n396), .B(new_n398), .C1(G179), .C2(new_n388), .ZN(new_n399));
  AND2_X1   g0199(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT18), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n401), .B(new_n378), .C1(new_n380), .C2(new_n381), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n375), .A2(new_n383), .A3(new_n400), .A4(new_n402), .ZN(new_n403));
  NOR3_X1   g0203(.A1(new_n300), .A2(new_n342), .A3(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n278), .A2(new_n280), .A3(G244), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT4), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n308), .A2(new_n310), .A3(G250), .A4(G1698), .ZN(new_n408));
  NAND2_X1  g0208(.A1(G33), .A2(G283), .ZN(new_n409));
  AND2_X1   g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n215), .B1(new_n275), .B2(new_n277), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n411), .A2(KEYINPUT4), .A3(new_n280), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n407), .A2(new_n410), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n272), .ZN(new_n414));
  INV_X1    g0214(.A(G41), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n263), .B(G45), .C1(new_n415), .C2(KEYINPUT5), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(KEYINPUT73), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT5), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(G41), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT73), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n419), .A2(new_n420), .A3(new_n263), .A4(G45), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n418), .A2(G41), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n422), .A2(new_n284), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n273), .A2(new_n417), .A3(new_n421), .A4(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(KEYINPUT74), .ZN(new_n425));
  NOR3_X1   g0225(.A1(new_n272), .A2(new_n284), .A3(new_n422), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT74), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n426), .A2(new_n427), .A3(new_n417), .A4(new_n421), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n416), .A2(new_n422), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n430), .A2(new_n272), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(G257), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n414), .A2(new_n429), .A3(G190), .A4(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT75), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n264), .A2(G97), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n263), .A2(G33), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n264), .A2(new_n437), .A3(new_n226), .A4(new_n248), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n438), .A2(new_n205), .ZN(new_n439));
  NOR3_X1   g0239(.A1(new_n280), .A2(new_n352), .A3(G20), .ZN(new_n440));
  AOI21_X1  g0240(.A(KEYINPUT7), .B1(new_n311), .B2(new_n227), .ZN(new_n441));
  OAI21_X1  g0241(.A(G107), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n256), .A2(G77), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n206), .A2(KEYINPUT6), .A3(G97), .ZN(new_n444));
  XOR2_X1   g0244(.A(G97), .B(G107), .Z(new_n445));
  OAI21_X1  g0245(.A(new_n444), .B1(new_n445), .B2(KEYINPUT6), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(G20), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n442), .A2(new_n443), .A3(new_n447), .ZN(new_n448));
  AOI211_X1 g0248(.A(new_n436), .B(new_n439), .C1(new_n448), .C2(new_n249), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n429), .A2(new_n432), .ZN(new_n450));
  AND3_X1   g0250(.A1(new_n411), .A2(KEYINPUT4), .A3(new_n280), .ZN(new_n451));
  AOI21_X1  g0251(.A(KEYINPUT4), .B1(new_n411), .B2(new_n280), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n273), .B1(new_n453), .B2(new_n410), .ZN(new_n454));
  OAI21_X1  g0254(.A(G200), .B1(new_n450), .B2(new_n454), .ZN(new_n455));
  AOI22_X1  g0255(.A1(new_n425), .A2(new_n428), .B1(G257), .B2(new_n431), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n456), .A2(new_n414), .A3(KEYINPUT75), .A4(G190), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n435), .A2(new_n449), .A3(new_n455), .A4(new_n457), .ZN(new_n458));
  OR3_X1    g0258(.A1(new_n264), .A2(KEYINPUT25), .A3(G107), .ZN(new_n459));
  OAI21_X1  g0259(.A(KEYINPUT25), .B1(new_n264), .B2(G107), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n459), .B(new_n460), .C1(new_n206), .C2(new_n438), .ZN(new_n461));
  XNOR2_X1  g0261(.A(new_n461), .B(KEYINPUT82), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n308), .A2(new_n310), .A3(new_n227), .A4(G87), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT80), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n464), .A2(KEYINPUT22), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT23), .ZN(new_n466));
  OAI21_X1  g0266(.A(KEYINPUT81), .B1(new_n227), .B2(G107), .ZN(new_n467));
  AOI22_X1  g0267(.A1(new_n463), .A2(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OR2_X1    g0268(.A1(new_n467), .A2(new_n466), .ZN(new_n469));
  AND2_X1   g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(G116), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n252), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n227), .ZN(new_n473));
  XOR2_X1   g0273(.A(KEYINPUT80), .B(KEYINPUT22), .Z(new_n474));
  OR2_X1    g0274(.A1(new_n463), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n470), .A2(KEYINPUT24), .A3(new_n473), .A4(new_n475), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n475), .A2(new_n468), .A3(new_n473), .A4(new_n469), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT24), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n476), .A2(new_n249), .A3(new_n479), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n308), .A2(new_n310), .A3(G257), .A4(G1698), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT83), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n280), .A2(KEYINPUT83), .A3(G257), .A4(G1698), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n278), .A2(new_n280), .A3(G250), .ZN(new_n485));
  NAND2_X1  g0285(.A1(G33), .A2(G294), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n483), .A2(new_n484), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n487), .A2(new_n272), .B1(G264), .B2(new_n431), .ZN(new_n488));
  AND3_X1   g0288(.A1(new_n488), .A2(new_n293), .A3(new_n429), .ZN(new_n489));
  AOI21_X1  g0289(.A(G200), .B1(new_n488), .B2(new_n429), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n462), .B(new_n480), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n456), .A2(new_n414), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n297), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n448), .A2(new_n249), .ZN(new_n494));
  INV_X1    g0294(.A(new_n436), .ZN(new_n495));
  INV_X1    g0295(.A(new_n439), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n456), .A2(new_n377), .A3(new_n414), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n493), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n458), .A2(new_n491), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n480), .A2(new_n462), .ZN(new_n501));
  AND2_X1   g0301(.A1(new_n488), .A2(new_n429), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n377), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n488), .A2(new_n429), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n297), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n501), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n500), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n438), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(G116), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n265), .A2(new_n471), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n248), .A2(new_n226), .B1(G20), .B2(new_n471), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n409), .B(new_n227), .C1(G33), .C2(new_n205), .ZN(new_n513));
  AND3_X1   g0313(.A1(new_n512), .A2(KEYINPUT20), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(KEYINPUT20), .B1(new_n512), .B2(new_n513), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n510), .B(new_n511), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  AND2_X1   g0316(.A1(new_n516), .A2(G179), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT77), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n431), .A2(G270), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n278), .A2(G257), .B1(G264), .B2(G1698), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n273), .B1(new_n520), .B2(new_n280), .ZN(new_n521));
  INV_X1    g0321(.A(G303), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n311), .A2(new_n522), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n428), .A2(new_n425), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n517), .A2(new_n518), .A3(new_n519), .A4(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n521), .A2(new_n523), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n429), .A2(new_n526), .A3(new_n519), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n516), .A2(G179), .ZN(new_n528));
  OAI21_X1  g0328(.A(KEYINPUT77), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  AND2_X1   g0329(.A1(new_n525), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n527), .A2(G169), .A3(new_n516), .ZN(new_n531));
  AND3_X1   g0331(.A1(new_n531), .A2(KEYINPUT78), .A3(KEYINPUT21), .ZN(new_n532));
  AOI21_X1  g0332(.A(KEYINPUT21), .B1(new_n531), .B2(KEYINPUT78), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n530), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n516), .B1(new_n527), .B2(G200), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n535), .A2(KEYINPUT79), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT79), .ZN(new_n537));
  AOI211_X1 g0337(.A(new_n537), .B(new_n516), .C1(new_n527), .C2(G200), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n527), .A2(new_n293), .ZN(new_n539));
  NOR3_X1   g0339(.A1(new_n536), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n534), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n280), .A2(new_n227), .A3(G68), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT19), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n543), .B1(new_n254), .B2(new_n205), .ZN(new_n544));
  AOI21_X1  g0344(.A(G20), .B1(new_n305), .B2(KEYINPUT19), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n207), .A2(G87), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n542), .B(new_n544), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n547), .A2(new_n249), .B1(new_n265), .B2(new_n393), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n509), .A2(new_n392), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n263), .A2(G45), .A3(G274), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n263), .A2(G45), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n273), .A2(G250), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(G244), .A2(G1698), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n554), .B1(new_n385), .B2(new_n384), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n472), .B1(new_n555), .B2(new_n280), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n551), .B(new_n553), .C1(new_n556), .C2(new_n273), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(G169), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n278), .A2(G238), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n311), .B1(new_n559), .B2(new_n554), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n272), .B1(new_n560), .B2(new_n472), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n561), .A2(G179), .A3(new_n551), .A4(new_n553), .ZN(new_n562));
  AND3_X1   g0362(.A1(new_n558), .A2(KEYINPUT76), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(KEYINPUT76), .B1(new_n558), .B2(new_n562), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n550), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n557), .A2(G200), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n561), .A2(G190), .A3(new_n551), .A4(new_n553), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n509), .A2(G87), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n566), .A2(new_n567), .A3(new_n548), .A4(new_n568), .ZN(new_n569));
  AND2_X1   g0369(.A1(new_n565), .A2(new_n569), .ZN(new_n570));
  AND4_X1   g0370(.A1(new_n404), .A2(new_n508), .A3(new_n541), .A4(new_n570), .ZN(G372));
  AND2_X1   g0371(.A1(new_n458), .A2(new_n499), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT86), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n558), .A2(new_n562), .B1(new_n548), .B2(new_n549), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n557), .A2(KEYINPUT84), .A3(G200), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n567), .ZN(new_n576));
  AOI21_X1  g0376(.A(KEYINPUT84), .B1(new_n557), .B2(G200), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n548), .A2(new_n568), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(KEYINPUT85), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT85), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n548), .A2(new_n581), .A3(new_n568), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n574), .B1(new_n578), .B2(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n572), .A2(new_n573), .A3(new_n491), .A4(new_n584), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n506), .B(new_n530), .C1(new_n532), .C2(new_n533), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT87), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n574), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n548), .A2(new_n581), .A3(new_n568), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n581), .B1(new_n548), .B2(new_n568), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT84), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n566), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n594), .A2(new_n567), .A3(new_n575), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n589), .B1(new_n592), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(KEYINPUT86), .B1(new_n500), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n531), .A2(KEYINPUT78), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT21), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n531), .A2(KEYINPUT78), .A3(KEYINPUT21), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n602), .A2(KEYINPUT87), .A3(new_n506), .A4(new_n530), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n585), .A2(new_n588), .A3(new_n597), .A4(new_n603), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n493), .A2(new_n497), .A3(new_n498), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n565), .A2(new_n605), .A3(new_n569), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(KEYINPUT26), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT26), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n584), .A2(new_n608), .A3(new_n605), .ZN(new_n609));
  AND3_X1   g0409(.A1(new_n607), .A2(new_n589), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n604), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n404), .A2(new_n611), .ZN(new_n612));
  XOR2_X1   g0412(.A(new_n399), .B(KEYINPUT88), .Z(new_n613));
  INV_X1    g0413(.A(new_n332), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n340), .A2(new_n331), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n615), .A2(new_n616), .B1(new_n374), .B2(new_n372), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n362), .A2(new_n367), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n378), .ZN(new_n619));
  XNOR2_X1  g0419(.A(new_n619), .B(new_n401), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n296), .B1(new_n617), .B2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT89), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n622), .A2(new_n623), .A3(new_n299), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n623), .B1(new_n622), .B2(new_n299), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n612), .B1(new_n624), .B2(new_n625), .ZN(G369));
  INV_X1    g0426(.A(G13), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n627), .A2(G20), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n263), .ZN(new_n629));
  OR2_X1    g0429(.A1(new_n629), .A2(KEYINPUT27), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(KEYINPUT27), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n630), .A2(G213), .A3(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(G343), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n516), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n541), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n534), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n636), .B1(new_n637), .B2(new_n635), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n638), .A2(G330), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n637), .A2(new_n634), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n501), .A2(new_n634), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n507), .B1(new_n491), .B2(new_n642), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n506), .A2(new_n634), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n641), .A2(new_n646), .ZN(new_n647));
  OR2_X1    g0447(.A1(new_n647), .A2(new_n644), .ZN(G399));
  NAND4_X1  g0448(.A1(new_n586), .A2(new_n572), .A3(new_n491), .A4(new_n584), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n570), .A2(new_n608), .A3(new_n605), .ZN(new_n650));
  OAI21_X1  g0450(.A(KEYINPUT26), .B1(new_n596), .B2(new_n499), .ZN(new_n651));
  XOR2_X1   g0451(.A(new_n574), .B(KEYINPUT92), .Z(new_n652));
  NAND4_X1  g0452(.A1(new_n649), .A2(new_n650), .A3(new_n651), .A4(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n634), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT29), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n634), .B1(new_n604), .B2(new_n610), .ZN(new_n658));
  XNOR2_X1  g0458(.A(new_n658), .B(KEYINPUT91), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n657), .B1(new_n659), .B2(new_n656), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n492), .A2(new_n527), .ZN(new_n661));
  INV_X1    g0461(.A(new_n562), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n661), .A2(new_n488), .A3(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT30), .ZN(new_n664));
  OR2_X1    g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n663), .A2(new_n664), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n502), .A2(G179), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n667), .A2(new_n492), .A3(new_n527), .A4(new_n557), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n665), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n634), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n670), .A2(KEYINPUT31), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n541), .A2(new_n508), .A3(new_n570), .A4(new_n654), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n672), .A2(KEYINPUT31), .A3(new_n670), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(G330), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n660), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT93), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n660), .A2(KEYINPUT93), .A3(new_n675), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(new_n263), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n210), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(G41), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NOR3_X1   g0483(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(G1), .A3(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n229), .B2(new_n683), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n686), .B(KEYINPUT90), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(KEYINPUT28), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n680), .A2(new_n688), .ZN(G364));
  AOI21_X1  g0489(.A(new_n226), .B1(G20), .B2(new_n297), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n227), .A2(G190), .ZN(new_n692));
  NOR2_X1   g0492(.A1(G179), .A2(G200), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(G190), .ZN(new_n697));
  XNOR2_X1  g0497(.A(KEYINPUT33), .B(G317), .ZN(new_n698));
  AOI22_X1  g0498(.A1(new_n695), .A2(G329), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(G311), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n692), .A2(G179), .A3(new_n321), .ZN(new_n701));
  OAI211_X1 g0501(.A(new_n699), .B(new_n311), .C1(new_n700), .C2(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n227), .A2(new_n293), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n321), .A2(G179), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(new_n522), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n692), .A2(new_n704), .ZN(new_n707));
  INV_X1    g0507(.A(G283), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n696), .A2(new_n293), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(G326), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NOR4_X1   g0513(.A1(new_n702), .A2(new_n706), .A3(new_n709), .A4(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(G294), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n227), .B1(new_n693), .B2(G190), .ZN(new_n716));
  AND2_X1   g0516(.A1(new_n716), .A2(KEYINPUT95), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n716), .A2(KEYINPUT95), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(G322), .ZN(new_n720));
  INV_X1    g0520(.A(new_n703), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n721), .A2(new_n377), .A3(G200), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  OAI221_X1 g0523(.A(new_n714), .B1(new_n715), .B2(new_n719), .C1(new_n720), .C2(new_n723), .ZN(new_n724));
  XOR2_X1   g0524(.A(new_n724), .B(KEYINPUT96), .Z(new_n725));
  OAI22_X1  g0525(.A1(new_n723), .A2(new_n201), .B1(new_n206), .B2(new_n707), .ZN(new_n726));
  INV_X1    g0526(.A(new_n719), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(G97), .ZN(new_n728));
  INV_X1    g0528(.A(new_n705), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n311), .B1(new_n729), .B2(G87), .ZN(new_n730));
  INV_X1    g0530(.A(G159), .ZN(new_n731));
  OAI21_X1  g0531(.A(KEYINPUT32), .B1(new_n694), .B2(new_n731), .ZN(new_n732));
  OR3_X1    g0532(.A1(new_n694), .A2(KEYINPUT32), .A3(new_n731), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n728), .A2(new_n730), .A3(new_n732), .A4(new_n733), .ZN(new_n734));
  AOI211_X1 g0534(.A(new_n726), .B(new_n734), .C1(G68), .C2(new_n697), .ZN(new_n735));
  OR2_X1    g0535(.A1(new_n701), .A2(KEYINPUT94), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n701), .A2(KEYINPUT94), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  OAI221_X1 g0538(.A(new_n735), .B1(new_n262), .B2(new_n711), .C1(new_n214), .C2(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n691), .B1(new_n725), .B2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(G13), .A2(G33), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(G20), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(new_n690), .ZN(new_n744));
  INV_X1    g0544(.A(G45), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n230), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n681), .A2(new_n280), .ZN(new_n747));
  OAI211_X1 g0547(.A(new_n746), .B(new_n747), .C1(new_n246), .C2(new_n745), .ZN(new_n748));
  INV_X1    g0548(.A(G355), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n280), .A2(new_n210), .ZN(new_n750));
  OAI221_X1 g0550(.A(new_n748), .B1(G116), .B2(new_n210), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n740), .B1(new_n744), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n628), .A2(G45), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n683), .A2(G1), .A3(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n743), .ZN(new_n756));
  OAI211_X1 g0556(.A(new_n752), .B(new_n755), .C1(new_n638), .C2(new_n756), .ZN(new_n757));
  XOR2_X1   g0557(.A(new_n757), .B(KEYINPUT97), .Z(new_n758));
  OR2_X1    g0558(.A1(new_n639), .A2(new_n755), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n638), .A2(G330), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n758), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(G396));
  NAND2_X1  g0563(.A1(new_n396), .A2(new_n634), .ZN(new_n764));
  MUX2_X1   g0564(.A(new_n613), .B(new_n400), .S(new_n764), .Z(new_n765));
  AOI21_X1  g0565(.A(KEYINPUT100), .B1(new_n658), .B2(new_n765), .ZN(new_n766));
  AND4_X1   g0566(.A1(KEYINPUT100), .A2(new_n611), .A3(new_n654), .A4(new_n765), .ZN(new_n767));
  OAI22_X1  g0567(.A1(new_n659), .A2(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n675), .ZN(new_n769));
  XNOR2_X1  g0569(.A(new_n768), .B(new_n769), .ZN(new_n770));
  AND2_X1   g0570(.A1(new_n770), .A2(new_n754), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n707), .A2(new_n344), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n728), .B1(new_n471), .B2(new_n738), .ZN(new_n773));
  AOI211_X1 g0573(.A(new_n772), .B(new_n773), .C1(G294), .C2(new_n722), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n710), .A2(G303), .ZN(new_n775));
  INV_X1    g0575(.A(new_n697), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n776), .A2(new_n708), .B1(new_n694), .B2(new_n700), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n777), .B1(G107), .B2(new_n729), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n774), .A2(new_n311), .A3(new_n775), .A4(new_n778), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n722), .A2(G143), .B1(G150), .B2(new_n697), .ZN(new_n780));
  INV_X1    g0580(.A(G137), .ZN(new_n781));
  OAI221_X1 g0581(.A(new_n780), .B1(new_n781), .B2(new_n711), .C1(new_n738), .C2(new_n731), .ZN(new_n782));
  XOR2_X1   g0582(.A(new_n782), .B(KEYINPUT34), .Z(new_n783));
  INV_X1    g0583(.A(new_n707), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G68), .ZN(new_n785));
  INV_X1    g0585(.A(G132), .ZN(new_n786));
  OAI221_X1 g0586(.A(new_n785), .B1(new_n262), .B2(new_n705), .C1(new_n786), .C2(new_n694), .ZN(new_n787));
  OR3_X1    g0587(.A1(new_n783), .A2(new_n311), .A3(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n719), .A2(new_n201), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n779), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT99), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(new_n690), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n765), .A2(new_n742), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n690), .A2(new_n741), .ZN(new_n795));
  XOR2_X1   g0595(.A(new_n795), .B(KEYINPUT98), .Z(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(new_n214), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NOR4_X1   g0598(.A1(new_n793), .A2(new_n794), .A3(new_n754), .A4(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n771), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(G384));
  INV_X1    g0601(.A(new_n632), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(new_n380), .B2(new_n381), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(KEYINPUT103), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n372), .A2(new_n805), .A3(new_n374), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(new_n620), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n805), .B1(new_n372), .B2(new_n374), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n804), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n619), .A2(new_n373), .ZN(new_n810));
  OAI21_X1  g0610(.A(KEYINPUT37), .B1(new_n804), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n369), .A2(KEYINPUT37), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n812), .A2(new_n382), .A3(new_n803), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(KEYINPUT38), .B1(new_n809), .B2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT38), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n632), .B1(new_n362), .B2(new_n367), .ZN(new_n817));
  OAI21_X1  g0617(.A(KEYINPUT37), .B1(new_n810), .B2(new_n817), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n375), .A2(new_n383), .A3(new_n402), .ZN(new_n819));
  AOI221_X4 g0619(.A(new_n816), .B1(new_n813), .B2(new_n818), .C1(new_n819), .C2(new_n817), .ZN(new_n820));
  OAI21_X1  g0620(.A(KEYINPUT105), .B1(new_n815), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT105), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n819), .A2(new_n817), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n813), .A2(new_n818), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n823), .A2(KEYINPUT38), .A3(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n374), .ZN(new_n826));
  NOR3_X1   g0626(.A1(new_n373), .A2(KEYINPUT72), .A3(KEYINPUT17), .ZN(new_n827));
  OAI21_X1  g0627(.A(KEYINPUT103), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n828), .A2(new_n620), .A3(new_n806), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n829), .A2(new_n804), .B1(new_n813), .B2(new_n811), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n822), .B(new_n825), .C1(new_n830), .C2(KEYINPUT38), .ZN(new_n831));
  AND3_X1   g0631(.A1(new_n821), .A2(new_n831), .A3(KEYINPUT40), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n671), .A2(new_n673), .A3(new_n765), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n331), .A2(new_n634), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n616), .A2(new_n614), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(KEYINPUT102), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT102), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n341), .A2(new_n837), .A3(new_n834), .ZN(new_n838));
  INV_X1    g0638(.A(new_n616), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n836), .A2(new_n838), .B1(new_n839), .B2(new_n634), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n833), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n836), .A2(new_n838), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n839), .A2(new_n634), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n674), .A2(new_n844), .A3(KEYINPUT104), .A4(new_n765), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n823), .A2(new_n824), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(new_n816), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(new_n825), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT104), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(new_n833), .B2(new_n840), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n845), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT40), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n832), .A2(new_n841), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n853), .A2(new_n404), .A3(new_n674), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n851), .A2(new_n852), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n821), .A2(new_n831), .A3(KEYINPUT40), .A4(new_n841), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n855), .A2(G330), .A3(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n769), .A2(new_n404), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n854), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n404), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n660), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n624), .A2(new_n625), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT39), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(new_n815), .B2(new_n820), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n847), .A2(KEYINPUT39), .A3(new_n825), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n616), .A2(new_n634), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n399), .A2(new_n634), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n873), .B1(new_n767), .B2(new_n766), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n874), .A2(new_n848), .A3(new_n844), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n621), .A2(new_n632), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n871), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  XOR2_X1   g0677(.A(new_n865), .B(new_n877), .Z(new_n878));
  OAI21_X1  g0678(.A(new_n861), .B1(new_n878), .B2(KEYINPUT106), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(KEYINPUT106), .ZN(new_n880));
  XOR2_X1   g0680(.A(new_n879), .B(new_n880), .Z(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n263), .B2(new_n628), .ZN(new_n882));
  OAI211_X1 g0682(.A(G116), .B(new_n228), .C1(new_n446), .C2(KEYINPUT35), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n883), .B(KEYINPUT101), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n446), .A2(KEYINPUT35), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n886), .B(KEYINPUT36), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n350), .A2(G77), .ZN(new_n888));
  OAI22_X1  g0688(.A1(new_n229), .A2(new_n888), .B1(G50), .B2(new_n202), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n889), .A2(G1), .A3(new_n627), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n882), .A2(new_n887), .A3(new_n890), .ZN(G367));
  NAND2_X1  g0691(.A1(new_n753), .A2(G1), .ZN(new_n892));
  XOR2_X1   g0692(.A(new_n892), .B(KEYINPUT111), .Z(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT45), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n645), .A2(new_n640), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n896), .A2(new_n644), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT110), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n458), .B(new_n499), .C1(new_n449), .C2(new_n654), .ZN(new_n899));
  OR2_X1    g0699(.A1(new_n899), .A2(KEYINPUT108), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n605), .A2(new_n634), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n899), .A2(KEYINPUT108), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n897), .A2(new_n898), .A3(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n898), .B1(new_n897), .B2(new_n903), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n895), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OR2_X1    g0707(.A1(new_n896), .A2(new_n644), .ZN(new_n908));
  INV_X1    g0708(.A(new_n903), .ZN(new_n909));
  OAI21_X1  g0709(.A(KEYINPUT110), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n910), .A2(KEYINPUT45), .A3(new_n904), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT44), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n912), .B1(new_n908), .B2(new_n909), .ZN(new_n913));
  NOR3_X1   g0713(.A1(new_n897), .A2(KEYINPUT44), .A3(new_n903), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n639), .A2(new_n645), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n907), .A2(new_n911), .A3(new_n915), .A4(new_n916), .ZN(new_n917));
  NOR3_X1   g0717(.A1(new_n639), .A2(new_n645), .A3(new_n640), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n647), .A2(new_n918), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n678), .A2(new_n679), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n682), .B(KEYINPUT41), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n894), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n903), .B(KEYINPUT109), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n507), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n499), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n654), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n896), .A2(new_n903), .ZN(new_n928));
  XOR2_X1   g0728(.A(new_n928), .B(KEYINPUT42), .Z(new_n929));
  NAND2_X1  g0729(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n592), .A2(new_n634), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n584), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n589), .B2(new_n931), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(KEYINPUT43), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n933), .B(KEYINPUT107), .Z(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n936), .A2(KEYINPUT43), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n930), .A2(new_n934), .A3(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n927), .A2(new_n929), .A3(new_n937), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n924), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n941), .B1(new_n916), .B2(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n942), .A2(new_n916), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n939), .A2(new_n944), .A3(new_n940), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n923), .A2(new_n943), .A3(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT46), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n705), .B2(new_n471), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n948), .A2(KEYINPUT112), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n722), .A2(G303), .B1(new_n710), .B2(G311), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n729), .A2(KEYINPUT46), .A3(G116), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n948), .A2(KEYINPUT112), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n949), .A2(new_n950), .A3(new_n951), .A4(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n707), .A2(new_n205), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(new_n727), .B2(G107), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n280), .B1(new_n695), .B2(G317), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n955), .B(new_n956), .C1(new_n715), .C2(new_n776), .ZN(new_n957));
  INV_X1    g0757(.A(new_n738), .ZN(new_n958));
  AOI211_X1 g0758(.A(new_n953), .B(new_n957), .C1(G283), .C2(new_n958), .ZN(new_n959));
  AOI22_X1  g0759(.A1(new_n958), .A2(G50), .B1(G77), .B2(new_n784), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n727), .A2(G68), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n960), .B(new_n961), .C1(new_n781), .C2(new_n694), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n710), .A2(G143), .ZN(new_n963));
  OAI221_X1 g0763(.A(new_n963), .B1(new_n201), .B2(new_n705), .C1(new_n723), .C2(new_n255), .ZN(new_n964));
  NOR3_X1   g0764(.A1(new_n962), .A2(new_n311), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n697), .A2(G159), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n959), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n967), .B(KEYINPUT47), .Z(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n690), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n933), .A2(new_n756), .ZN(new_n970));
  INV_X1    g0770(.A(new_n747), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n744), .B1(new_n210), .B2(new_n393), .C1(new_n238), .C2(new_n971), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n969), .A2(new_n970), .A3(new_n755), .A4(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n946), .A2(new_n973), .ZN(G387));
  NAND2_X1  g0774(.A1(new_n678), .A2(new_n679), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n919), .ZN(new_n976));
  INV_X1    g0776(.A(new_n919), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n678), .A2(new_n679), .A3(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n976), .A2(new_n682), .A3(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n747), .B1(new_n235), .B2(new_n745), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n684), .B2(new_n750), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n251), .A2(G50), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT50), .ZN(new_n983));
  AOI21_X1  g0783(.A(G45), .B1(G68), .B2(G77), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n983), .A2(new_n684), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n981), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(G107), .B2(new_n210), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n744), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n645), .B2(new_n756), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n722), .A2(G317), .B1(G311), .B2(new_n697), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n990), .B1(new_n720), .B2(new_n711), .C1(new_n738), .C2(new_n522), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT48), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n992), .B1(new_n708), .B2(new_n719), .C1(new_n715), .C2(new_n705), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT113), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT49), .ZN(new_n995));
  OR2_X1    g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n994), .A2(new_n995), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n784), .A2(G116), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n996), .A2(new_n997), .A3(new_n311), .A4(new_n998), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n694), .A2(new_n712), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n280), .B1(new_n776), .B2(new_n251), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n719), .A2(new_n393), .ZN(new_n1002));
  AOI211_X1 g0802(.A(new_n1001), .B(new_n1002), .C1(G150), .C2(new_n695), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n1003), .B1(new_n202), .B2(new_n701), .C1(new_n214), .C2(new_n705), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n954), .B1(new_n722), .B2(G50), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n731), .B2(new_n711), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n999), .A2(new_n1000), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n989), .B1(new_n1007), .B2(new_n690), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n1008), .A2(new_n755), .B1(new_n919), .B2(new_n893), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n979), .A2(new_n1009), .ZN(G393));
  AOI21_X1  g0810(.A(new_n977), .B1(new_n678), .B2(new_n679), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n917), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n907), .A2(new_n915), .A3(new_n911), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(new_n916), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1012), .B(new_n682), .C1(new_n1014), .C2(new_n1011), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n942), .A2(new_n743), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n744), .B1(new_n243), .B2(new_n971), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(G97), .B2(new_n681), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n722), .A2(G311), .B1(new_n710), .B2(G317), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT52), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n727), .A2(G116), .B1(G303), .B2(new_n697), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1021), .A2(KEYINPUT115), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n1020), .B(new_n1022), .C1(G107), .C2(new_n784), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n311), .B1(new_n705), .B2(new_n708), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(new_n1021), .B2(KEYINPUT115), .ZN(new_n1025));
  AND2_X1   g0825(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1026), .B1(new_n715), .B2(new_n701), .C1(new_n720), .C2(new_n694), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n727), .A2(G77), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1028), .B1(new_n262), .B2(new_n776), .C1(new_n251), .C2(new_n738), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT114), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n772), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n311), .B1(new_n695), .B2(G143), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n729), .A2(G68), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .A4(new_n1033), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n722), .A2(G159), .B1(new_n710), .B2(G150), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT51), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1027), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT116), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n754), .B(new_n1018), .C1(new_n1038), .C2(new_n690), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n1014), .A2(new_n893), .B1(new_n1016), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1015), .A2(new_n1040), .ZN(G390));
  NAND3_X1  g0841(.A1(new_n765), .A2(new_n654), .A3(new_n653), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n873), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n870), .B1(new_n1043), .B2(new_n844), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1044), .A2(new_n821), .A3(new_n831), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n870), .B1(new_n874), .B2(new_n844), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1045), .B1(new_n1046), .B2(new_n869), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(KEYINPUT117), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n841), .A2(G330), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT117), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1051), .B(new_n1045), .C1(new_n1046), .C2(new_n869), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1048), .A2(new_n1050), .A3(new_n1052), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1047), .A2(KEYINPUT117), .A3(new_n1049), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NOR3_X1   g0855(.A1(new_n863), .A2(new_n864), .A3(new_n860), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n674), .A2(G330), .A3(new_n765), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(new_n840), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(new_n1049), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n874), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n1043), .B2(new_n1059), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1056), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1055), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1053), .A2(new_n1054), .A3(new_n1062), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1064), .A2(new_n682), .A3(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n894), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1067));
  OR2_X1    g0867(.A1(new_n869), .A2(new_n742), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n280), .B1(new_n707), .B2(new_n262), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n729), .A2(G150), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT53), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n1069), .B(new_n1071), .C1(G159), .C2(new_n727), .ZN(new_n1072));
  XOR2_X1   g0872(.A(KEYINPUT54), .B(G143), .Z(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n738), .A2(new_n1074), .B1(new_n781), .B2(new_n776), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT118), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n710), .A2(G128), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n722), .A2(G132), .B1(G125), .B2(new_n695), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n1072), .A2(new_n1076), .A3(new_n1077), .A4(new_n1078), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n958), .A2(G97), .B1(G107), .B2(new_n697), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n1080), .A2(KEYINPUT119), .B1(G68), .B2(new_n784), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n1081), .B1(new_n471), .B2(new_n723), .C1(new_n708), .C2(new_n711), .ZN(new_n1082));
  OR2_X1    g0882(.A1(new_n1082), .A2(new_n280), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1080), .A2(KEYINPUT119), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(G77), .B2(new_n727), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n1085), .B1(new_n344), .B2(new_n705), .C1(new_n715), .C2(new_n694), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1079), .B1(new_n1083), .B2(new_n1086), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT120), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n690), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1068), .A2(new_n755), .A3(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(new_n251), .B2(new_n796), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1067), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1066), .A2(new_n1092), .ZN(G378));
  NAND3_X1  g0893(.A1(new_n300), .A2(new_n269), .A3(new_n802), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n269), .A2(new_n802), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n296), .A2(new_n299), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1094), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1101));
  AND2_X1   g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n741), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n707), .A2(new_n201), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n727), .A2(G68), .B1(G107), .B2(new_n722), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n1105), .B1(new_n205), .B2(new_n776), .C1(new_n393), .C2(new_n701), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n1104), .B(new_n1106), .C1(G283), .C2(new_n695), .ZN(new_n1107));
  AOI211_X1 g0907(.A(G41), .B(new_n280), .C1(new_n729), .C2(G77), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1107), .B(new_n1108), .C1(new_n471), .C2(new_n711), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1109), .B(KEYINPUT58), .ZN(new_n1110));
  AOI21_X1  g0910(.A(G50), .B1(new_n311), .B2(new_n415), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(G33), .A2(G41), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT121), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n1074), .A2(new_n705), .B1(new_n786), .B2(new_n776), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1115), .B1(G125), .B2(new_n710), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n701), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n722), .A2(G128), .B1(G137), .B2(new_n1117), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1116), .B(new_n1118), .C1(new_n255), .C2(new_n719), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT59), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1113), .B1(G124), .B2(new_n695), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1121), .B1(new_n731), .B2(new_n707), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1110), .B(new_n1114), .C1(new_n1120), .C2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n690), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n754), .B1(new_n262), .B2(new_n795), .ZN(new_n1125));
  XOR2_X1   g0925(.A(new_n1125), .B(KEYINPUT122), .Z(new_n1126));
  AND3_X1   g0926(.A1(new_n1103), .A2(new_n1124), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(new_n853), .B2(G330), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n857), .A2(new_n1102), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n877), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n853), .A2(G330), .A3(new_n1128), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n877), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n857), .A2(new_n1102), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1131), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1127), .B1(new_n1136), .B2(new_n893), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1064), .A2(new_n1056), .ZN(new_n1138));
  AOI21_X1  g0938(.A(KEYINPUT57), .B1(new_n1138), .B2(new_n1136), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1062), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1056), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1136), .A2(KEYINPUT57), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n682), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1137), .B1(new_n1139), .B2(new_n1144), .ZN(G375));
  INV_X1    g0945(.A(new_n1061), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1141), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1147), .A2(new_n921), .A3(new_n1062), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n840), .A2(new_n741), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1104), .B1(G150), .B2(new_n1117), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n311), .B1(new_n695), .B2(G128), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1150), .B(new_n1151), .C1(new_n731), .C2(new_n705), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1152), .B1(G50), .B2(new_n727), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT123), .ZN(new_n1154));
  OAI221_X1 g0954(.A(new_n1154), .B1(new_n786), .B2(new_n711), .C1(new_n776), .C2(new_n1074), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(G137), .B2(new_n722), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1002), .B1(G283), .B2(new_n722), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n1157), .B1(new_n206), .B2(new_n738), .C1(new_n715), .C2(new_n711), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n694), .A2(new_n522), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n311), .B1(new_n707), .B2(new_n214), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n776), .A2(new_n471), .B1(new_n705), .B2(new_n205), .ZN(new_n1161));
  NOR4_X1   g0961(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .A4(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n690), .B1(new_n1156), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n796), .A2(new_n202), .ZN(new_n1164));
  AND4_X1   g0964(.A1(new_n755), .A2(new_n1149), .A3(new_n1163), .A4(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(new_n1061), .B2(new_n893), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1148), .A2(new_n1166), .ZN(G381));
  INV_X1    g0967(.A(new_n1137), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT57), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(new_n1131), .B2(new_n1135), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n683), .B1(new_n1138), .B2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1136), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(new_n1169), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1168), .B1(new_n1171), .B2(new_n1173), .ZN(new_n1174));
  AND3_X1   g0974(.A1(new_n1053), .A2(new_n1054), .A3(new_n1062), .ZN(new_n1175));
  NOR3_X1   g0975(.A1(new_n1175), .A2(new_n1140), .A3(new_n683), .ZN(new_n1176));
  OR2_X1    g0976(.A1(new_n1067), .A2(new_n1091), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1174), .A2(new_n1178), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n946), .A2(new_n1015), .A3(new_n973), .A4(new_n1040), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n979), .A2(new_n762), .A3(new_n1009), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1181), .A2(G384), .ZN(new_n1182));
  XOR2_X1   g0982(.A(new_n1182), .B(KEYINPUT124), .Z(new_n1183));
  OR4_X1    g0983(.A1(G381), .A2(new_n1179), .A3(new_n1180), .A4(new_n1183), .ZN(G407));
  OAI211_X1 g0984(.A(G407), .B(G213), .C1(G343), .C2(new_n1179), .ZN(G409));
  OAI211_X1 g0985(.A(new_n1136), .B(new_n921), .C1(new_n1140), .C2(new_n1141), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1186), .A2(new_n1137), .ZN(new_n1187));
  INV_X1    g0987(.A(G213), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n1187), .A2(G378), .B1(new_n1188), .B2(G343), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(G378), .B2(G375), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1188), .A2(G343), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT60), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n683), .B1(new_n1147), .B2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1141), .A2(KEYINPUT60), .A3(new_n1146), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1193), .A2(new_n1062), .A3(new_n1194), .ZN(new_n1195));
  AND3_X1   g0995(.A1(new_n1195), .A2(G384), .A3(new_n1166), .ZN(new_n1196));
  AOI21_X1  g0996(.A(G384), .B1(new_n1195), .B2(new_n1166), .ZN(new_n1197));
  OAI211_X1 g0997(.A(G2897), .B(new_n1191), .C1(new_n1196), .C2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1197), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1195), .A2(G384), .A3(new_n1166), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1191), .A2(G2897), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1198), .A2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(KEYINPUT63), .B1(new_n1190), .B2(new_n1203), .ZN(new_n1204));
  AND2_X1   g1004(.A1(new_n1186), .A2(new_n1137), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1191), .B1(new_n1205), .B2(new_n1178), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1206), .B(new_n1207), .C1(new_n1178), .C2(new_n1174), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1204), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(G393), .A2(G396), .ZN(new_n1210));
  AND2_X1   g1010(.A1(new_n1210), .A2(new_n1181), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1180), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n946), .A2(new_n973), .B1(new_n1015), .B2(new_n1040), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1211), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(G387), .A2(G390), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1210), .A2(new_n1181), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1215), .A2(new_n1216), .A3(new_n1180), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1214), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1208), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1218), .B1(new_n1219), .B2(KEYINPUT63), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT61), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1209), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  AND3_X1   g1022(.A1(new_n1208), .A2(KEYINPUT125), .A3(KEYINPUT62), .ZN(new_n1223));
  AOI21_X1  g1023(.A(KEYINPUT62), .B1(new_n1208), .B2(KEYINPUT125), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1221), .B1(new_n1190), .B2(new_n1203), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(new_n1223), .A2(new_n1224), .A3(new_n1225), .ZN(new_n1226));
  AND3_X1   g1026(.A1(new_n1214), .A2(KEYINPUT126), .A3(new_n1217), .ZN(new_n1227));
  AOI21_X1  g1027(.A(KEYINPUT126), .B1(new_n1214), .B2(new_n1217), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1222), .B1(new_n1226), .B2(new_n1230), .ZN(G405));
  NOR2_X1   g1031(.A1(G375), .A2(G378), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1171), .A2(new_n1173), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1178), .B1(new_n1233), .B2(new_n1137), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n1232), .A2(new_n1234), .B1(new_n1197), .B2(new_n1196), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(G375), .A2(G378), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1236), .A2(new_n1179), .A3(new_n1207), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1235), .A2(new_n1229), .A3(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT127), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1235), .A2(new_n1237), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n1230), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1235), .A2(new_n1229), .A3(KEYINPUT127), .A4(new_n1237), .ZN(new_n1243));
  AND3_X1   g1043(.A1(new_n1240), .A2(new_n1242), .A3(new_n1243), .ZN(G402));
endmodule


