//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 0 1 0 0 0 1 1 0 1 0 0 1 1 0 1 0 1 0 1 1 1 0 0 1 1 1 1 0 0 1 0 1 0 1 1 0 0 0 1 1 1 1 0 1 0 1 1 0 0 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:21 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1220, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1272, new_n1273, new_n1274;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT64), .Z(new_n209));
  INV_X1    g0009(.A(G58), .ZN(new_n210));
  INV_X1    g0010(.A(G232), .ZN(new_n211));
  INV_X1    g0011(.A(G244), .ZN(new_n212));
  OAI22_X1  g0012(.A1(new_n210), .A2(new_n211), .B1(new_n202), .B2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(G68), .ZN(new_n214));
  INV_X1    g0014(.A(G238), .ZN(new_n215));
  INV_X1    g0015(.A(G87), .ZN(new_n216));
  INV_X1    g0016(.A(G250), .ZN(new_n217));
  OAI22_X1  g0017(.A1(new_n214), .A2(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(G97), .ZN(new_n219));
  INV_X1    g0019(.A(G257), .ZN(new_n220));
  INV_X1    g0020(.A(G107), .ZN(new_n221));
  INV_X1    g0021(.A(G264), .ZN(new_n222));
  OAI22_X1  g0022(.A1(new_n219), .A2(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NOR3_X1   g0023(.A1(new_n213), .A2(new_n218), .A3(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n207), .B1(new_n209), .B2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(KEYINPUT1), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT65), .Z(new_n228));
  INV_X1    g0028(.A(G13), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n207), .A2(new_n229), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n231), .B(G250), .C1(G257), .C2(G264), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT0), .ZN(new_n233));
  OAI21_X1  g0033(.A(G50), .B1(G58), .B2(G68), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g0035(.A1(G1), .A2(G13), .ZN(new_n236));
  NOR2_X1   g0036(.A1(new_n236), .A2(new_n206), .ZN(new_n237));
  NAND2_X1  g0037(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  OAI211_X1 g0038(.A(new_n233), .B(new_n238), .C1(new_n226), .C2(new_n225), .ZN(new_n239));
  NOR2_X1   g0039(.A1(new_n228), .A2(new_n239), .ZN(G361));
  XNOR2_X1  g0040(.A(G238), .B(G244), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G232), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT2), .B(G226), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G250), .B(G257), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G264), .B(G270), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G358));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XOR2_X1   g0049(.A(G107), .B(G116), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G50), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G68), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n214), .A2(G50), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(G58), .B(G77), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XOR2_X1   g0057(.A(new_n251), .B(new_n257), .Z(G351));
  INV_X1    g0058(.A(G150), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G20), .A2(G33), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  OAI22_X1  g0061(.A1(new_n259), .A2(new_n261), .B1(new_n201), .B2(new_n206), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT8), .B(G58), .ZN(new_n263));
  XNOR2_X1  g0063(.A(new_n263), .B(KEYINPUT67), .ZN(new_n264));
  INV_X1    g0064(.A(G33), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(G20), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n262), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(new_n236), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  NOR3_X1   g0071(.A1(new_n229), .A2(new_n206), .A3(G1), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(new_n252), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n205), .A2(G20), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n270), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n273), .B1(new_n275), .B2(new_n252), .ZN(new_n276));
  OR2_X1    g0076(.A1(new_n271), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT9), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n271), .A2(new_n276), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(KEYINPUT9), .ZN(new_n281));
  AND2_X1   g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT10), .ZN(new_n283));
  INV_X1    g0083(.A(G41), .ZN(new_n284));
  OAI211_X1 g0084(.A(G1), .B(G13), .C1(new_n265), .C2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G274), .ZN(new_n286));
  INV_X1    g0086(.A(G45), .ZN(new_n287));
  AOI21_X1  g0087(.A(G1), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n285), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n290), .B1(G226), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n265), .A2(KEYINPUT3), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT3), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G33), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G1698), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G222), .ZN(new_n300));
  OAI22_X1  g0100(.A1(new_n299), .A2(new_n300), .B1(new_n202), .B2(new_n297), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n294), .A2(new_n296), .A3(G1698), .ZN(new_n302));
  XNOR2_X1  g0102(.A(new_n302), .B(KEYINPUT66), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n301), .B1(G223), .B2(new_n303), .ZN(new_n304));
  OAI211_X1 g0104(.A(G190), .B(new_n293), .C1(new_n304), .C2(new_n285), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n293), .B1(new_n304), .B2(new_n285), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G200), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n282), .A2(new_n283), .A3(new_n305), .A4(new_n307), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n279), .A2(new_n305), .A3(new_n307), .A4(new_n281), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(KEYINPUT10), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n266), .A2(G77), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n214), .A2(G20), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n313), .B(new_n314), .C1(new_n252), .C2(new_n261), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(new_n269), .ZN(new_n316));
  XNOR2_X1  g0116(.A(new_n316), .B(KEYINPUT11), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n229), .A2(G1), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G20), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT68), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n272), .A2(KEYINPUT68), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n324), .A2(new_n269), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n325), .A2(G68), .A3(new_n274), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT12), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n327), .B1(new_n324), .B2(new_n214), .ZN(new_n328));
  NOR4_X1   g0128(.A1(new_n314), .A2(KEYINPUT12), .A3(G1), .A4(new_n229), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n317), .B(new_n326), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n294), .A2(new_n296), .A3(G232), .A4(G1698), .ZN(new_n331));
  OR2_X1    g0131(.A1(new_n331), .A2(KEYINPUT69), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(KEYINPUT69), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n294), .A2(new_n296), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n335), .A2(G1698), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n336), .A2(G226), .B1(G33), .B2(G97), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n285), .B1(new_n334), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n290), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n339), .B1(new_n215), .B2(new_n291), .ZN(new_n340));
  OAI21_X1  g0140(.A(KEYINPUT13), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n290), .B1(G238), .B2(new_n292), .ZN(new_n342));
  XNOR2_X1  g0142(.A(KEYINPUT70), .B(KEYINPUT13), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n297), .A2(G226), .A3(new_n298), .ZN(new_n344));
  NAND2_X1  g0144(.A1(G33), .A2(G97), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n346), .B1(new_n332), .B2(new_n333), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n342), .B(new_n343), .C1(new_n347), .C2(new_n285), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n341), .A2(new_n348), .A3(G179), .ZN(new_n349));
  INV_X1    g0149(.A(G169), .ZN(new_n350));
  INV_X1    g0150(.A(new_n343), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n351), .B1(new_n338), .B2(new_n340), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n350), .B1(new_n352), .B2(new_n348), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT14), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n349), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  AOI211_X1 g0155(.A(KEYINPUT14), .B(new_n350), .C1(new_n352), .C2(new_n348), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n330), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n352), .A2(new_n348), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n330), .B1(new_n358), .B2(G200), .ZN(new_n359));
  INV_X1    g0159(.A(G190), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n338), .A2(new_n340), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n360), .B1(new_n361), .B2(new_n343), .ZN(new_n362));
  AND3_X1   g0162(.A1(new_n362), .A2(KEYINPUT71), .A3(new_n341), .ZN(new_n363));
  AOI21_X1  g0163(.A(KEYINPUT71), .B1(new_n362), .B2(new_n341), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n359), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n357), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n280), .B1(new_n306), .B2(new_n350), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(G179), .B2(new_n306), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n290), .B1(G244), .B2(new_n292), .ZN(new_n369));
  OAI22_X1  g0169(.A1(new_n299), .A2(new_n211), .B1(new_n221), .B2(new_n297), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n370), .B1(G238), .B2(new_n303), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n369), .B1(new_n371), .B2(new_n285), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(G200), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n325), .A2(G77), .A3(new_n274), .ZN(new_n374));
  XOR2_X1   g0174(.A(KEYINPUT15), .B(G87), .Z(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(new_n266), .ZN(new_n376));
  OAI221_X1 g0176(.A(new_n376), .B1(new_n206), .B2(new_n202), .C1(new_n261), .C2(new_n263), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n377), .A2(new_n269), .B1(new_n202), .B2(new_n324), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n374), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n373), .B(new_n380), .C1(new_n360), .C2(new_n372), .ZN(new_n381));
  INV_X1    g0181(.A(new_n370), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n303), .A2(G238), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n285), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n369), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n350), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(G179), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n387), .B(new_n369), .C1(new_n371), .C2(new_n285), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n386), .A2(new_n388), .A3(new_n379), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n368), .A2(new_n381), .A3(new_n389), .ZN(new_n390));
  NOR3_X1   g0190(.A1(new_n312), .A2(new_n366), .A3(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(KEYINPUT72), .B1(new_n295), .B2(G33), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT72), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n393), .A2(new_n265), .A3(KEYINPUT3), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NOR2_X1   g0195(.A1(G223), .A2(G1698), .ZN(new_n396));
  INV_X1    g0196(.A(G226), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n396), .B1(new_n397), .B2(G1698), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n395), .A2(new_n398), .A3(new_n296), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n265), .A2(new_n216), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT75), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n399), .A2(KEYINPUT75), .A3(new_n401), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n285), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(KEYINPUT76), .B1(new_n291), .B2(new_n211), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT76), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n289), .A2(new_n408), .A3(G232), .A4(new_n285), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n339), .ZN(new_n411));
  OAI21_X1  g0211(.A(G169), .B1(new_n406), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n236), .B1(G33), .B2(G41), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n265), .A2(KEYINPUT3), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n414), .B1(new_n392), .B2(new_n394), .ZN(new_n415));
  AOI211_X1 g0215(.A(new_n403), .B(new_n400), .C1(new_n415), .C2(new_n398), .ZN(new_n416));
  AOI21_X1  g0216(.A(KEYINPUT75), .B1(new_n399), .B2(new_n401), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n413), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n290), .B1(new_n407), .B2(new_n409), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n418), .A2(G179), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n412), .A2(new_n420), .ZN(new_n421));
  OR2_X1    g0221(.A1(new_n264), .A2(new_n272), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n264), .A2(new_n275), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n395), .A2(new_n296), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT7), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n425), .A2(new_n426), .A3(new_n206), .ZN(new_n427));
  OAI21_X1  g0227(.A(KEYINPUT7), .B1(new_n415), .B2(G20), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n427), .A2(G68), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(G58), .A2(G68), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(KEYINPUT73), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT73), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n432), .A2(G58), .A3(G68), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n431), .B(new_n433), .C1(G58), .C2(G68), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n434), .A2(G20), .B1(G159), .B2(new_n260), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n429), .A2(KEYINPUT16), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n269), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n294), .A2(KEYINPUT74), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT74), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n439), .A2(new_n265), .A3(KEYINPUT3), .ZN(new_n440));
  AND3_X1   g0240(.A1(new_n438), .A2(new_n440), .A3(new_n296), .ZN(new_n441));
  OAI21_X1  g0241(.A(KEYINPUT7), .B1(new_n441), .B2(G20), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n335), .A2(new_n426), .A3(new_n206), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n442), .A2(G68), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(KEYINPUT16), .B1(new_n444), .B2(new_n435), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n424), .B1(new_n437), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(KEYINPUT18), .B1(new_n421), .B2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n421), .A2(new_n446), .A3(KEYINPUT18), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n448), .A2(KEYINPUT77), .A3(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT77), .ZN(new_n451));
  INV_X1    g0251(.A(new_n449), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n451), .B1(new_n452), .B2(new_n447), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n446), .ZN(new_n455));
  AND3_X1   g0255(.A1(new_n418), .A2(new_n360), .A3(new_n419), .ZN(new_n456));
  AOI21_X1  g0256(.A(G200), .B1(new_n418), .B2(new_n419), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT78), .ZN(new_n458));
  NOR3_X1   g0258(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(G200), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n460), .B1(new_n406), .B2(new_n411), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n418), .A2(new_n360), .A3(new_n419), .ZN(new_n462));
  AOI21_X1  g0262(.A(KEYINPUT78), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n455), .B1(new_n459), .B2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT79), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n458), .B1(new_n456), .B2(new_n457), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n461), .A2(KEYINPUT78), .A3(new_n462), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n446), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(KEYINPUT79), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n466), .A2(new_n470), .A3(KEYINPUT17), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT17), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n472), .B(new_n455), .C1(new_n459), .C2(new_n463), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT80), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n469), .A2(KEYINPUT80), .A3(new_n472), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n454), .B1(new_n471), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n391), .A2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  AND2_X1   g0280(.A1(KEYINPUT4), .A2(G244), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n297), .A2(KEYINPUT83), .A3(new_n298), .A4(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n297), .A2(G250), .A3(G1698), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n294), .A2(new_n296), .A3(new_n481), .A4(new_n298), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT83), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(G33), .A2(G283), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n482), .A2(new_n483), .A3(new_n486), .A4(new_n487), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n212), .A2(G1698), .ZN(new_n489));
  AOI21_X1  g0289(.A(KEYINPUT4), .B1(new_n415), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n413), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(G274), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n413), .A2(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n287), .A2(G1), .ZN(new_n494));
  XNOR2_X1  g0294(.A(KEYINPUT5), .B(G41), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n413), .B1(new_n494), .B2(new_n495), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(G257), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n491), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  OR2_X1    g0299(.A1(new_n499), .A2(G179), .ZN(new_n500));
  XNOR2_X1  g0300(.A(G97), .B(G107), .ZN(new_n501));
  NOR2_X1   g0301(.A1(KEYINPUT81), .A2(KEYINPUT6), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n502), .B1(KEYINPUT6), .B2(new_n219), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n504), .B1(new_n501), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(KEYINPUT82), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT82), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n504), .B(new_n508), .C1(new_n501), .C2(new_n505), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n507), .A2(G20), .A3(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n442), .A2(G107), .A3(new_n443), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n260), .A2(G77), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n269), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n272), .A2(new_n219), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n205), .A2(G33), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n270), .A2(new_n319), .A3(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n515), .B1(new_n517), .B2(new_n219), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n514), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n499), .A2(new_n350), .ZN(new_n521));
  AND3_X1   g0321(.A1(new_n500), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n518), .B1(new_n513), .B2(new_n269), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n499), .A2(G200), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n491), .A2(G190), .A3(new_n496), .A4(new_n498), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT84), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n523), .A2(new_n524), .A3(KEYINPUT84), .A4(new_n525), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n522), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT89), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT23), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n532), .A2(new_n221), .A3(G20), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(KEYINPUT88), .ZN(new_n534));
  NAND2_X1  g0334(.A1(KEYINPUT23), .A2(G107), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n537));
  OAI22_X1  g0337(.A1(new_n533), .A2(KEYINPUT88), .B1(new_n537), .B2(G20), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n415), .A2(KEYINPUT22), .A3(new_n206), .A4(G87), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT22), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n206), .A2(G87), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n541), .B1(new_n335), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n539), .A2(new_n540), .A3(new_n543), .ZN(new_n544));
  OR2_X1    g0344(.A1(new_n544), .A2(KEYINPUT24), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(KEYINPUT24), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n270), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n272), .A2(new_n221), .ZN(new_n548));
  XOR2_X1   g0348(.A(new_n548), .B(KEYINPUT25), .Z(new_n549));
  OAI21_X1  g0349(.A(new_n549), .B1(new_n221), .B2(new_n517), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n495), .A2(new_n494), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n285), .ZN(new_n553));
  NOR2_X1   g0353(.A1(G250), .A2(G1698), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n554), .B1(new_n220), .B2(G1698), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n415), .A2(new_n555), .B1(G33), .B2(G294), .ZN(new_n556));
  OAI221_X1 g0356(.A(new_n496), .B1(new_n553), .B2(new_n222), .C1(new_n556), .C2(new_n285), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n387), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n557), .A2(new_n350), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n551), .A2(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n496), .B1(new_n222), .B2(new_n553), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n556), .A2(new_n285), .ZN(new_n564));
  OAI21_X1  g0364(.A(G200), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(new_n557), .B2(new_n360), .ZN(new_n566));
  NOR3_X1   g0366(.A1(new_n547), .A2(new_n566), .A3(new_n550), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n531), .B1(new_n562), .B2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(new_n566), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n551), .A2(new_n569), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n560), .B(new_n559), .C1(new_n547), .C2(new_n550), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n570), .A2(KEYINPUT89), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n487), .B(new_n206), .C1(G33), .C2(new_n219), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n574), .B(new_n269), .C1(new_n206), .C2(G116), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT20), .ZN(new_n576));
  XNOR2_X1  g0376(.A(new_n575), .B(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(G116), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n324), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n323), .A2(G116), .A3(new_n270), .A4(new_n516), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n577), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(G270), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n496), .B1(new_n582), .B2(new_n553), .ZN(new_n583));
  NOR2_X1   g0383(.A1(G257), .A2(G1698), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n584), .B1(new_n222), .B2(G1698), .ZN(new_n585));
  XOR2_X1   g0385(.A(KEYINPUT86), .B(G303), .Z(new_n586));
  AOI22_X1  g0386(.A1(new_n415), .A2(new_n585), .B1(new_n586), .B2(new_n335), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n587), .A2(new_n285), .ZN(new_n588));
  OR2_X1    g0388(.A1(new_n583), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n581), .B1(new_n589), .B2(G200), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT87), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n583), .A2(new_n588), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n590), .A2(new_n591), .B1(G190), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n592), .A2(new_n460), .ZN(new_n594));
  OAI21_X1  g0394(.A(KEYINPUT87), .B1(new_n594), .B2(new_n581), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n589), .A2(G169), .A3(new_n581), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT21), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n589), .A2(KEYINPUT21), .A3(new_n581), .A4(G169), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n581), .A2(new_n592), .A3(G179), .ZN(new_n601));
  AND3_X1   g0401(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT85), .ZN(new_n603));
  AOI21_X1  g0403(.A(KEYINPUT19), .B1(new_n266), .B2(G97), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT19), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n206), .B1(new_n345), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n216), .A2(new_n219), .A3(new_n221), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n604), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n415), .A2(new_n206), .A3(G68), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n269), .ZN(new_n611));
  INV_X1    g0411(.A(new_n375), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n324), .A2(new_n612), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n611), .B(new_n613), .C1(new_n612), .C2(new_n517), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n494), .A2(new_n217), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n493), .A2(new_n494), .B1(new_n285), .B2(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(G238), .A2(G1698), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n617), .B1(new_n212), .B2(G1698), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n415), .A2(new_n618), .B1(G33), .B2(G116), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n616), .B1(new_n619), .B2(new_n285), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(G179), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n620), .A2(G169), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n603), .A2(new_n614), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  OR2_X1    g0424(.A1(new_n614), .A2(new_n603), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n621), .A2(G190), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n620), .A2(G200), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n611), .A2(new_n613), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n517), .A2(new_n216), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n624), .A2(new_n625), .B1(new_n628), .B2(new_n632), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n596), .A2(new_n602), .A3(new_n633), .ZN(new_n634));
  AND4_X1   g0434(.A1(new_n480), .A2(new_n530), .A3(new_n573), .A4(new_n634), .ZN(G372));
  XNOR2_X1  g0435(.A(new_n311), .B(KEYINPUT90), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n467), .A2(new_n468), .ZN(new_n637));
  AOI21_X1  g0437(.A(KEYINPUT79), .B1(new_n637), .B2(new_n455), .ZN(new_n638));
  AOI211_X1 g0438(.A(new_n465), .B(new_n446), .C1(new_n467), .C2(new_n468), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  AOI22_X1  g0440(.A1(new_n640), .A2(KEYINPUT17), .B1(new_n475), .B2(new_n476), .ZN(new_n641));
  INV_X1    g0441(.A(new_n389), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n365), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n641), .B1(new_n357), .B2(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n452), .A2(new_n447), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n636), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n528), .A2(new_n529), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n622), .A2(new_n623), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(new_n614), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n626), .A2(new_n629), .A3(new_n631), .A4(new_n627), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n651), .A2(new_n567), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n571), .A2(new_n599), .A3(new_n600), .A4(new_n601), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n500), .A2(new_n520), .A3(new_n521), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n647), .A2(new_n652), .A3(new_n653), .A4(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n522), .A2(new_n633), .A3(KEYINPUT26), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT26), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n657), .B1(new_n654), .B2(new_n651), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n655), .A2(new_n659), .A3(new_n649), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n646), .B(new_n368), .C1(new_n479), .C2(new_n661), .ZN(G369));
  INV_X1    g0462(.A(new_n573), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n318), .A2(new_n206), .ZN(new_n664));
  OR2_X1    g0464(.A1(new_n664), .A2(KEYINPUT27), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(KEYINPUT27), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n665), .A2(G213), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n667), .B(KEYINPUT91), .ZN(new_n668));
  INV_X1    g0468(.A(G343), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n602), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n663), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n670), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n672), .B1(new_n562), .B2(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n670), .B1(new_n547), .B2(new_n550), .ZN(new_n675));
  AOI22_X1  g0475(.A1(new_n573), .A2(new_n675), .B1(new_n562), .B2(new_n670), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n670), .A2(new_n581), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n596), .A2(new_n602), .A3(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n678), .B1(new_n602), .B2(new_n677), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(G330), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n676), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n674), .A2(new_n681), .ZN(new_n682));
  XOR2_X1   g0482(.A(new_n682), .B(KEYINPUT92), .Z(G399));
  NOR2_X1   g0483(.A1(new_n230), .A2(G41), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n607), .A2(G116), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(G1), .A3(new_n686), .ZN(new_n687));
  OAI22_X1  g0487(.A1(new_n687), .A2(KEYINPUT93), .B1(new_n234), .B2(new_n685), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n688), .B1(KEYINPUT93), .B2(new_n687), .ZN(new_n689));
  XOR2_X1   g0489(.A(new_n689), .B(KEYINPUT28), .Z(new_n690));
  NOR3_X1   g0490(.A1(new_n661), .A2(KEYINPUT29), .A3(new_n670), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT29), .ZN(new_n692));
  OAI21_X1  g0492(.A(KEYINPUT26), .B1(new_n654), .B2(new_n651), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n522), .A2(new_n633), .A3(new_n657), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n655), .A2(new_n649), .A3(new_n693), .A4(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n692), .B1(new_n695), .B2(new_n673), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n691), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n573), .A2(new_n634), .A3(new_n530), .A4(new_n673), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n558), .A2(new_n592), .A3(G179), .A4(new_n621), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT30), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n491), .A2(new_n498), .ZN(new_n701));
  OR3_X1    g0501(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n700), .B1(new_n699), .B2(new_n701), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n499), .A2(new_n557), .ZN(new_n705));
  OR2_X1    g0505(.A1(new_n705), .A2(KEYINPUT95), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(KEYINPUT95), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n592), .A2(new_n621), .A3(G179), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n706), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n673), .B1(new_n704), .B2(new_n709), .ZN(new_n710));
  XOR2_X1   g0510(.A(KEYINPUT94), .B(KEYINPUT31), .Z(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  OAI211_X1 g0513(.A(new_n698), .B(new_n713), .C1(KEYINPUT31), .C2(new_n710), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(G330), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n697), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n690), .B1(new_n717), .B2(G1), .ZN(G364));
  NOR2_X1   g0518(.A1(new_n229), .A2(G20), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n205), .B1(new_n719), .B2(G45), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n684), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n722), .B1(new_n679), .B2(G330), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n723), .B1(G330), .B2(new_n679), .ZN(new_n724));
  INV_X1    g0524(.A(new_n722), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n230), .A2(new_n335), .ZN(new_n726));
  AOI22_X1  g0526(.A1(new_n726), .A2(G355), .B1(new_n578), .B2(new_n230), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n257), .A2(new_n287), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n415), .A2(new_n230), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n729), .B1(G45), .B2(new_n234), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n727), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n229), .A2(new_n265), .A3(KEYINPUT96), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT96), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n733), .B1(G13), .B2(G33), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(G20), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n236), .B1(G20), .B2(new_n350), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n725), .B1(new_n731), .B2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT97), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n738), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n206), .A2(new_n387), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n744), .A2(G190), .A3(new_n460), .ZN(new_n745));
  NOR2_X1   g0545(.A1(G190), .A2(G200), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  OAI22_X1  g0547(.A1(new_n745), .A2(new_n210), .B1(new_n747), .B2(new_n202), .ZN(new_n748));
  NOR3_X1   g0548(.A1(new_n360), .A2(G179), .A3(G200), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(new_n206), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n744), .A2(G200), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(new_n360), .ZN(new_n753));
  AOI22_X1  g0553(.A1(G97), .A2(new_n751), .B1(new_n753), .B2(G50), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT32), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n206), .A2(G179), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(new_n746), .ZN(new_n757));
  INV_X1    g0557(.A(G159), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n754), .B1(new_n755), .B2(new_n759), .ZN(new_n760));
  AOI211_X1 g0560(.A(new_n748), .B(new_n760), .C1(new_n755), .C2(new_n759), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n756), .A2(new_n360), .A3(G200), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(new_n221), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n756), .A2(G190), .A3(G200), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n335), .B(new_n763), .C1(G87), .C2(new_n765), .ZN(new_n766));
  XOR2_X1   g0566(.A(new_n766), .B(KEYINPUT98), .Z(new_n767));
  NAND3_X1  g0567(.A1(new_n744), .A2(new_n360), .A3(G200), .ZN(new_n768));
  AND2_X1   g0568(.A1(new_n768), .A2(KEYINPUT99), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n768), .A2(KEYINPUT99), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  OAI211_X1 g0571(.A(new_n761), .B(new_n767), .C1(new_n214), .C2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n745), .ZN(new_n773));
  INV_X1    g0573(.A(new_n757), .ZN(new_n774));
  AOI22_X1  g0574(.A1(new_n773), .A2(G322), .B1(new_n774), .B2(G329), .ZN(new_n775));
  INV_X1    g0575(.A(G311), .ZN(new_n776));
  OAI211_X1 g0576(.A(new_n775), .B(new_n335), .C1(new_n776), .C2(new_n747), .ZN(new_n777));
  INV_X1    g0577(.A(G283), .ZN(new_n778));
  INV_X1    g0578(.A(G303), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n778), .A2(new_n762), .B1(new_n764), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n777), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n753), .A2(G326), .ZN(new_n782));
  INV_X1    g0582(.A(G294), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n782), .B1(new_n783), .B2(new_n750), .ZN(new_n784));
  OR2_X1    g0584(.A1(new_n784), .A2(KEYINPUT100), .ZN(new_n785));
  INV_X1    g0585(.A(new_n771), .ZN(new_n786));
  XNOR2_X1  g0586(.A(KEYINPUT33), .B(G317), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n784), .A2(KEYINPUT100), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n781), .A2(new_n785), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n743), .B1(new_n772), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n740), .A2(new_n741), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n737), .B(KEYINPUT101), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n742), .B(new_n793), .C1(new_n679), .C2(new_n794), .ZN(new_n795));
  AND2_X1   g0595(.A1(new_n724), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(G396));
  INV_X1    g0597(.A(KEYINPUT103), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n670), .A2(new_n379), .ZN(new_n799));
  AND3_X1   g0599(.A1(new_n389), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n799), .B1(new_n389), .B2(new_n798), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n381), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(KEYINPUT104), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  OAI211_X1 g0604(.A(KEYINPUT104), .B(new_n381), .C1(new_n800), .C2(new_n801), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(new_n661), .B2(new_n670), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n806), .A2(new_n660), .A3(new_n673), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n722), .B1(new_n810), .B2(new_n715), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n811), .B1(new_n715), .B2(new_n810), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n735), .A2(new_n738), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n722), .B1(G77), .B2(new_n814), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n335), .B1(new_n757), .B2(new_n776), .C1(new_n578), .C2(new_n747), .ZN(new_n816));
  INV_X1    g0616(.A(new_n753), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n817), .A2(new_n779), .B1(new_n762), .B2(new_n216), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n816), .B(new_n818), .C1(G107), .C2(new_n765), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(new_n778), .B2(new_n771), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n750), .A2(new_n219), .B1(new_n745), .B2(new_n783), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT102), .ZN(new_n822));
  INV_X1    g0622(.A(G132), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n415), .B1(new_n823), .B2(new_n757), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n750), .A2(new_n210), .B1(new_n764), .B2(new_n252), .ZN(new_n825));
  INV_X1    g0625(.A(new_n762), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n824), .B(new_n825), .C1(G68), .C2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n747), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n773), .A2(G143), .B1(new_n828), .B2(G159), .ZN(new_n829));
  INV_X1    g0629(.A(G137), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n829), .B1(new_n830), .B2(new_n817), .C1(new_n771), .C2(new_n259), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n827), .B1(new_n832), .B2(KEYINPUT34), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT34), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n820), .A2(new_n822), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n815), .B1(new_n836), .B2(new_n738), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n806), .B2(new_n736), .ZN(new_n838));
  AND2_X1   g0638(.A1(new_n812), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(G384));
  NOR2_X1   g0640(.A1(new_n719), .A2(new_n205), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT38), .ZN(new_n842));
  AOI21_X1  g0642(.A(KEYINPUT16), .B1(new_n429), .B2(new_n435), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n424), .B1(new_n437), .B2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n668), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n471), .A2(new_n477), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n450), .A2(new_n453), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n846), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n412), .A2(new_n420), .A3(new_n668), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(new_n844), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n466), .A2(new_n470), .A3(new_n851), .ZN(new_n852));
  AND2_X1   g0652(.A1(new_n850), .A2(new_n446), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n853), .A2(KEYINPUT37), .ZN(new_n854));
  AOI22_X1  g0654(.A1(KEYINPUT37), .A2(new_n852), .B1(new_n640), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n842), .B1(new_n849), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n852), .A2(KEYINPUT37), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n640), .A2(new_n854), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OAI211_X1 g0659(.A(KEYINPUT38), .B(new_n859), .C1(new_n478), .C2(new_n846), .ZN(new_n860));
  AND3_X1   g0660(.A1(new_n856), .A2(new_n860), .A3(KEYINPUT39), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n455), .A2(new_n668), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n645), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n863), .B1(new_n847), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(KEYINPUT37), .B1(new_n469), .B2(new_n853), .ZN(new_n866));
  AND2_X1   g0666(.A1(new_n858), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n842), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(KEYINPUT39), .B1(new_n868), .B2(new_n860), .ZN(new_n869));
  OR2_X1    g0669(.A1(new_n357), .A2(new_n670), .ZN(new_n870));
  NOR3_X1   g0670(.A1(new_n861), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n330), .A2(new_n670), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n366), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n357), .A2(new_n365), .A3(new_n872), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n389), .A2(new_n670), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n877), .B1(new_n809), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n846), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n641), .B2(new_n454), .ZN(new_n882));
  AOI21_X1  g0682(.A(KEYINPUT38), .B1(new_n882), .B2(new_n859), .ZN(new_n883));
  NOR3_X1   g0683(.A1(new_n849), .A2(new_n842), .A3(new_n855), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n880), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n885), .B1(new_n864), .B2(new_n845), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n871), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n480), .B1(new_n691), .B2(new_n696), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n888), .A2(new_n368), .A3(new_n646), .ZN(new_n889));
  XOR2_X1   g0689(.A(new_n887), .B(new_n889), .Z(new_n890));
  INV_X1    g0690(.A(G330), .ZN(new_n891));
  INV_X1    g0691(.A(new_n709), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n702), .A2(new_n703), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n670), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n711), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n710), .A2(KEYINPUT31), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n698), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n874), .A2(new_n875), .B1(new_n804), .B2(new_n805), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n900), .B1(new_n883), .B2(new_n884), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT40), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n901), .A2(KEYINPUT106), .A3(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT106), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n899), .B1(new_n856), .B2(new_n860), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n904), .B1(new_n905), .B2(KEYINPUT40), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n868), .A2(new_n860), .ZN(new_n907));
  AND3_X1   g0707(.A1(new_n897), .A2(KEYINPUT40), .A3(new_n898), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n903), .A2(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n480), .A2(new_n897), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n891), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n909), .B2(new_n910), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n841), .B1(new_n890), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n890), .B2(new_n912), .ZN(new_n914));
  NAND4_X1  g0714(.A1(new_n235), .A2(G77), .A3(new_n433), .A4(new_n431), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n253), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n916), .A2(G1), .A3(new_n229), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n507), .A2(new_n509), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  OR2_X1    g0719(.A1(new_n919), .A2(KEYINPUT35), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(KEYINPUT35), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n920), .A2(new_n921), .A3(G116), .A4(new_n237), .ZN(new_n922));
  XNOR2_X1  g0722(.A(KEYINPUT105), .B(KEYINPUT36), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n922), .B(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n914), .A2(new_n917), .A3(new_n924), .ZN(new_n925));
  XOR2_X1   g0725(.A(new_n925), .B(KEYINPUT107), .Z(G367));
  INV_X1    g0726(.A(new_n672), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n530), .B1(new_n523), .B2(new_n673), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n522), .A2(new_n670), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(KEYINPUT42), .B1(new_n927), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n571), .B1(new_n528), .B2(new_n529), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n673), .B1(new_n933), .B2(new_n522), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NOR3_X1   g0735(.A1(new_n927), .A2(new_n931), .A3(KEYINPUT42), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT43), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n673), .A2(new_n632), .ZN(new_n938));
  MUX2_X1   g0738(.A(new_n651), .B(new_n649), .S(new_n938), .Z(new_n939));
  OAI22_X1  g0739(.A1(new_n935), .A2(new_n936), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n937), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n940), .B(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n681), .A2(new_n931), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n942), .B1(KEYINPUT108), .B2(new_n943), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n943), .B(KEYINPUT108), .Z(new_n945));
  OR2_X1    g0745(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n684), .B(KEYINPUT41), .Z(new_n947));
  NAND2_X1  g0747(.A1(new_n674), .A2(new_n930), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n948), .B(KEYINPUT45), .Z(new_n949));
  NOR2_X1   g0749(.A1(new_n674), .A2(new_n930), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT44), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(new_n681), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n676), .A2(new_n671), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n927), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(new_n680), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n956), .A2(new_n716), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n953), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n947), .B1(new_n958), .B2(new_n717), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n944), .B(new_n946), .C1(new_n959), .C2(new_n721), .ZN(new_n960));
  INV_X1    g0760(.A(new_n794), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n939), .A2(new_n961), .ZN(new_n962));
  AOI211_X1 g0762(.A(new_n738), .B(new_n737), .C1(new_n230), .C2(new_n375), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n247), .A2(new_n729), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n725), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n750), .A2(new_n214), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(G77), .B2(new_n826), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n335), .B1(new_n773), .B2(G150), .ZN(new_n968));
  AOI22_X1  g0768(.A1(G50), .A2(new_n828), .B1(new_n774), .B2(G137), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n753), .A2(G143), .B1(new_n765), .B2(G58), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n967), .A2(new_n968), .A3(new_n969), .A4(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n771), .A2(new_n758), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n415), .B1(new_n753), .B2(G311), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n751), .A2(G107), .B1(new_n826), .B2(G97), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n973), .B(new_n974), .C1(new_n771), .C2(new_n783), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n773), .A2(new_n586), .B1(new_n774), .B2(G317), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n765), .A2(KEYINPUT46), .A3(G116), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT46), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n764), .B2(new_n578), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n828), .A2(G283), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n976), .A2(new_n977), .A3(new_n979), .A4(new_n980), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n971), .A2(new_n972), .B1(new_n975), .B2(new_n981), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT109), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n983), .B(KEYINPUT47), .Z(new_n984));
  OAI211_X1 g0784(.A(new_n962), .B(new_n965), .C1(new_n984), .C2(new_n743), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n960), .A2(new_n985), .ZN(G387));
  NOR2_X1   g0786(.A1(new_n957), .A2(new_n685), .ZN(new_n987));
  INV_X1    g0787(.A(new_n956), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n987), .B1(new_n717), .B2(new_n988), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n786), .A2(new_n264), .B1(G68), .B2(new_n828), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT112), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n415), .B1(new_n745), .B2(new_n252), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n612), .A2(new_n750), .B1(new_n219), .B2(new_n762), .ZN(new_n993));
  AOI211_X1 g0793(.A(new_n992), .B(new_n993), .C1(G159), .C2(new_n753), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n764), .A2(new_n202), .B1(new_n757), .B2(new_n259), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT111), .Z(new_n996));
  NAND3_X1  g0796(.A1(new_n991), .A2(new_n994), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n753), .A2(G322), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n773), .A2(G317), .B1(new_n828), .B2(new_n586), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n998), .B(new_n999), .C1(new_n771), .C2(new_n776), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT48), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n751), .A2(G283), .B1(new_n765), .B2(G294), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT49), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(KEYINPUT113), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n415), .B1(G326), .B2(new_n774), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n1007), .B(new_n1008), .C1(new_n578), .C2(new_n762), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1006), .A2(KEYINPUT113), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n997), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n738), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n676), .A2(new_n961), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n686), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n726), .A2(new_n1014), .B1(new_n221), .B2(new_n230), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n244), .A2(new_n287), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n263), .A2(G50), .ZN(new_n1017));
  XOR2_X1   g0817(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n1018));
  XNOR2_X1  g0818(.A(new_n1017), .B(new_n1018), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n686), .B(new_n287), .C1(new_n214), .C2(new_n202), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n729), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1015), .B1(new_n1016), .B2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n725), .B1(new_n1022), .B2(new_n739), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1012), .A2(new_n1013), .A3(new_n1023), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n989), .B(new_n1024), .C1(new_n720), .C2(new_n956), .ZN(G393));
  AOI21_X1  g0825(.A(new_n685), .B1(new_n953), .B2(new_n957), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n957), .B2(new_n953), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n817), .A2(new_n259), .B1(new_n758), .B2(new_n745), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT51), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n214), .A2(new_n764), .B1(new_n762), .B2(new_n216), .ZN(new_n1030));
  INV_X1    g0830(.A(G143), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n415), .B1(new_n757), .B2(new_n1031), .C1(new_n263), .C2(new_n747), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n1030), .B(new_n1032), .C1(G77), .C2(new_n751), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1029), .B(new_n1033), .C1(new_n252), .C2(new_n771), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT114), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(G317), .A2(new_n753), .B1(new_n773), .B2(G311), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT52), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n786), .A2(new_n586), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n335), .B1(new_n747), .B2(new_n783), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(G322), .B2(new_n774), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n764), .A2(new_n778), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n763), .B(new_n1042), .C1(G116), .C2(new_n751), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1039), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1036), .B1(new_n1038), .B2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n738), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n251), .A2(new_n729), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1048), .B(new_n739), .C1(new_n219), .C2(new_n231), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1047), .A2(new_n722), .A3(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(new_n931), .B2(new_n737), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(new_n953), .B2(new_n721), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1027), .A2(new_n1052), .ZN(G390));
  NAND3_X1  g0853(.A1(new_n897), .A2(new_n898), .A3(G330), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n870), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n880), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT39), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n862), .B1(new_n641), .B2(new_n645), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n858), .A2(new_n866), .ZN(new_n1060));
  AOI21_X1  g0860(.A(KEYINPUT38), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1058), .B1(new_n1061), .B2(new_n884), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n856), .A2(new_n860), .A3(KEYINPUT39), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1057), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT115), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n876), .B(new_n1065), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n695), .A2(new_n806), .A3(new_n673), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(new_n879), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1069));
  AND3_X1   g0869(.A1(new_n1069), .A2(new_n907), .A3(new_n870), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1055), .B1(new_n1064), .B2(new_n1070), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n861), .A2(new_n869), .B1(new_n880), .B2(new_n1056), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1069), .A2(new_n907), .A3(new_n870), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n714), .A2(G330), .A3(new_n806), .A4(new_n876), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n480), .A2(G330), .A3(new_n897), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n888), .A2(new_n1076), .A3(new_n368), .A4(new_n646), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n809), .A2(new_n879), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n714), .A2(G330), .A3(new_n806), .ZN(new_n1079));
  AND2_X1   g0879(.A1(new_n1079), .A2(new_n877), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1078), .B1(new_n1080), .B2(new_n1055), .ZN(new_n1081));
  AND2_X1   g0881(.A1(new_n1067), .A2(new_n879), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n897), .A2(G330), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1083), .A2(new_n807), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1082), .B(new_n1074), .C1(new_n1084), .C2(new_n1066), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1077), .B1(new_n1081), .B2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1071), .A2(new_n1075), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(KEYINPUT116), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT116), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n1071), .A2(new_n1075), .A3(new_n1086), .A4(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  AND2_X1   g0891(.A1(new_n1071), .A2(new_n1075), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1091), .B(new_n684), .C1(new_n1092), .C2(new_n1086), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n735), .B1(new_n861), .B2(new_n869), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n722), .B1(new_n264), .B2(new_n814), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n753), .A2(G128), .B1(new_n826), .B2(G50), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n1096), .B1(new_n758), .B2(new_n750), .C1(new_n771), .C2(new_n830), .ZN(new_n1097));
  XOR2_X1   g0897(.A(KEYINPUT54), .B(G143), .Z(new_n1098));
  AOI22_X1  g0898(.A1(new_n828), .A2(new_n1098), .B1(new_n774), .B2(G125), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n335), .B1(new_n773), .B2(G132), .ZN(new_n1100));
  OR3_X1    g0900(.A1(new_n764), .A2(KEYINPUT53), .A3(new_n259), .ZN(new_n1101));
  OAI21_X1  g0901(.A(KEYINPUT53), .B1(new_n764), .B2(new_n259), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .A4(new_n1102), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n771), .A2(new_n221), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(G77), .A2(new_n751), .B1(new_n753), .B2(G283), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n297), .B1(new_n828), .B2(G97), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n773), .A2(G116), .B1(new_n774), .B2(G294), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n765), .A2(G87), .B1(new_n826), .B2(G68), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .A4(new_n1108), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n1097), .A2(new_n1103), .B1(new_n1104), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT117), .ZN(new_n1111));
  OR2_X1    g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n743), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1095), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n1092), .A2(new_n721), .B1(new_n1094), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1093), .A2(new_n1115), .ZN(G378));
  AOI21_X1  g0916(.A(new_n891), .B1(new_n907), .B2(new_n908), .ZN(new_n1117));
  AOI21_X1  g0917(.A(KEYINPUT106), .B1(new_n901), .B2(new_n902), .ZN(new_n1118));
  NOR3_X1   g0918(.A1(new_n905), .A2(new_n904), .A3(KEYINPUT40), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1117), .B(KEYINPUT118), .C1(new_n1118), .C2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n636), .A2(new_n368), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n277), .A2(new_n845), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1121), .B(new_n1122), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1124));
  XOR2_X1   g0924(.A(new_n1123), .B(new_n1124), .Z(new_n1125));
  NAND2_X1  g0925(.A1(new_n1120), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n907), .A2(new_n908), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(G330), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(new_n903), .B2(new_n906), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1129), .A2(KEYINPUT118), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1126), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n887), .ZN(new_n1132));
  NOR3_X1   g0932(.A1(new_n1125), .A2(new_n1129), .A3(KEYINPUT118), .ZN(new_n1133));
  NOR3_X1   g0933(.A1(new_n1131), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1126), .A2(new_n1130), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1117), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT118), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1138), .A2(new_n1120), .A3(new_n1125), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n887), .B1(new_n1135), .B2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1077), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1141));
  NOR3_X1   g0941(.A1(new_n1134), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(KEYINPUT119), .B1(new_n1142), .B2(KEYINPUT57), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1077), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1091), .A2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1132), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1135), .A2(new_n1139), .A3(new_n887), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1145), .A2(new_n1146), .A3(KEYINPUT57), .A4(new_n1147), .ZN(new_n1148));
  AND2_X1   g0948(.A1(new_n1148), .A2(new_n684), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT119), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT57), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1150), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1143), .A2(new_n1149), .A3(new_n1153), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n817), .A2(new_n578), .B1(new_n762), .B2(new_n210), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n966), .B(new_n1155), .C1(G77), .C2(new_n765), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n745), .A2(new_n221), .B1(new_n757), .B2(new_n778), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n425), .A2(new_n284), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n1157), .B(new_n1158), .C1(new_n375), .C2(new_n828), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1156), .B(new_n1159), .C1(new_n219), .C2(new_n771), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT58), .ZN(new_n1161));
  AOI21_X1  g0961(.A(G50), .B1(new_n265), .B2(new_n284), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n1160), .A2(new_n1161), .B1(new_n1158), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(G128), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n745), .A2(new_n1164), .B1(new_n747), .B2(new_n830), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(G150), .B2(new_n751), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n753), .A2(G125), .B1(new_n765), .B2(new_n1098), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1166), .B(new_n1167), .C1(new_n771), .C2(new_n823), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1168), .A2(KEYINPUT59), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(KEYINPUT59), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n826), .A2(G159), .ZN(new_n1171));
  AOI211_X1 g0971(.A(G33), .B(G41), .C1(new_n774), .C2(G124), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  OAI221_X1 g0973(.A(new_n1163), .B1(new_n1161), .B2(new_n1160), .C1(new_n1169), .C2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(new_n738), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1175), .B(new_n722), .C1(G50), .C2(new_n814), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(new_n1125), .B2(new_n735), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1134), .A2(new_n1140), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1177), .B1(new_n1178), .B2(new_n721), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1154), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT120), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1184));
  AND2_X1   g0984(.A1(new_n1183), .A2(new_n1184), .ZN(G375));
  NOR2_X1   g0985(.A1(new_n1086), .A2(new_n947), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1081), .A2(new_n1085), .A3(new_n1077), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1081), .A2(new_n1085), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1066), .A2(new_n736), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1190), .B(KEYINPUT121), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n814), .A2(G68), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n817), .A2(new_n823), .B1(new_n252), .B2(new_n750), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(G159), .B2(new_n765), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n786), .A2(new_n1098), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n747), .A2(new_n259), .B1(new_n757), .B2(new_n1164), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(G137), .B2(new_n773), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n425), .B1(G58), .B2(new_n826), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1194), .A2(new_n1195), .A3(new_n1197), .A4(new_n1198), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n817), .A2(new_n783), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n335), .B1(new_n747), .B2(new_n221), .C1(new_n778), .C2(new_n745), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n612), .A2(new_n750), .B1(new_n202), .B2(new_n762), .ZN(new_n1202));
  NOR3_X1   g1002(.A1(new_n1200), .A2(new_n1201), .A3(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n578), .B2(new_n771), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n764), .A2(new_n219), .B1(new_n757), .B2(new_n779), .ZN(new_n1205));
  XOR2_X1   g1005(.A(new_n1205), .B(KEYINPUT122), .Z(new_n1206));
  OAI21_X1  g1006(.A(new_n1199), .B1(new_n1204), .B2(new_n1206), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n725), .B(new_n1192), .C1(new_n1207), .C2(new_n738), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n721), .A2(new_n1189), .B1(new_n1191), .B2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1188), .A2(new_n1209), .ZN(G381));
  INV_X1    g1010(.A(G390), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(new_n839), .ZN(new_n1212));
  OR2_X1    g1012(.A1(G393), .A2(G396), .ZN(new_n1213));
  NOR4_X1   g1013(.A1(new_n1212), .A2(G387), .A3(G381), .A4(new_n1213), .ZN(new_n1214));
  XOR2_X1   g1014(.A(new_n1214), .B(KEYINPUT123), .Z(new_n1215));
  AOI21_X1  g1015(.A(G378), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n1215), .A2(KEYINPUT124), .A3(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(KEYINPUT124), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1218));
  OR2_X1    g1018(.A1(new_n1217), .A2(new_n1218), .ZN(G407));
  NAND2_X1  g1019(.A1(new_n1216), .A2(new_n669), .ZN(new_n1220));
  OAI211_X1 g1020(.A(G213), .B(new_n1220), .C1(new_n1217), .C2(new_n1218), .ZN(G409));
  XNOR2_X1  g1021(.A(G393), .B(new_n796), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n960), .A2(new_n985), .A3(G390), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(G390), .B1(new_n960), .B2(new_n985), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1223), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1226), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1228), .A2(new_n1222), .A3(new_n1224), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1227), .A2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1154), .A2(G378), .A3(new_n1179), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1179), .B1(new_n947), .B2(new_n1150), .ZN(new_n1232));
  INV_X1    g1032(.A(G378), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1231), .A2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n669), .A2(G213), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT60), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1187), .B1(new_n1086), .B2(new_n1237), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1081), .A2(KEYINPUT60), .A3(new_n1077), .A4(new_n1085), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1238), .A2(new_n684), .A3(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(new_n1209), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(new_n1241), .B(G384), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1235), .A2(new_n1236), .A3(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(KEYINPUT62), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT125), .ZN(new_n1246));
  INV_X1    g1046(.A(G2897), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1236), .A2(new_n1247), .ZN(new_n1248));
  OR3_X1    g1048(.A1(new_n1242), .A2(new_n1246), .A3(new_n1248), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1248), .B1(new_n1242), .B2(new_n1246), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n1249), .A2(new_n1250), .B1(new_n1246), .B2(new_n1242), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1245), .A2(new_n1251), .ZN(new_n1252));
  XOR2_X1   g1052(.A(KEYINPUT127), .B(KEYINPUT61), .Z(new_n1253));
  NAND3_X1  g1053(.A1(new_n1244), .A2(new_n1252), .A3(new_n1253), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1243), .A2(KEYINPUT62), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1230), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT61), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1227), .A2(new_n1229), .A3(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1258), .B1(new_n1245), .B2(new_n1251), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT126), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n1231), .A2(new_n1234), .B1(G213), .B2(new_n669), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT63), .ZN(new_n1262));
  AND3_X1   g1062(.A1(new_n1261), .A2(new_n1262), .A3(new_n1242), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1262), .B1(new_n1261), .B2(new_n1242), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1259), .B(new_n1260), .C1(new_n1263), .C2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1243), .A2(KEYINPUT63), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1261), .A2(new_n1262), .A3(new_n1242), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1260), .B1(new_n1269), .B2(new_n1259), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1256), .B1(new_n1266), .B2(new_n1270), .ZN(G405));
  AOI21_X1  g1071(.A(new_n1233), .B1(new_n1154), .B2(new_n1179), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1216), .A2(new_n1272), .ZN(new_n1273));
  XNOR2_X1  g1073(.A(new_n1230), .B(new_n1242), .ZN(new_n1274));
  XNOR2_X1  g1074(.A(new_n1273), .B(new_n1274), .ZN(G402));
endmodule


