

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733;

  NAND2_X1 U369 ( .A1(n527), .A2(n492), .ZN(n687) );
  OR2_X1 U370 ( .A1(n633), .A2(n447), .ZN(n452) );
  OR2_X1 U371 ( .A1(n704), .A2(G902), .ZN(n356) );
  OR2_X1 U372 ( .A1(n699), .A2(G902), .ZN(n406) );
  XNOR2_X1 U373 ( .A(n436), .B(n383), .ZN(n455) );
  XNOR2_X2 U374 ( .A(n549), .B(n548), .ZN(n369) );
  XNOR2_X1 U375 ( .A(n346), .B(KEYINPUT69), .ZN(n537) );
  NAND2_X1 U376 ( .A1(n513), .A2(n514), .ZN(n346) );
  AND2_X1 U377 ( .A1(n494), .A2(n550), .ZN(n645) );
  AND2_X1 U378 ( .A1(n592), .A2(n562), .ZN(n564) );
  AND2_X4 U379 ( .A1(n606), .A2(n607), .ZN(n698) );
  NOR2_X2 U380 ( .A1(n655), .A2(n487), .ZN(n491) );
  NAND2_X2 U381 ( .A1(n485), .A2(n657), .ZN(n655) );
  OR2_X2 U382 ( .A1(n572), .A2(n648), .ZN(n540) );
  INV_X1 U383 ( .A(n581), .ZN(n485) );
  NOR2_X2 U384 ( .A1(n557), .A2(n556), .ZN(n559) );
  XNOR2_X2 U385 ( .A(n496), .B(n495), .ZN(n557) );
  XNOR2_X2 U386 ( .A(n559), .B(n558), .ZN(n592) );
  INV_X2 U387 ( .A(G953), .ZN(n723) );
  NOR2_X1 U388 ( .A1(n645), .A2(n557), .ZN(n497) );
  INV_X1 U389 ( .A(n516), .ZN(n544) );
  NAND2_X1 U390 ( .A1(n372), .A2(n370), .ZN(n606) );
  NAND2_X1 U391 ( .A1(n371), .A2(KEYINPUT83), .ZN(n370) );
  NAND2_X1 U392 ( .A1(n547), .A2(n546), .ZN(n549) );
  XNOR2_X1 U393 ( .A(n600), .B(KEYINPUT45), .ZN(n715) );
  NOR2_X1 U394 ( .A1(n731), .A2(n621), .ZN(n578) );
  AND2_X1 U395 ( .A1(n687), .A2(n497), .ZN(n503) );
  OR2_X1 U396 ( .A1(n589), .A2(n648), .ZN(n489) );
  OR2_X1 U397 ( .A1(n588), .A2(n486), .ZN(n487) );
  BUF_X1 U398 ( .A(n588), .Z(n348) );
  XNOR2_X1 U399 ( .A(n482), .B(G469), .ZN(n588) );
  XNOR2_X1 U400 ( .A(G116), .B(G113), .ZN(n431) );
  XNOR2_X1 U401 ( .A(KEYINPUT66), .B(G101), .ZN(n461) );
  XNOR2_X1 U402 ( .A(KEYINPUT3), .B(G119), .ZN(n430) );
  AND2_X2 U403 ( .A1(n722), .A2(n715), .ZN(n347) );
  INV_X1 U404 ( .A(n347), .ZN(n640) );
  NAND2_X1 U405 ( .A1(n581), .A2(n428), .ZN(n429) );
  XNOR2_X1 U406 ( .A(n480), .B(n479), .ZN(n721) );
  INV_X1 U407 ( .A(G902), .ZN(n449) );
  INV_X1 U408 ( .A(KEYINPUT70), .ZN(n359) );
  NAND2_X1 U409 ( .A1(n498), .A2(n662), .ZN(n358) );
  XNOR2_X1 U410 ( .A(KEYINPUT0), .B(KEYINPUT90), .ZN(n558) );
  XNOR2_X1 U411 ( .A(n481), .B(n721), .ZN(n694) );
  NOR2_X1 U412 ( .A1(n678), .A2(n677), .ZN(n366) );
  INV_X1 U413 ( .A(KEYINPUT47), .ZN(n360) );
  AND2_X1 U414 ( .A1(n512), .A2(n511), .ZN(n513) );
  NAND2_X1 U415 ( .A1(G234), .A2(G237), .ZN(n421) );
  XOR2_X1 U416 ( .A(KEYINPUT68), .B(KEYINPUT8), .Z(n378) );
  XOR2_X1 U417 ( .A(G137), .B(G140), .Z(n478) );
  XNOR2_X1 U418 ( .A(n588), .B(KEYINPUT1), .ZN(n570) );
  INV_X1 U419 ( .A(G237), .ZN(n448) );
  XNOR2_X1 U420 ( .A(G116), .B(G107), .ZN(n381) );
  XNOR2_X1 U421 ( .A(G131), .B(G140), .ZN(n398) );
  XNOR2_X1 U422 ( .A(G110), .B(G107), .ZN(n434) );
  INV_X1 U423 ( .A(KEYINPUT76), .ZN(n602) );
  XNOR2_X1 U424 ( .A(n376), .B(n552), .ZN(n601) );
  XNOR2_X1 U425 ( .A(n358), .B(n499), .ZN(n502) );
  XNOR2_X1 U426 ( .A(n355), .B(KEYINPUT25), .ZN(n354) );
  NAND2_X1 U427 ( .A1(n419), .A2(G217), .ZN(n355) );
  XNOR2_X1 U428 ( .A(n367), .B(n352), .ZN(n731) );
  BUF_X1 U429 ( .A(n530), .Z(n617) );
  XNOR2_X1 U430 ( .A(n696), .B(n695), .ZN(n697) );
  XNOR2_X1 U431 ( .A(n694), .B(n693), .ZN(n695) );
  INV_X1 U432 ( .A(KEYINPUT53), .ZN(n363) );
  XNOR2_X1 U433 ( .A(n366), .B(KEYINPUT124), .ZN(n365) );
  XNOR2_X1 U434 ( .A(n362), .B(KEYINPUT33), .ZN(n644) );
  AND2_X1 U435 ( .A1(n524), .A2(n507), .ZN(n349) );
  AND2_X1 U436 ( .A1(n614), .A2(KEYINPUT2), .ZN(n350) );
  XNOR2_X1 U437 ( .A(KEYINPUT34), .B(KEYINPUT79), .ZN(n351) );
  XOR2_X1 U438 ( .A(KEYINPUT85), .B(KEYINPUT35), .Z(n352) );
  XOR2_X1 U439 ( .A(KEYINPUT88), .B(KEYINPUT48), .Z(n353) );
  XNOR2_X1 U440 ( .A(KEYINPUT15), .B(G902), .ZN(n604) );
  XNOR2_X2 U441 ( .A(n356), .B(n354), .ZN(n581) );
  XNOR2_X1 U442 ( .A(n357), .B(n416), .ZN(n704) );
  XNOR2_X1 U443 ( .A(n409), .B(n410), .ZN(n357) );
  XNOR2_X2 U444 ( .A(n429), .B(n359), .ZN(n498) );
  AND2_X2 U445 ( .A1(n490), .A2(n491), .ZN(n527) );
  NAND2_X1 U446 ( .A1(n687), .A2(n360), .ZN(n504) );
  INV_X1 U447 ( .A(n570), .ZN(n575) );
  NAND2_X1 U448 ( .A1(n575), .A2(n571), .ZN(n586) );
  NAND2_X1 U449 ( .A1(n361), .A2(n575), .ZN(n362) );
  NOR2_X1 U450 ( .A1(n655), .A2(n572), .ZN(n361) );
  XNOR2_X1 U451 ( .A(n364), .B(n363), .ZN(G75) );
  NAND2_X1 U452 ( .A1(n365), .A2(n723), .ZN(n364) );
  NAND2_X1 U453 ( .A1(n368), .A2(n574), .ZN(n367) );
  XNOR2_X1 U454 ( .A(n573), .B(n351), .ZN(n368) );
  NAND2_X1 U455 ( .A1(n369), .A2(n350), .ZN(n376) );
  AND2_X2 U456 ( .A1(n369), .A2(n614), .ZN(n722) );
  NAND2_X1 U457 ( .A1(n347), .A2(n447), .ZN(n371) );
  NAND2_X1 U458 ( .A1(n373), .A2(n447), .ZN(n372) );
  NAND2_X1 U459 ( .A1(n375), .A2(n374), .ZN(n373) );
  INV_X1 U460 ( .A(KEYINPUT2), .ZN(n374) );
  NAND2_X1 U461 ( .A1(n347), .A2(n605), .ZN(n375) );
  NOR2_X2 U462 ( .A1(G953), .A2(G237), .ZN(n456) );
  INV_X1 U463 ( .A(KEYINPUT84), .ZN(n552) );
  INV_X1 U464 ( .A(n478), .ZN(n479) );
  NOR2_X1 U465 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U466 ( .A(n415), .B(n414), .ZN(n416) );
  INV_X1 U467 ( .A(n707), .ZN(n611) );
  BUF_X1 U468 ( .A(n622), .Z(n625) );
  XOR2_X1 U469 ( .A(KEYINPUT105), .B(KEYINPUT7), .Z(n380) );
  NAND2_X1 U470 ( .A1(G234), .A2(n723), .ZN(n377) );
  XNOR2_X1 U471 ( .A(n378), .B(n377), .ZN(n411) );
  NAND2_X1 U472 ( .A1(G217), .A2(n411), .ZN(n379) );
  XNOR2_X1 U473 ( .A(n380), .B(n379), .ZN(n387) );
  XOR2_X1 U474 ( .A(KEYINPUT9), .B(G122), .Z(n382) );
  XNOR2_X1 U475 ( .A(n382), .B(n381), .ZN(n385) );
  XNOR2_X2 U476 ( .A(G143), .B(G128), .ZN(n436) );
  INV_X1 U477 ( .A(G134), .ZN(n383) );
  INV_X1 U478 ( .A(n455), .ZN(n384) );
  XNOR2_X1 U479 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U480 ( .A(n387), .B(n386), .ZN(n608) );
  NAND2_X1 U481 ( .A1(n608), .A2(n449), .ZN(n389) );
  XNOR2_X1 U482 ( .A(G478), .B(KEYINPUT106), .ZN(n388) );
  XNOR2_X1 U483 ( .A(n389), .B(n388), .ZN(n493) );
  INV_X1 U484 ( .A(n493), .ZN(n407) );
  NAND2_X1 U485 ( .A1(n456), .A2(G214), .ZN(n390) );
  XNOR2_X1 U486 ( .A(n390), .B(KEYINPUT102), .ZN(n392) );
  XNOR2_X1 U487 ( .A(KEYINPUT12), .B(KEYINPUT101), .ZN(n391) );
  XNOR2_X1 U488 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X2 U489 ( .A(G146), .B(G125), .ZN(n438) );
  XNOR2_X2 U490 ( .A(n438), .B(KEYINPUT10), .ZN(n720) );
  XNOR2_X1 U491 ( .A(n393), .B(n720), .ZN(n402) );
  INV_X1 U492 ( .A(G113), .ZN(n394) );
  XNOR2_X1 U493 ( .A(n394), .B(G122), .ZN(n396) );
  XNOR2_X1 U494 ( .A(G143), .B(G104), .ZN(n395) );
  XNOR2_X1 U495 ( .A(n396), .B(n395), .ZN(n400) );
  XNOR2_X1 U496 ( .A(KEYINPUT103), .B(KEYINPUT11), .ZN(n397) );
  XNOR2_X1 U497 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U498 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U499 ( .A(n402), .B(n401), .ZN(n699) );
  XNOR2_X1 U500 ( .A(KEYINPUT13), .B(G475), .ZN(n404) );
  INV_X1 U501 ( .A(KEYINPUT104), .ZN(n403) );
  XNOR2_X1 U502 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U503 ( .A(n406), .B(n405), .ZN(n517) );
  NAND2_X1 U504 ( .A1(n407), .A2(n517), .ZN(n408) );
  XNOR2_X2 U505 ( .A(n408), .B(KEYINPUT107), .ZN(n530) );
  XOR2_X1 U506 ( .A(G110), .B(n478), .Z(n410) );
  XNOR2_X1 U507 ( .A(n720), .B(G128), .ZN(n409) );
  AND2_X1 U508 ( .A1(G221), .A2(n411), .ZN(n415) );
  XOR2_X1 U509 ( .A(KEYINPUT98), .B(KEYINPUT23), .Z(n413) );
  XNOR2_X1 U510 ( .A(G119), .B(KEYINPUT24), .ZN(n412) );
  XNOR2_X1 U511 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U512 ( .A(KEYINPUT99), .B(KEYINPUT20), .Z(n418) );
  NAND2_X1 U513 ( .A1(G234), .A2(n604), .ZN(n417) );
  XNOR2_X1 U514 ( .A(n418), .B(n417), .ZN(n419) );
  NAND2_X1 U515 ( .A1(n419), .A2(G221), .ZN(n420) );
  XOR2_X1 U516 ( .A(n420), .B(KEYINPUT21), .Z(n657) );
  XNOR2_X1 U517 ( .A(n421), .B(KEYINPUT14), .ZN(n424) );
  NAND2_X1 U518 ( .A1(n424), .A2(G952), .ZN(n423) );
  INV_X1 U519 ( .A(KEYINPUT96), .ZN(n422) );
  XNOR2_X1 U520 ( .A(n423), .B(n422), .ZN(n672) );
  AND2_X1 U521 ( .A1(n672), .A2(n723), .ZN(n555) );
  NAND2_X1 U522 ( .A1(G902), .A2(n424), .ZN(n553) );
  OR2_X1 U523 ( .A1(n723), .A2(n553), .ZN(n425) );
  NOR2_X1 U524 ( .A1(n425), .A2(G900), .ZN(n426) );
  NOR2_X1 U525 ( .A1(n555), .A2(n426), .ZN(n486) );
  INV_X1 U526 ( .A(n486), .ZN(n427) );
  AND2_X1 U527 ( .A1(n657), .A2(n427), .ZN(n428) );
  XNOR2_X1 U528 ( .A(n431), .B(n430), .ZN(n462) );
  XNOR2_X1 U529 ( .A(KEYINPUT74), .B(KEYINPUT16), .ZN(n432) );
  XNOR2_X1 U530 ( .A(n432), .B(G122), .ZN(n433) );
  XNOR2_X1 U531 ( .A(n462), .B(n433), .ZN(n435) );
  XNOR2_X1 U532 ( .A(n434), .B(G104), .ZN(n474) );
  XNOR2_X1 U533 ( .A(n435), .B(n474), .ZN(n708) );
  XNOR2_X1 U534 ( .A(n436), .B(n461), .ZN(n440) );
  XNOR2_X1 U535 ( .A(KEYINPUT78), .B(KEYINPUT91), .ZN(n437) );
  XNOR2_X1 U536 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U537 ( .A(n440), .B(n439), .ZN(n445) );
  XOR2_X1 U538 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n443) );
  NAND2_X1 U539 ( .A1(G224), .A2(n723), .ZN(n441) );
  XNOR2_X1 U540 ( .A(n441), .B(KEYINPUT4), .ZN(n442) );
  XNOR2_X1 U541 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U542 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U543 ( .A(n708), .B(n446), .ZN(n633) );
  INV_X1 U544 ( .A(n604), .ZN(n447) );
  NAND2_X1 U545 ( .A1(n449), .A2(n448), .ZN(n470) );
  NAND2_X1 U546 ( .A1(n470), .A2(G210), .ZN(n450) );
  XNOR2_X1 U547 ( .A(n450), .B(KEYINPUT95), .ZN(n451) );
  XNOR2_X2 U548 ( .A(n452), .B(n451), .ZN(n516) );
  AND2_X1 U549 ( .A1(n498), .A2(n516), .ZN(n453) );
  NAND2_X1 U550 ( .A1(n530), .A2(n453), .ZN(n471) );
  XNOR2_X1 U551 ( .A(KEYINPUT4), .B(G131), .ZN(n454) );
  XNOR2_X2 U552 ( .A(n455), .B(n454), .ZN(n480) );
  NAND2_X1 U553 ( .A1(n456), .A2(G210), .ZN(n457) );
  XNOR2_X1 U554 ( .A(n457), .B(KEYINPUT100), .ZN(n459) );
  XNOR2_X1 U555 ( .A(KEYINPUT5), .B(G137), .ZN(n458) );
  XNOR2_X1 U556 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U557 ( .A(n480), .B(n460), .ZN(n465) );
  XNOR2_X1 U558 ( .A(n461), .B(G146), .ZN(n477) );
  INV_X1 U559 ( .A(n462), .ZN(n463) );
  XNOR2_X1 U560 ( .A(n477), .B(n463), .ZN(n464) );
  XNOR2_X1 U561 ( .A(n465), .B(n464), .ZN(n626) );
  OR2_X2 U562 ( .A1(n626), .A2(G902), .ZN(n467) );
  XNOR2_X1 U563 ( .A(KEYINPUT73), .B(G472), .ZN(n466) );
  XNOR2_X2 U564 ( .A(n467), .B(n466), .ZN(n589) );
  INV_X1 U565 ( .A(n589), .ZN(n469) );
  XNOR2_X1 U566 ( .A(KEYINPUT108), .B(KEYINPUT6), .ZN(n468) );
  XNOR2_X1 U567 ( .A(n469), .B(n468), .ZN(n572) );
  NAND2_X1 U568 ( .A1(n470), .A2(G214), .ZN(n519) );
  INV_X1 U569 ( .A(n519), .ZN(n648) );
  NOR2_X2 U570 ( .A1(n471), .A2(n540), .ZN(n472) );
  XNOR2_X1 U571 ( .A(n472), .B(KEYINPUT36), .ZN(n483) );
  NAND2_X1 U572 ( .A1(G227), .A2(n723), .ZN(n473) );
  XOR2_X1 U573 ( .A(n473), .B(KEYINPUT77), .Z(n475) );
  XNOR2_X1 U574 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U575 ( .A(n477), .B(n476), .ZN(n481) );
  NOR2_X1 U576 ( .A1(G902), .A2(n694), .ZN(n482) );
  XNOR2_X1 U577 ( .A(n570), .B(KEYINPUT93), .ZN(n566) );
  NAND2_X1 U578 ( .A1(n483), .A2(n566), .ZN(n484) );
  XNOR2_X2 U579 ( .A(n484), .B(KEYINPUT117), .ZN(n622) );
  INV_X1 U580 ( .A(n622), .ZN(n514) );
  XNOR2_X1 U581 ( .A(KEYINPUT111), .B(KEYINPUT30), .ZN(n488) );
  XNOR2_X1 U582 ( .A(n489), .B(n488), .ZN(n490) );
  AND2_X1 U583 ( .A1(n493), .A2(n517), .ZN(n574) );
  AND2_X1 U584 ( .A1(n574), .A2(n516), .ZN(n492) );
  INV_X1 U585 ( .A(n530), .ZN(n494) );
  OR2_X1 U586 ( .A1(n407), .A2(n517), .ZN(n550) );
  NAND2_X1 U587 ( .A1(n516), .A2(n519), .ZN(n496) );
  INV_X1 U588 ( .A(KEYINPUT19), .ZN(n495) );
  INV_X1 U589 ( .A(n557), .ZN(n507) );
  INV_X1 U590 ( .A(n589), .ZN(n662) );
  XNOR2_X1 U591 ( .A(KEYINPUT113), .B(KEYINPUT28), .ZN(n499) );
  INV_X1 U592 ( .A(KEYINPUT112), .ZN(n500) );
  XNOR2_X1 U593 ( .A(n348), .B(n500), .ZN(n501) );
  AND2_X2 U594 ( .A1(n502), .A2(n501), .ZN(n524) );
  NAND2_X1 U595 ( .A1(n503), .A2(n524), .ZN(n505) );
  NAND2_X1 U596 ( .A1(n505), .A2(n504), .ZN(n506) );
  XNOR2_X1 U597 ( .A(n506), .B(KEYINPUT82), .ZN(n512) );
  INV_X1 U598 ( .A(n645), .ZN(n593) );
  XNOR2_X1 U599 ( .A(KEYINPUT67), .B(KEYINPUT47), .ZN(n508) );
  NAND2_X1 U600 ( .A1(n593), .A2(n508), .ZN(n509) );
  XNOR2_X1 U601 ( .A(n509), .B(KEYINPUT75), .ZN(n510) );
  NAND2_X1 U602 ( .A1(n349), .A2(n510), .ZN(n511) );
  XNOR2_X2 U603 ( .A(n544), .B(KEYINPUT38), .ZN(n646) );
  INV_X1 U604 ( .A(n646), .ZN(n649) );
  INV_X1 U605 ( .A(n517), .ZN(n518) );
  AND2_X1 U606 ( .A1(n407), .A2(n518), .ZN(n650) );
  NAND2_X1 U607 ( .A1(n650), .A2(n519), .ZN(n520) );
  OR2_X1 U608 ( .A1(n649), .A2(n520), .ZN(n523) );
  INV_X1 U609 ( .A(KEYINPUT115), .ZN(n521) );
  XNOR2_X1 U610 ( .A(n521), .B(KEYINPUT41), .ZN(n522) );
  XNOR2_X2 U611 ( .A(n523), .B(n522), .ZN(n674) );
  NAND2_X1 U612 ( .A1(n674), .A2(n524), .ZN(n526) );
  XNOR2_X1 U613 ( .A(KEYINPUT116), .B(KEYINPUT42), .ZN(n525) );
  XNOR2_X1 U614 ( .A(n526), .B(n525), .ZN(n620) );
  NAND2_X1 U615 ( .A1(n527), .A2(n646), .ZN(n529) );
  XNOR2_X1 U616 ( .A(KEYINPUT72), .B(KEYINPUT39), .ZN(n528) );
  XNOR2_X1 U617 ( .A(n529), .B(n528), .ZN(n551) );
  NAND2_X1 U618 ( .A1(n551), .A2(n617), .ZN(n532) );
  XNOR2_X1 U619 ( .A(KEYINPUT114), .B(KEYINPUT40), .ZN(n531) );
  XNOR2_X1 U620 ( .A(n532), .B(n531), .ZN(n619) );
  NAND2_X1 U621 ( .A1(n620), .A2(n619), .ZN(n535) );
  XNOR2_X1 U622 ( .A(KEYINPUT89), .B(KEYINPUT46), .ZN(n533) );
  XNOR2_X1 U623 ( .A(n533), .B(KEYINPUT64), .ZN(n534) );
  XNOR2_X1 U624 ( .A(n535), .B(n534), .ZN(n536) );
  NAND2_X1 U625 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U626 ( .A(n538), .B(n353), .ZN(n547) );
  AND2_X1 U627 ( .A1(n570), .A2(n498), .ZN(n539) );
  NAND2_X1 U628 ( .A1(n539), .A2(n617), .ZN(n541) );
  OR2_X1 U629 ( .A1(n541), .A2(n540), .ZN(n543) );
  XNOR2_X1 U630 ( .A(KEYINPUT110), .B(KEYINPUT43), .ZN(n542) );
  XNOR2_X1 U631 ( .A(n543), .B(n542), .ZN(n545) );
  AND2_X1 U632 ( .A1(n545), .A2(n544), .ZN(n691) );
  INV_X1 U633 ( .A(n691), .ZN(n546) );
  INV_X1 U634 ( .A(KEYINPUT86), .ZN(n548) );
  INV_X1 U635 ( .A(n550), .ZN(n688) );
  NAND2_X1 U636 ( .A1(n551), .A2(n688), .ZN(n614) );
  XNOR2_X1 U637 ( .A(G898), .B(KEYINPUT97), .ZN(n713) );
  NAND2_X1 U638 ( .A1(G953), .A2(n713), .ZN(n709) );
  NOR2_X1 U639 ( .A1(n709), .A2(n553), .ZN(n554) );
  NOR2_X1 U640 ( .A1(n555), .A2(n554), .ZN(n556) );
  INV_X1 U641 ( .A(n650), .ZN(n561) );
  INV_X1 U642 ( .A(n657), .ZN(n560) );
  XNOR2_X1 U643 ( .A(KEYINPUT65), .B(KEYINPUT22), .ZN(n563) );
  XNOR2_X1 U644 ( .A(n564), .B(n563), .ZN(n576) );
  INV_X1 U645 ( .A(n572), .ZN(n582) );
  NOR2_X1 U646 ( .A1(n485), .A2(n582), .ZN(n565) );
  NAND2_X1 U647 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U648 ( .A(n567), .B(KEYINPUT80), .ZN(n568) );
  NOR2_X1 U649 ( .A1(n576), .A2(n568), .ZN(n569) );
  XOR2_X1 U650 ( .A(KEYINPUT32), .B(n569), .Z(n733) );
  INV_X1 U651 ( .A(n655), .ZN(n571) );
  NAND2_X1 U652 ( .A1(n644), .A2(n592), .ZN(n573) );
  NOR2_X2 U653 ( .A1(n576), .A2(n575), .ZN(n584) );
  NAND2_X1 U654 ( .A1(n581), .A2(n584), .ZN(n577) );
  NOR2_X2 U655 ( .A1(n662), .A2(n577), .ZN(n621) );
  NAND2_X1 U656 ( .A1(n733), .A2(n578), .ZN(n580) );
  NOR2_X1 U657 ( .A1(KEYINPUT44), .A2(KEYINPUT71), .ZN(n579) );
  XNOR2_X1 U658 ( .A(n580), .B(n579), .ZN(n599) );
  NAND2_X1 U659 ( .A1(KEYINPUT44), .A2(KEYINPUT71), .ZN(n597) );
  NOR2_X1 U660 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U661 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U662 ( .A(KEYINPUT109), .B(n585), .ZN(n732) );
  NOR2_X1 U663 ( .A1(n586), .A2(n589), .ZN(n665) );
  NAND2_X1 U664 ( .A1(n592), .A2(n665), .ZN(n587) );
  XNOR2_X1 U665 ( .A(n587), .B(KEYINPUT31), .ZN(n689) );
  NOR2_X1 U666 ( .A1(n655), .A2(n348), .ZN(n590) );
  AND2_X1 U667 ( .A1(n590), .A2(n589), .ZN(n591) );
  AND2_X1 U668 ( .A1(n592), .A2(n591), .ZN(n679) );
  OR2_X1 U669 ( .A1(n689), .A2(n679), .ZN(n594) );
  AND2_X1 U670 ( .A1(n594), .A2(n593), .ZN(n595) );
  NOR2_X1 U671 ( .A1(n732), .A2(n595), .ZN(n596) );
  AND2_X1 U672 ( .A1(n597), .A2(n596), .ZN(n598) );
  NAND2_X1 U673 ( .A1(n599), .A2(n598), .ZN(n600) );
  NAND2_X1 U674 ( .A1(n601), .A2(n715), .ZN(n603) );
  XNOR2_X1 U675 ( .A(n603), .B(n602), .ZN(n643) );
  INV_X1 U676 ( .A(n643), .ZN(n607) );
  INV_X1 U677 ( .A(KEYINPUT83), .ZN(n605) );
  NAND2_X1 U678 ( .A1(n698), .A2(G478), .ZN(n609) );
  XNOR2_X1 U679 ( .A(n609), .B(n608), .ZN(n612) );
  INV_X1 U680 ( .A(G952), .ZN(n610) );
  AND2_X1 U681 ( .A1(n610), .A2(G953), .ZN(n707) );
  NAND2_X1 U682 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U683 ( .A(n613), .B(KEYINPUT125), .ZN(G63) );
  XNOR2_X1 U684 ( .A(n614), .B(G134), .ZN(G36) );
  NAND2_X1 U685 ( .A1(n679), .A2(n617), .ZN(n615) );
  XNOR2_X1 U686 ( .A(n615), .B(G104), .ZN(G6) );
  NAND2_X1 U687 ( .A1(n349), .A2(n617), .ZN(n616) );
  XNOR2_X1 U688 ( .A(n616), .B(G146), .ZN(G48) );
  NAND2_X1 U689 ( .A1(n689), .A2(n617), .ZN(n618) );
  XNOR2_X1 U690 ( .A(n618), .B(G113), .ZN(G15) );
  XNOR2_X1 U691 ( .A(n619), .B(G131), .ZN(G33) );
  XNOR2_X1 U692 ( .A(n620), .B(G137), .ZN(G39) );
  XOR2_X1 U693 ( .A(G110), .B(n621), .Z(G12) );
  XOR2_X1 U694 ( .A(KEYINPUT120), .B(KEYINPUT37), .Z(n623) );
  XOR2_X1 U695 ( .A(n623), .B(G125), .Z(n624) );
  XNOR2_X1 U696 ( .A(n625), .B(n624), .ZN(G27) );
  NAND2_X1 U697 ( .A1(n698), .A2(G472), .ZN(n629) );
  XNOR2_X1 U698 ( .A(KEYINPUT92), .B(KEYINPUT62), .ZN(n627) );
  XNOR2_X1 U699 ( .A(n626), .B(n627), .ZN(n628) );
  XNOR2_X1 U700 ( .A(n629), .B(n628), .ZN(n630) );
  NOR2_X2 U701 ( .A1(n630), .A2(n707), .ZN(n632) );
  XOR2_X1 U702 ( .A(KEYINPUT94), .B(KEYINPUT63), .Z(n631) );
  XNOR2_X1 U703 ( .A(n632), .B(n631), .ZN(G57) );
  NAND2_X1 U704 ( .A1(n698), .A2(G210), .ZN(n636) );
  XOR2_X1 U705 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n634) );
  XNOR2_X1 U706 ( .A(n633), .B(n634), .ZN(n635) );
  XNOR2_X1 U707 ( .A(n636), .B(n635), .ZN(n637) );
  NOR2_X2 U708 ( .A1(n637), .A2(n707), .ZN(n639) );
  XOR2_X1 U709 ( .A(KEYINPUT87), .B(KEYINPUT56), .Z(n638) );
  XNOR2_X1 U710 ( .A(n639), .B(n638), .ZN(G51) );
  NAND2_X1 U711 ( .A1(n640), .A2(n374), .ZN(n641) );
  XNOR2_X1 U712 ( .A(n641), .B(KEYINPUT81), .ZN(n642) );
  NOR2_X1 U713 ( .A1(n643), .A2(n642), .ZN(n678) );
  NOR2_X1 U714 ( .A1(n645), .A2(n648), .ZN(n647) );
  NAND2_X1 U715 ( .A1(n647), .A2(n646), .ZN(n653) );
  NAND2_X1 U716 ( .A1(n649), .A2(n648), .ZN(n651) );
  NAND2_X1 U717 ( .A1(n651), .A2(n650), .ZN(n652) );
  NAND2_X1 U718 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U719 ( .A1(n644), .A2(n654), .ZN(n669) );
  NAND2_X1 U720 ( .A1(n570), .A2(n655), .ZN(n656) );
  XNOR2_X1 U721 ( .A(KEYINPUT50), .B(n656), .ZN(n661) );
  NOR2_X1 U722 ( .A1(n485), .A2(n657), .ZN(n659) );
  XNOR2_X1 U723 ( .A(KEYINPUT122), .B(KEYINPUT49), .ZN(n658) );
  XNOR2_X1 U724 ( .A(n659), .B(n658), .ZN(n660) );
  NAND2_X1 U725 ( .A1(n661), .A2(n660), .ZN(n663) );
  NOR2_X1 U726 ( .A1(n663), .A2(n662), .ZN(n664) );
  NOR2_X1 U727 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U728 ( .A(n666), .B(KEYINPUT51), .ZN(n667) );
  NAND2_X1 U729 ( .A1(n667), .A2(n674), .ZN(n668) );
  NAND2_X1 U730 ( .A1(n669), .A2(n668), .ZN(n671) );
  XOR2_X1 U731 ( .A(KEYINPUT123), .B(KEYINPUT52), .Z(n670) );
  XNOR2_X1 U732 ( .A(n671), .B(n670), .ZN(n673) );
  NAND2_X1 U733 ( .A1(n673), .A2(n672), .ZN(n676) );
  NAND2_X1 U734 ( .A1(n644), .A2(n674), .ZN(n675) );
  NAND2_X1 U735 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U736 ( .A(G107), .B(KEYINPUT27), .ZN(n683) );
  XOR2_X1 U737 ( .A(KEYINPUT118), .B(KEYINPUT26), .Z(n681) );
  NAND2_X1 U738 ( .A1(n679), .A2(n688), .ZN(n680) );
  XNOR2_X1 U739 ( .A(n681), .B(n680), .ZN(n682) );
  XNOR2_X1 U740 ( .A(n683), .B(n682), .ZN(G9) );
  XOR2_X1 U741 ( .A(G128), .B(KEYINPUT29), .Z(n685) );
  NAND2_X1 U742 ( .A1(n349), .A2(n688), .ZN(n684) );
  XNOR2_X1 U743 ( .A(n685), .B(n684), .ZN(G30) );
  XOR2_X1 U744 ( .A(G143), .B(KEYINPUT119), .Z(n686) );
  XNOR2_X1 U745 ( .A(n687), .B(n686), .ZN(G45) );
  NAND2_X1 U746 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U747 ( .A(n690), .B(G116), .ZN(G18) );
  XNOR2_X1 U748 ( .A(n691), .B(G140), .ZN(n692) );
  XNOR2_X1 U749 ( .A(n692), .B(KEYINPUT121), .ZN(G42) );
  NAND2_X1 U750 ( .A1(n698), .A2(G469), .ZN(n696) );
  XOR2_X1 U751 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n693) );
  NOR2_X1 U752 ( .A1(n707), .A2(n697), .ZN(G54) );
  NAND2_X1 U753 ( .A1(n698), .A2(G475), .ZN(n701) );
  XOR2_X1 U754 ( .A(KEYINPUT59), .B(n699), .Z(n700) );
  XNOR2_X1 U755 ( .A(n701), .B(n700), .ZN(n702) );
  NOR2_X2 U756 ( .A1(n702), .A2(n707), .ZN(n703) );
  XNOR2_X1 U757 ( .A(n703), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U758 ( .A1(n698), .A2(G217), .ZN(n705) );
  XNOR2_X1 U759 ( .A(n704), .B(n705), .ZN(n706) );
  NOR2_X1 U760 ( .A1(n707), .A2(n706), .ZN(G66) );
  XOR2_X1 U761 ( .A(n708), .B(G101), .Z(n710) );
  NAND2_X1 U762 ( .A1(n710), .A2(n709), .ZN(n719) );
  XOR2_X1 U763 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n712) );
  NAND2_X1 U764 ( .A1(G224), .A2(G953), .ZN(n711) );
  XNOR2_X1 U765 ( .A(n712), .B(n711), .ZN(n714) );
  NOR2_X1 U766 ( .A1(n714), .A2(n713), .ZN(n717) );
  AND2_X1 U767 ( .A1(n723), .A2(n715), .ZN(n716) );
  NOR2_X1 U768 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U769 ( .A(n719), .B(n718), .ZN(G69) );
  XNOR2_X1 U770 ( .A(n721), .B(n720), .ZN(n725) );
  XOR2_X1 U771 ( .A(n725), .B(n722), .Z(n724) );
  NAND2_X1 U772 ( .A1(n724), .A2(n723), .ZN(n730) );
  XNOR2_X1 U773 ( .A(G227), .B(n725), .ZN(n726) );
  NAND2_X1 U774 ( .A1(n726), .A2(G900), .ZN(n727) );
  NAND2_X1 U775 ( .A1(n727), .A2(G953), .ZN(n728) );
  XOR2_X1 U776 ( .A(KEYINPUT127), .B(n728), .Z(n729) );
  NAND2_X1 U777 ( .A1(n730), .A2(n729), .ZN(G72) );
  XOR2_X1 U778 ( .A(n731), .B(G122), .Z(G24) );
  XOR2_X1 U779 ( .A(G101), .B(n732), .Z(G3) );
  XNOR2_X1 U780 ( .A(G119), .B(n733), .ZN(G21) );
endmodule

