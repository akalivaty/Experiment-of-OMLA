//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 0 1 1 0 0 0 1 0 1 1 0 0 1 1 1 0 1 1 0 1 0 0 1 1 1 1 0 1 1 1 0 0 0 0 1 0 0 1 1 1 1 0 1 0 0 0 0 1 0 1 0 1 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:51 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1253, new_n1254, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT64), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n211));
  NAND3_X1  g0011(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  OAI21_X1  g0012(.A(new_n206), .B1(new_n208), .B2(new_n212), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT1), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n206), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  INV_X1    g0016(.A(KEYINPUT0), .ZN(new_n217));
  INV_X1    g0017(.A(new_n201), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G50), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  INV_X1    g0021(.A(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(new_n216), .A2(new_n217), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n224), .B1(new_n217), .B2(new_n216), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n214), .A2(new_n225), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT2), .B(G226), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(G250), .B(G257), .Z(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n230), .B(new_n233), .ZN(G358));
  XNOR2_X1  g0034(.A(G50), .B(G68), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G58), .B(G77), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n235), .B(new_n236), .Z(new_n237));
  XOR2_X1   g0037(.A(G87), .B(G116), .Z(new_n238));
  XNOR2_X1  g0038(.A(G97), .B(G107), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G351));
  INV_X1    g0041(.A(G1), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(KEYINPUT65), .ZN(new_n243));
  INV_X1    g0043(.A(KEYINPUT65), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(G1), .ZN(new_n245));
  AOI21_X1  g0045(.A(new_n222), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(new_n221), .ZN(new_n248));
  NOR2_X1   g0048(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G50), .ZN(new_n250));
  XNOR2_X1  g0050(.A(KEYINPUT65), .B(G1), .ZN(new_n251));
  INV_X1    g0051(.A(G13), .ZN(new_n252));
  NOR3_X1   g0052(.A1(new_n251), .A2(new_n252), .A3(new_n222), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n202), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n250), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n248), .ZN(new_n257));
  XOR2_X1   g0057(.A(KEYINPUT8), .B(G58), .Z(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(G20), .ZN(new_n260));
  NOR2_X1   g0060(.A1(G20), .A2(G33), .ZN(new_n261));
  AOI22_X1  g0061(.A1(new_n258), .A2(new_n260), .B1(G150), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n203), .A2(G20), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n257), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  OR2_X1    g0065(.A1(KEYINPUT70), .A2(KEYINPUT9), .ZN(new_n266));
  NAND2_X1  g0066(.A1(KEYINPUT70), .A2(KEYINPUT9), .ZN(new_n267));
  NAND4_X1  g0067(.A1(new_n256), .A2(new_n265), .A3(new_n266), .A4(new_n267), .ZN(new_n268));
  OAI211_X1 g0068(.A(KEYINPUT70), .B(KEYINPUT9), .C1(new_n255), .C2(new_n264), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(G41), .A2(G45), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n272), .A2(new_n242), .A3(G274), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  XNOR2_X1  g0074(.A(KEYINPUT3), .B(G33), .ZN(new_n275));
  INV_X1    g0075(.A(G1698), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n275), .A2(G222), .A3(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G77), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n275), .A2(G1698), .ZN(new_n279));
  INV_X1    g0079(.A(G223), .ZN(new_n280));
  OAI221_X1 g0080(.A(new_n277), .B1(new_n278), .B2(new_n275), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(G33), .A2(G41), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n282), .A2(G1), .A3(G13), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n274), .B1(new_n281), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT66), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n286), .B1(new_n251), .B2(new_n271), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n244), .A2(G1), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n242), .A2(KEYINPUT65), .ZN(new_n289));
  OAI211_X1 g0089(.A(KEYINPUT66), .B(new_n272), .C1(new_n288), .C2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n284), .B1(new_n287), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G226), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n285), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G200), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n285), .A2(G190), .A3(new_n292), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n270), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  XNOR2_X1  g0096(.A(new_n296), .B(KEYINPUT10), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT71), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n275), .A2(G226), .A3(new_n276), .ZN(new_n299));
  NAND2_X1  g0099(.A1(G33), .A2(G97), .ZN(new_n300));
  INV_X1    g0100(.A(G232), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n299), .B(new_n300), .C1(new_n279), .C2(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n274), .B1(new_n302), .B2(new_n284), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT13), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n291), .A2(G238), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n304), .B1(new_n303), .B2(new_n305), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G200), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n298), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G68), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n253), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g0113(.A(new_n313), .B(KEYINPUT12), .ZN(new_n314));
  AOI22_X1  g0114(.A1(new_n260), .A2(G77), .B1(G20), .B2(new_n312), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n261), .A2(G50), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n257), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  OR2_X1    g0117(.A1(new_n317), .A2(KEYINPUT11), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n249), .A2(G68), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n317), .A2(KEYINPUT11), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n314), .A2(new_n318), .A3(new_n319), .A4(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n321), .B1(new_n309), .B2(G190), .ZN(new_n322));
  OAI211_X1 g0122(.A(KEYINPUT71), .B(G200), .C1(new_n307), .C2(new_n308), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n311), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n255), .A2(new_n264), .ZN(new_n325));
  INV_X1    g0125(.A(G169), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n325), .B1(new_n293), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G179), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n285), .A2(new_n328), .A3(new_n292), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n253), .A2(new_n278), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT68), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n331), .A2(new_n332), .B1(G77), .B2(new_n249), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n253), .A2(KEYINPUT68), .A3(new_n278), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(KEYINPUT15), .A2(G87), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT67), .ZN(new_n338));
  NAND2_X1  g0138(.A1(KEYINPUT15), .A2(G87), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n339), .ZN(new_n341));
  OAI21_X1  g0141(.A(KEYINPUT67), .B1(new_n341), .B2(new_n336), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n260), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n258), .A2(new_n261), .B1(G20), .B2(G77), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n257), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  OR2_X1    g0147(.A1(new_n335), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT69), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n275), .A2(G238), .A3(G1698), .ZN(new_n350));
  INV_X1    g0150(.A(G107), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n275), .A2(new_n276), .ZN(new_n352));
  OAI221_X1 g0152(.A(new_n350), .B1(new_n351), .B2(new_n275), .C1(new_n352), .C2(new_n301), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n274), .B1(new_n353), .B2(new_n284), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n291), .A2(G244), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n348), .A2(new_n349), .B1(G200), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n356), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n335), .A2(new_n347), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n358), .A2(G190), .B1(new_n359), .B2(KEYINPUT69), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n297), .A2(new_n324), .A3(new_n330), .A4(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n308), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n363), .A2(G179), .A3(new_n306), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n326), .B1(new_n363), .B2(new_n306), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT14), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(G169), .B1(new_n307), .B2(new_n308), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n368), .A2(KEYINPUT14), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n321), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n358), .A2(new_n328), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n356), .A2(new_n326), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n371), .A2(new_n348), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT72), .ZN(new_n375));
  AOI211_X1 g0175(.A(new_n301), .B(new_n284), .C1(new_n287), .C2(new_n290), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n375), .B1(new_n376), .B2(new_n274), .ZN(new_n377));
  NOR3_X1   g0177(.A1(new_n251), .A2(new_n286), .A3(new_n271), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n243), .A2(new_n245), .ZN(new_n379));
  AOI21_X1  g0179(.A(KEYINPUT66), .B1(new_n379), .B2(new_n272), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n283), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  OAI211_X1 g0181(.A(KEYINPUT72), .B(new_n273), .C1(new_n381), .C2(new_n301), .ZN(new_n382));
  INV_X1    g0182(.A(G190), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n275), .A2(G226), .A3(G1698), .ZN(new_n384));
  INV_X1    g0184(.A(G87), .ZN(new_n385));
  OAI221_X1 g0185(.A(new_n384), .B1(new_n259), .B2(new_n385), .C1(new_n352), .C2(new_n280), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(new_n284), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n377), .A2(new_n382), .A3(new_n383), .A4(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n274), .B1(new_n291), .B2(G232), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n387), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(new_n310), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT17), .ZN(new_n393));
  OAI211_X1 g0193(.A(G13), .B(G20), .C1(new_n288), .C2(new_n289), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n394), .A2(new_n258), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n395), .B1(new_n249), .B2(new_n258), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT3), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(G33), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(KEYINPUT7), .B1(new_n401), .B2(new_n222), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT7), .ZN(new_n403));
  AOI211_X1 g0203(.A(new_n403), .B(G20), .C1(new_n398), .C2(new_n400), .ZN(new_n404));
  OAI21_X1  g0204(.A(G68), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(G58), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n406), .A2(new_n312), .ZN(new_n407));
  OAI21_X1  g0207(.A(G20), .B1(new_n407), .B2(new_n201), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n261), .A2(G159), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n405), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT16), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n257), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n405), .A2(KEYINPUT16), .A3(new_n411), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n397), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  AND3_X1   g0216(.A1(new_n392), .A2(new_n393), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n393), .B1(new_n392), .B2(new_n416), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n403), .B1(new_n275), .B2(G20), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n401), .A2(KEYINPUT7), .A3(new_n222), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n312), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n413), .B1(new_n421), .B2(new_n410), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n415), .A2(new_n422), .A3(new_n248), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n396), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n377), .A2(new_n382), .A3(new_n328), .A4(new_n387), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n390), .A2(new_n326), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT18), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n423), .A2(new_n396), .B1(new_n390), .B2(new_n326), .ZN(new_n430));
  AOI21_X1  g0230(.A(KEYINPUT18), .B1(new_n430), .B2(new_n425), .ZN(new_n431));
  OAI22_X1  g0231(.A1(new_n417), .A2(new_n418), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  NOR3_X1   g0232(.A1(new_n362), .A2(new_n374), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n379), .A2(G33), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n394), .A2(new_n434), .A3(G116), .A4(new_n257), .ZN(new_n435));
  INV_X1    g0235(.A(G116), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n253), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n247), .A2(new_n221), .B1(G20), .B2(new_n436), .ZN(new_n439));
  NAND2_X1  g0239(.A1(G33), .A2(G283), .ZN(new_n440));
  INV_X1    g0240(.A(G97), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n440), .B(new_n222), .C1(G33), .C2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n439), .A2(KEYINPUT20), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(KEYINPUT20), .B1(new_n439), .B2(new_n442), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(KEYINPUT77), .B1(new_n438), .B2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n445), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(new_n443), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT77), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n449), .A2(new_n450), .A3(new_n435), .A4(new_n437), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n447), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n398), .A2(new_n400), .A3(G257), .A4(new_n276), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n398), .A2(new_n400), .A3(G264), .A4(G1698), .ZN(new_n454));
  INV_X1    g0254(.A(G303), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n453), .B(new_n454), .C1(new_n455), .C2(new_n275), .ZN(new_n456));
  AND2_X1   g0256(.A1(new_n456), .A2(new_n284), .ZN(new_n457));
  XNOR2_X1  g0257(.A(KEYINPUT5), .B(G41), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n379), .A2(new_n458), .A3(G45), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n459), .A2(G270), .A3(new_n283), .ZN(new_n460));
  INV_X1    g0260(.A(G45), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n461), .B1(new_n243), .B2(new_n245), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n462), .A2(G274), .A3(new_n283), .A4(new_n458), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(G169), .B1(new_n457), .B2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n452), .A2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT21), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n467), .A2(KEYINPUT78), .A3(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n464), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n456), .A2(new_n284), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n472), .A2(new_n383), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n310), .B1(new_n470), .B2(new_n471), .ZN(new_n474));
  OR3_X1    g0274(.A1(new_n473), .A2(new_n452), .A3(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n472), .A2(new_n328), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n452), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n465), .B1(new_n451), .B2(new_n447), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT78), .ZN(new_n479));
  OAI21_X1  g0279(.A(KEYINPUT21), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AND4_X1   g0280(.A1(new_n469), .A2(new_n475), .A3(new_n477), .A4(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT76), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n394), .A2(new_n434), .A3(new_n257), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(G87), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT75), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n222), .A2(G33), .A3(G97), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT19), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT74), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n222), .B1(new_n300), .B2(new_n488), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n385), .A2(new_n441), .A3(new_n351), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n398), .A2(new_n400), .A3(new_n222), .A4(G68), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT74), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n487), .A2(new_n495), .A3(new_n488), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n490), .A2(new_n493), .A3(new_n494), .A4(new_n496), .ZN(new_n497));
  AOI221_X4 g0297(.A(new_n486), .B1(new_n343), .B2(new_n253), .C1(new_n497), .C2(new_n248), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n248), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n343), .A2(new_n253), .ZN(new_n500));
  AOI21_X1  g0300(.A(KEYINPUT75), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n485), .B1(new_n498), .B2(new_n501), .ZN(new_n502));
  OAI211_X1 g0302(.A(G250), .B(new_n283), .C1(new_n251), .C2(new_n461), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n379), .A2(new_n283), .A3(G45), .A4(G274), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n398), .A2(new_n400), .A3(G244), .A4(G1698), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n398), .A2(new_n400), .A3(G238), .A4(new_n276), .ZN(new_n507));
  NAND2_X1  g0307(.A1(G33), .A2(G116), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n505), .B1(new_n284), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(G190), .ZN(new_n511));
  AND2_X1   g0311(.A1(new_n503), .A2(new_n504), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n509), .A2(new_n284), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(G200), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n502), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n512), .A2(new_n328), .A3(new_n513), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(new_n510), .B2(G169), .ZN(new_n519));
  AND2_X1   g0319(.A1(new_n493), .A2(new_n494), .ZN(new_n520));
  AND3_X1   g0320(.A1(new_n487), .A2(new_n495), .A3(new_n488), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n495), .B1(new_n487), .B2(new_n488), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n257), .B1(new_n520), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n500), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n486), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n499), .A2(KEYINPUT75), .A3(new_n500), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n484), .A2(new_n344), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n519), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n482), .B1(new_n517), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n529), .B1(new_n498), .B2(new_n501), .ZN(new_n532));
  INV_X1    g0332(.A(new_n519), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n528), .A2(new_n485), .A3(new_n515), .A4(new_n511), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n534), .A2(new_n535), .A3(KEYINPUT76), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n531), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n398), .A2(new_n400), .A3(G244), .A4(new_n276), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT4), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n275), .A2(KEYINPUT4), .A3(G244), .A4(new_n276), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n275), .A2(G250), .A3(G1698), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n540), .A2(new_n541), .A3(new_n440), .A4(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n284), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n284), .B1(new_n462), .B2(new_n458), .ZN(new_n545));
  AND2_X1   g0345(.A1(G33), .A2(G41), .ZN(new_n546));
  OAI21_X1  g0346(.A(G274), .B1(new_n546), .B2(new_n221), .ZN(new_n547));
  NOR3_X1   g0347(.A1(new_n547), .A2(new_n251), .A3(new_n461), .ZN(new_n548));
  AOI22_X1  g0348(.A1(G257), .A2(new_n545), .B1(new_n548), .B2(new_n458), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n544), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n326), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n544), .A2(new_n549), .A3(new_n328), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n261), .A2(G77), .ZN(new_n553));
  AND3_X1   g0353(.A1(new_n351), .A2(KEYINPUT6), .A3(G97), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT6), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n554), .B1(new_n239), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n553), .B1(new_n556), .B2(new_n222), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT73), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n419), .A2(new_n420), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n557), .A2(new_n558), .B1(new_n559), .B2(G107), .ZN(new_n560));
  OAI211_X1 g0360(.A(KEYINPUT73), .B(new_n553), .C1(new_n556), .C2(new_n222), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n257), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n394), .A2(G97), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n564), .B1(new_n483), .B2(new_n441), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n551), .B(new_n552), .C1(new_n562), .C2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n351), .A2(G97), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n441), .A2(G107), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n567), .A2(new_n568), .A3(new_n555), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n351), .A2(KEYINPUT6), .A3(G97), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n222), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n553), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n558), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  OAI21_X1  g0373(.A(G107), .B1(new_n402), .B2(new_n404), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n573), .A2(new_n561), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n565), .B1(new_n575), .B2(new_n248), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n550), .A2(G200), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n544), .A2(new_n549), .A3(G190), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n566), .A2(new_n579), .ZN(new_n580));
  OAI21_X1  g0380(.A(KEYINPUT80), .B1(new_n394), .B2(G107), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT80), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n246), .A2(new_n582), .A3(G13), .A4(new_n351), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n581), .A2(KEYINPUT25), .A3(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n394), .A2(new_n434), .A3(G107), .A4(new_n257), .ZN(new_n585));
  AND2_X1   g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n581), .A2(new_n583), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT25), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n260), .A2(G116), .ZN(new_n590));
  OR3_X1    g0390(.A1(new_n222), .A2(KEYINPUT23), .A3(G107), .ZN(new_n591));
  OAI21_X1  g0391(.A(KEYINPUT23), .B1(new_n222), .B2(G107), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n385), .B1(KEYINPUT79), .B2(KEYINPUT22), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n275), .A2(new_n222), .A3(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(KEYINPUT79), .A2(KEYINPUT22), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n275), .A2(new_n594), .A3(new_n222), .A4(new_n596), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n593), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  AND2_X1   g0400(.A1(new_n600), .A2(KEYINPUT24), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n248), .B1(new_n600), .B2(KEYINPUT24), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n586), .B(new_n589), .C1(new_n601), .C2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n275), .A2(G250), .A3(new_n276), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n275), .A2(G257), .A3(G1698), .ZN(new_n605));
  NAND2_X1  g0405(.A1(G33), .A2(G294), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  AND2_X1   g0407(.A1(new_n607), .A2(new_n284), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n545), .A2(G264), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n463), .ZN(new_n610));
  OAI21_X1  g0410(.A(G169), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n607), .A2(new_n284), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT81), .ZN(new_n613));
  AND3_X1   g0413(.A1(new_n545), .A2(new_n613), .A3(G264), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n613), .B1(new_n545), .B2(G264), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n463), .B(new_n612), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n611), .B1(new_n616), .B2(new_n328), .ZN(new_n617));
  AND2_X1   g0417(.A1(new_n603), .A2(new_n617), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n612), .A2(new_n463), .A3(new_n609), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n616), .A2(new_n310), .B1(new_n619), .B2(new_n383), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n620), .A2(new_n603), .ZN(new_n621));
  NOR3_X1   g0421(.A1(new_n580), .A2(new_n618), .A3(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n433), .A2(new_n481), .A3(new_n537), .A4(new_n622), .ZN(new_n623));
  XOR2_X1   g0423(.A(new_n623), .B(KEYINPUT82), .Z(G372));
  NAND2_X1  g0424(.A1(new_n427), .A2(new_n428), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n430), .A2(KEYINPUT18), .A3(new_n425), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n392), .A2(new_n416), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(KEYINPUT17), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n424), .B1(new_n391), .B2(new_n388), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n393), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n633), .A2(new_n324), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n628), .B1(new_n634), .B2(new_n374), .ZN(new_n635));
  INV_X1    g0435(.A(new_n297), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n330), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n566), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n531), .A2(new_n536), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(KEYINPUT26), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n603), .A2(new_n617), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n480), .A2(new_n469), .A3(new_n477), .A4(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n580), .A2(new_n621), .ZN(new_n643));
  AOI21_X1  g0443(.A(KEYINPUT83), .B1(new_n534), .B2(new_n535), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n534), .A2(new_n535), .A3(KEYINPUT83), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n642), .B(new_n643), .C1(new_n644), .C2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT84), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n459), .A2(G257), .A3(new_n283), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(new_n463), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n649), .B1(new_n284), .B2(new_n543), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n552), .B1(new_n650), .B2(G169), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n647), .B1(new_n651), .B2(new_n576), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n575), .A2(new_n248), .ZN(new_n653));
  INV_X1    g0453(.A(new_n565), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n655), .A2(KEYINPUT84), .A3(new_n551), .A4(new_n552), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT26), .ZN(new_n658));
  OAI211_X1 g0458(.A(new_n657), .B(new_n658), .C1(new_n645), .C2(new_n644), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n640), .A2(new_n646), .A3(new_n534), .A4(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n637), .B1(new_n433), .B2(new_n660), .ZN(new_n661));
  XOR2_X1   g0461(.A(new_n661), .B(KEYINPUT85), .Z(G369));
  NAND2_X1  g0462(.A1(new_n222), .A2(G13), .ZN(new_n663));
  OR3_X1    g0463(.A1(new_n251), .A2(KEYINPUT27), .A3(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(KEYINPUT27), .B1(new_n251), .B2(new_n663), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(new_n665), .A3(G213), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(G343), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n452), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n481), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n479), .B1(new_n452), .B2(new_n466), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n477), .B1(new_n672), .B2(new_n468), .ZN(new_n673));
  NOR3_X1   g0473(.A1(new_n478), .A2(new_n479), .A3(KEYINPUT21), .ZN(new_n674));
  OAI211_X1 g0474(.A(new_n452), .B(new_n669), .C1(new_n673), .C2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(KEYINPUT86), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT86), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n671), .A2(new_n678), .A3(new_n675), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n618), .A2(KEYINPUT87), .A3(new_n669), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT87), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n682), .B1(new_n641), .B2(new_n668), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n603), .A2(new_n669), .ZN(new_n685));
  OAI211_X1 g0485(.A(new_n641), .B(new_n685), .C1(new_n603), .C2(new_n620), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n680), .A2(G330), .A3(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n641), .A2(new_n669), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n668), .B1(new_n673), .B2(new_n674), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n689), .B1(new_n687), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n688), .A2(new_n692), .ZN(G399));
  INV_X1    g0493(.A(new_n215), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(G41), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n492), .A2(G116), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n696), .A2(G1), .A3(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(new_n219), .B2(new_n696), .ZN(new_n699));
  XNOR2_X1  g0499(.A(new_n699), .B(KEYINPUT28), .ZN(new_n700));
  INV_X1    g0500(.A(G330), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n612), .B1(new_n614), .B2(new_n615), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(new_n514), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n703), .A2(new_n476), .A3(new_n650), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT30), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n510), .A2(G179), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n707), .A2(new_n616), .A3(new_n472), .A4(new_n550), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n476), .A2(new_n703), .A3(KEYINPUT30), .A4(new_n650), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n706), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT31), .ZN(new_n711));
  AND3_X1   g0511(.A1(new_n710), .A2(new_n711), .A3(new_n669), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n537), .A2(new_n481), .A3(new_n622), .A4(new_n668), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n711), .B1(new_n710), .B2(new_n669), .ZN(new_n714));
  AOI211_X1 g0514(.A(new_n701), .B(new_n712), .C1(new_n713), .C2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n646), .A2(new_n534), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n531), .A2(new_n638), .A3(new_n536), .A4(new_n658), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n652), .A2(new_n656), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT83), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n720), .B1(new_n517), .B2(new_n530), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n534), .A2(new_n535), .A3(KEYINPUT83), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n719), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n718), .B1(new_n723), .B2(new_n658), .ZN(new_n724));
  OAI211_X1 g0524(.A(KEYINPUT29), .B(new_n668), .C1(new_n717), .C2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(KEYINPUT29), .B1(new_n660), .B2(new_n668), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n716), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n700), .B1(new_n729), .B2(G1), .ZN(G364));
  NAND3_X1  g0530(.A1(new_n677), .A2(new_n701), .A3(new_n679), .ZN(new_n731));
  INV_X1    g0531(.A(new_n679), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n678), .B1(new_n671), .B2(new_n675), .ZN(new_n733));
  OAI21_X1  g0533(.A(G330), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n663), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n242), .B1(new_n735), .B2(G45), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(new_n695), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n731), .A2(new_n734), .A3(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n221), .B1(G20), .B2(new_n326), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n222), .A2(new_n383), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n310), .A2(G179), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n222), .A2(G190), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(new_n744), .ZN(new_n747));
  INV_X1    g0547(.A(G283), .ZN(new_n748));
  OAI22_X1  g0548(.A1(new_n745), .A2(new_n455), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n328), .A2(G200), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n746), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  AOI211_X1 g0552(.A(new_n275), .B(new_n749), .C1(G311), .C2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n328), .A2(new_n310), .ZN(new_n754));
  AND2_X1   g0554(.A1(new_n743), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(G326), .ZN(new_n757));
  NOR2_X1   g0557(.A1(G179), .A2(G200), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n222), .B1(new_n758), .B2(G190), .ZN(new_n759));
  INV_X1    g0559(.A(G294), .ZN(new_n760));
  OAI22_X1  g0560(.A1(new_n756), .A2(new_n757), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OR2_X1    g0561(.A1(new_n761), .A2(KEYINPUT91), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(KEYINPUT91), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n743), .A2(new_n750), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n746), .A2(new_n758), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI22_X1  g0567(.A1(G322), .A2(new_n765), .B1(new_n767), .B2(G329), .ZN(new_n768));
  AND2_X1   g0568(.A1(new_n754), .A2(new_n746), .ZN(new_n769));
  XNOR2_X1  g0569(.A(KEYINPUT33), .B(G317), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AND2_X1   g0571(.A1(new_n768), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g0572(.A1(new_n753), .A2(new_n762), .A3(new_n763), .A4(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n769), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n774), .A2(new_n312), .B1(new_n751), .B2(new_n278), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n775), .B1(G58), .B2(new_n765), .ZN(new_n776));
  INV_X1    g0576(.A(new_n745), .ZN(new_n777));
  AOI22_X1  g0577(.A1(new_n777), .A2(G87), .B1(new_n755), .B2(G50), .ZN(new_n778));
  INV_X1    g0578(.A(new_n747), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G107), .ZN(new_n780));
  AND3_X1   g0580(.A1(new_n778), .A2(new_n275), .A3(new_n780), .ZN(new_n781));
  XNOR2_X1  g0581(.A(KEYINPUT90), .B(KEYINPUT32), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n767), .A2(G159), .A3(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n782), .B1(new_n767), .B2(G159), .ZN(new_n784));
  INV_X1    g0584(.A(new_n759), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n784), .B1(G97), .B2(new_n785), .ZN(new_n786));
  NAND4_X1  g0586(.A1(new_n776), .A2(new_n781), .A3(new_n783), .A4(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n742), .B1(new_n773), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(G13), .A2(G33), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(G20), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT89), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n741), .ZN(new_n794));
  OR2_X1    g0594(.A1(new_n237), .A2(new_n461), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n694), .A2(new_n275), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n797), .B1(new_n461), .B2(new_n220), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n694), .A2(new_n401), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n799), .A2(G355), .B1(new_n436), .B2(new_n694), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n795), .A2(new_n798), .B1(KEYINPUT88), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(KEYINPUT88), .B2(new_n801), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n739), .B(new_n788), .C1(new_n794), .C2(new_n803), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n804), .B1(new_n676), .B2(new_n792), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n740), .A2(new_n805), .ZN(G396));
  OAI22_X1  g0606(.A1(new_n774), .A2(new_n748), .B1(new_n760), .B2(new_n764), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n275), .B(new_n807), .C1(G116), .C2(new_n752), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n785), .A2(G97), .ZN(new_n809));
  AOI22_X1  g0609(.A1(G87), .A2(new_n779), .B1(new_n767), .B2(G311), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n777), .A2(G107), .B1(new_n755), .B2(G303), .ZN(new_n811));
  NAND4_X1  g0611(.A1(new_n808), .A2(new_n809), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  AOI22_X1  g0612(.A1(G137), .A2(new_n755), .B1(new_n769), .B2(G150), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT92), .ZN(new_n814));
  AOI22_X1  g0614(.A1(G143), .A2(new_n765), .B1(new_n752), .B2(G159), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n816), .B(KEYINPUT93), .Z(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(KEYINPUT34), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n401), .B1(new_n767), .B2(G132), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT94), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n779), .A2(G68), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n822), .B1(new_n202), .B2(new_n745), .C1(new_n406), .C2(new_n759), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n819), .A2(new_n820), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n818), .A2(new_n821), .A3(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n817), .A2(KEYINPUT34), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n812), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  AND2_X1   g0628(.A1(new_n828), .A2(KEYINPUT95), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n828), .A2(KEYINPUT95), .ZN(new_n830));
  NOR3_X1   g0630(.A1(new_n829), .A2(new_n830), .A3(new_n742), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n741), .A2(new_n789), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n373), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n834), .A2(new_n668), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n357), .A2(new_n360), .B1(new_n348), .B2(new_n669), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n835), .B1(new_n836), .B2(new_n834), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n738), .B1(G77), .B2(new_n833), .C1(new_n838), .C2(new_n790), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n831), .A2(new_n839), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n660), .A2(new_n668), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n841), .B(new_n838), .ZN(new_n842));
  OR2_X1    g0642(.A1(new_n842), .A2(new_n716), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n738), .B1(new_n842), .B2(new_n716), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n840), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(G384));
  OAI21_X1  g0646(.A(G77), .B1(new_n406), .B2(new_n312), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n219), .A2(new_n847), .B1(G50), .B2(new_n312), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n848), .A2(new_n252), .A3(new_n251), .ZN(new_n849));
  INV_X1    g0649(.A(new_n556), .ZN(new_n850));
  OAI211_X1 g0650(.A(G116), .B(new_n223), .C1(new_n850), .C2(KEYINPUT35), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n851), .B1(KEYINPUT35), .B2(new_n850), .ZN(new_n852));
  XOR2_X1   g0652(.A(new_n852), .B(KEYINPUT96), .Z(new_n853));
  INV_X1    g0653(.A(KEYINPUT36), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n849), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(new_n854), .B2(new_n853), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT38), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n666), .B1(new_n423), .B2(new_n396), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n859), .B1(new_n633), .B2(new_n627), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n629), .A2(new_n427), .A3(new_n859), .ZN(new_n861));
  OAI21_X1  g0661(.A(KEYINPUT37), .B1(new_n858), .B2(KEYINPUT97), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n858), .B1(new_n430), .B2(new_n425), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT97), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(new_n416), .B2(new_n666), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n864), .A2(KEYINPUT37), .A3(new_n629), .A4(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n863), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n857), .B1(new_n860), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n432), .A2(new_n858), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n427), .A2(new_n859), .ZN(new_n871));
  NOR3_X1   g0671(.A1(new_n871), .A2(new_n862), .A3(new_n631), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n864), .A2(new_n629), .B1(new_n866), .B2(KEYINPUT37), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n870), .A2(new_n874), .A3(KEYINPUT38), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n869), .A2(new_n875), .A3(KEYINPUT98), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n712), .B1(new_n713), .B2(new_n714), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT98), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n878), .B(new_n857), .C1(new_n860), .C2(new_n868), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n321), .A2(new_n669), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n365), .A2(new_n366), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n368), .A2(KEYINPUT14), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n881), .A2(new_n882), .A3(new_n364), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n324), .A2(new_n880), .B1(new_n883), .B2(new_n321), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n370), .A2(new_n669), .ZN(new_n885));
  NOR3_X1   g0685(.A1(new_n884), .A2(new_n885), .A3(new_n837), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n876), .A2(new_n877), .A3(new_n879), .A4(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT40), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AND2_X1   g0689(.A1(new_n886), .A2(new_n877), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT37), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n861), .B(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n857), .B1(new_n892), .B2(new_n860), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n888), .B1(new_n893), .B2(new_n875), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n890), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n889), .A2(new_n895), .A3(G330), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n877), .A2(new_n433), .A3(G330), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AOI22_X1  g0698(.A1(new_n887), .A2(new_n888), .B1(new_n890), .B2(new_n894), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n899), .A2(new_n433), .A3(new_n877), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n433), .B(new_n725), .C1(new_n841), .C2(KEYINPUT29), .ZN(new_n902));
  INV_X1    g0702(.A(new_n637), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  XOR2_X1   g0704(.A(new_n901), .B(new_n904), .Z(new_n905));
  NAND3_X1  g0705(.A1(new_n876), .A2(KEYINPUT39), .A3(new_n879), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT39), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n893), .A2(new_n907), .A3(new_n875), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n885), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n628), .A2(new_n666), .ZN(new_n911));
  AND2_X1   g0711(.A1(new_n876), .A2(new_n879), .ZN(new_n912));
  INV_X1    g0712(.A(new_n884), .ZN(new_n913));
  INV_X1    g0713(.A(new_n885), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n660), .A2(new_n668), .A3(new_n838), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n915), .B1(new_n916), .B2(new_n835), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n912), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n910), .A2(new_n911), .A3(new_n918), .ZN(new_n919));
  OAI22_X1  g0719(.A1(new_n905), .A2(new_n919), .B1(new_n379), .B2(new_n735), .ZN(new_n920));
  AND2_X1   g0720(.A1(new_n905), .A2(new_n919), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n856), .B1(new_n920), .B2(new_n921), .ZN(G367));
  OAI221_X1 g0722(.A(new_n794), .B1(new_n215), .B2(new_n343), .C1(new_n233), .C2(new_n797), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n739), .B1(new_n923), .B2(KEYINPUT104), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(KEYINPUT104), .B2(new_n923), .ZN(new_n925));
  OAI22_X1  g0725(.A1(new_n441), .A2(new_n747), .B1(new_n751), .B2(new_n748), .ZN(new_n926));
  AOI211_X1 g0726(.A(new_n275), .B(new_n926), .C1(G303), .C2(new_n765), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n755), .A2(G311), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n774), .B2(new_n760), .ZN(new_n929));
  XOR2_X1   g0729(.A(KEYINPUT105), .B(G317), .Z(new_n930));
  AOI21_X1  g0730(.A(new_n929), .B1(new_n767), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n777), .A2(KEYINPUT46), .A3(G116), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT46), .B1(new_n777), .B2(G116), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n933), .B1(G107), .B2(new_n785), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n927), .A2(new_n931), .A3(new_n932), .A4(new_n934), .ZN(new_n935));
  OAI22_X1  g0735(.A1(new_n745), .A2(new_n406), .B1(new_n751), .B2(new_n202), .ZN(new_n936));
  AOI211_X1 g0736(.A(new_n401), .B(new_n936), .C1(G159), .C2(new_n769), .ZN(new_n937));
  XNOR2_X1  g0737(.A(KEYINPUT106), .B(G137), .ZN(new_n938));
  AOI22_X1  g0738(.A1(G150), .A2(new_n765), .B1(new_n767), .B2(new_n938), .ZN(new_n939));
  AOI22_X1  g0739(.A1(G77), .A2(new_n779), .B1(new_n755), .B2(G143), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n785), .A2(G68), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n937), .A2(new_n939), .A3(new_n940), .A4(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n935), .A2(new_n942), .A3(KEYINPUT47), .ZN(new_n943));
  AOI21_X1  g0743(.A(KEYINPUT47), .B1(new_n935), .B2(new_n942), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n944), .A2(new_n742), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n925), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n502), .A2(new_n669), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n645), .B2(new_n644), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n530), .A2(new_n502), .A3(new_n669), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n946), .B1(new_n950), .B2(new_n792), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n687), .A2(new_n691), .ZN(new_n952));
  INV_X1    g0752(.A(new_n689), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n566), .B(new_n579), .C1(new_n576), .C2(new_n668), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT99), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n955), .B(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n638), .A2(new_n669), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(KEYINPUT44), .B1(new_n954), .B2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT44), .ZN(new_n962));
  NOR3_X1   g0762(.A1(new_n692), .A2(new_n959), .A3(new_n962), .ZN(new_n963));
  AND3_X1   g0763(.A1(new_n692), .A2(KEYINPUT45), .A3(new_n959), .ZN(new_n964));
  AOI21_X1  g0764(.A(KEYINPUT45), .B1(new_n692), .B2(new_n959), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n961), .A2(new_n963), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n688), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n965), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n692), .A2(KEYINPUT45), .A3(new_n959), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n954), .A2(new_n960), .A3(KEYINPUT44), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n962), .B1(new_n692), .B2(new_n959), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n971), .A2(new_n688), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n968), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n687), .A2(new_n691), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n690), .B1(new_n684), .B2(new_n686), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n734), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n680), .A2(new_n979), .A3(G330), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n729), .B1(new_n976), .B2(new_n983), .ZN(new_n984));
  XNOR2_X1  g0784(.A(KEYINPUT103), .B(KEYINPUT41), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n695), .B(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n737), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT42), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n692), .B2(new_n957), .ZN(new_n989));
  INV_X1    g0789(.A(new_n957), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n990), .A2(KEYINPUT42), .A3(new_n978), .A4(new_n641), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n989), .A2(new_n991), .B1(new_n638), .B2(new_n668), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT101), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT43), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n948), .A2(new_n995), .A3(new_n949), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n950), .A2(KEYINPUT43), .ZN(new_n998));
  AND2_X1   g0798(.A1(new_n998), .A2(KEYINPUT100), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n998), .A2(KEYINPUT100), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n993), .A2(new_n994), .A3(new_n997), .A4(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n997), .A2(new_n994), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n996), .A2(KEYINPUT101), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1001), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n1003), .B(new_n1004), .C1(new_n1005), .C2(new_n992), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1002), .A2(new_n1006), .ZN(new_n1007));
  OR3_X1    g0807(.A1(new_n688), .A2(KEYINPUT102), .A3(new_n960), .ZN(new_n1008));
  OAI21_X1  g0808(.A(KEYINPUT102), .B1(new_n688), .B2(new_n960), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n1002), .A2(new_n1006), .A3(new_n1008), .A4(new_n1009), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n951), .B1(new_n987), .B2(new_n1013), .ZN(G387));
  NOR2_X1   g0814(.A1(new_n734), .A2(new_n980), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n979), .B1(new_n680), .B2(G330), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n729), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n983), .A2(new_n728), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1018), .A2(new_n695), .A3(new_n1019), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n684), .A2(new_n686), .A3(new_n793), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n765), .A2(new_n930), .B1(new_n752), .B2(G303), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(G322), .A2(new_n755), .B1(new_n769), .B2(G311), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT48), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n745), .A2(new_n760), .B1(new_n759), .B2(new_n748), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT109), .Z(new_n1027));
  AND2_X1   g0827(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  AND2_X1   g0828(.A1(new_n1028), .A2(KEYINPUT49), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n1028), .A2(KEYINPUT49), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n401), .B1(new_n766), .B2(new_n757), .C1(new_n436), .C2(new_n747), .ZN(new_n1031));
  OR3_X1    g0831(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n764), .A2(new_n202), .B1(new_n751), .B2(new_n312), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n401), .B(new_n1033), .C1(G97), .C2(new_n779), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n344), .A2(new_n785), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(KEYINPUT108), .B(G150), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(G159), .A2(new_n755), .B1(new_n767), .B2(new_n1036), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(G77), .A2(new_n777), .B1(new_n769), .B2(new_n258), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n1034), .A2(new_n1035), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n742), .B1(new_n1032), .B2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n230), .A2(new_n461), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n258), .A2(new_n202), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT50), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n697), .B(new_n461), .C1(new_n312), .C2(new_n278), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n796), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1041), .B1(KEYINPUT107), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(KEYINPUT107), .B2(new_n1045), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n799), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1047), .B1(G107), .B2(new_n215), .C1(new_n697), .C2(new_n1048), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n739), .B(new_n1040), .C1(new_n794), .C2(new_n1049), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n1017), .A2(new_n737), .B1(new_n1021), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1020), .A2(new_n1051), .ZN(G393));
  OAI21_X1  g0852(.A(new_n794), .B1(new_n441), .B2(new_n215), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n240), .A2(new_n797), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n738), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT110), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n765), .A2(G311), .B1(new_n755), .B2(G317), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT52), .Z(new_n1058));
  OAI22_X1  g0858(.A1(new_n745), .A2(new_n748), .B1(new_n751), .B2(new_n760), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(G322), .B2(new_n767), .ZN(new_n1060));
  NAND4_X1  g0860(.A1(new_n1058), .A2(new_n401), .A3(new_n780), .A4(new_n1060), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n769), .A2(G303), .B1(new_n785), .B2(G116), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT112), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(G68), .A2(new_n777), .B1(new_n752), .B2(new_n258), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n769), .A2(G50), .B1(new_n767), .B2(G143), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n785), .A2(G77), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n401), .B1(new_n779), .B2(G87), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .A4(new_n1067), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n765), .A2(G159), .B1(new_n755), .B2(G150), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(KEYINPUT111), .B(KEYINPUT51), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1069), .B(new_n1070), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n1061), .A2(new_n1063), .B1(new_n1068), .B2(new_n1071), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1072), .A2(KEYINPUT113), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1072), .A2(KEYINPUT113), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n741), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1056), .B1(new_n1073), .B2(new_n1075), .C1(new_n959), .C2(new_n792), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n976), .B2(new_n736), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n968), .A2(new_n975), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n983), .A2(new_n728), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n696), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n976), .A2(new_n1018), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1077), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(G390));
  OAI211_X1 g0883(.A(new_n906), .B(new_n908), .C1(new_n917), .C2(new_n885), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n348), .A2(new_n669), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n361), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(new_n373), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n668), .B(new_n1087), .C1(new_n717), .C2(new_n724), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1088), .A2(new_n835), .A3(new_n914), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n913), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n893), .A2(new_n875), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1084), .A2(new_n1092), .ZN(new_n1093));
  AND3_X1   g0893(.A1(new_n886), .A2(new_n877), .A3(G330), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT114), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n715), .A2(new_n886), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(KEYINPUT114), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1093), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n1084), .A2(new_n1092), .A3(new_n1095), .A4(new_n1094), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n897), .A2(KEYINPUT115), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT115), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n715), .A2(new_n1103), .A3(new_n433), .ZN(new_n1104));
  AND2_X1   g0904(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n884), .A2(new_n885), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(new_n715), .B2(new_n838), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1088), .A2(new_n835), .ZN(new_n1108));
  NOR3_X1   g0908(.A1(new_n1107), .A2(new_n1094), .A3(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n877), .A2(G330), .A3(new_n838), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n915), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n1111), .A2(new_n1097), .B1(new_n835), .B2(new_n916), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n904), .B(new_n1105), .C1(new_n1109), .C2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1101), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1099), .A2(new_n1113), .A3(new_n1100), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1115), .A2(new_n695), .A3(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n906), .A2(new_n789), .A3(new_n908), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n738), .B1(new_n258), .B2(new_n833), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT116), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n777), .A2(new_n1036), .ZN(new_n1121));
  XOR2_X1   g0921(.A(new_n1121), .B(KEYINPUT53), .Z(new_n1122));
  XOR2_X1   g0922(.A(KEYINPUT54), .B(G143), .Z(new_n1123));
  AOI22_X1  g0923(.A1(new_n752), .A2(new_n1123), .B1(new_n779), .B2(G50), .ZN(new_n1124));
  INV_X1    g0924(.A(G128), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1122), .B(new_n1124), .C1(new_n1125), .C2(new_n756), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(G132), .A2(new_n765), .B1(new_n769), .B2(new_n938), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n785), .A2(G159), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n401), .B1(new_n767), .B2(G125), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1127), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(G116), .A2(new_n765), .B1(new_n769), .B2(G107), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n1131), .B1(new_n441), .B2(new_n751), .C1(new_n748), .C2(new_n756), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n275), .B1(new_n777), .B2(G87), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n767), .A2(G294), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1133), .A2(new_n822), .A3(new_n1066), .A4(new_n1134), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n1126), .A2(new_n1130), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1120), .B1(new_n1136), .B2(new_n741), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n1101), .A2(new_n737), .B1(new_n1118), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1117), .A2(new_n1138), .ZN(G378));
  INV_X1    g0939(.A(KEYINPUT119), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n902), .A2(new_n903), .A3(new_n1102), .A4(new_n1104), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(new_n1101), .B2(new_n1114), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n325), .A2(new_n666), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n297), .A2(KEYINPUT118), .A3(new_n330), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(KEYINPUT118), .B1(new_n297), .B2(new_n330), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1143), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1146), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1143), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1148), .A2(new_n1149), .A3(new_n1144), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1147), .A2(new_n1150), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1147), .A2(new_n1150), .A3(new_n1152), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  AND4_X1   g0956(.A1(G330), .A2(new_n1156), .A3(new_n889), .A4(new_n895), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1156), .B1(new_n899), .B2(G330), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n919), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1156), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n896), .A2(new_n1160), .ZN(new_n1161));
  AND2_X1   g0961(.A1(new_n918), .A2(new_n911), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n899), .A2(G330), .A3(new_n1156), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1161), .A2(new_n910), .A3(new_n1162), .A4(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1159), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT57), .ZN(new_n1166));
  NOR3_X1   g0966(.A1(new_n1142), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1140), .B1(new_n1167), .B2(new_n696), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1113), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1164), .B(new_n1159), .C1(new_n1169), .C2(new_n1141), .ZN(new_n1170));
  OAI211_X1 g0970(.A(KEYINPUT119), .B(new_n695), .C1(new_n1170), .C2(new_n1166), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1141), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1115), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1165), .ZN(new_n1174));
  AOI21_X1  g0974(.A(KEYINPUT57), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1168), .A2(new_n1171), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1174), .A2(new_n737), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n739), .B1(new_n202), .B2(new_n832), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n275), .A2(G41), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n278), .B2(new_n745), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n756), .A2(new_n436), .B1(new_n764), .B2(new_n351), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n1181), .B(new_n1182), .C1(G68), .C2(new_n785), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n344), .A2(new_n752), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n779), .A2(G58), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n769), .A2(G97), .B1(new_n767), .B2(G283), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .A4(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n1188), .A2(KEYINPUT58), .B1(new_n1180), .B2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT117), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1188), .A2(KEYINPUT58), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n755), .A2(G125), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n777), .A2(new_n1123), .B1(new_n752), .B2(G137), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(G128), .A2(new_n765), .B1(new_n769), .B2(G132), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n785), .A2(G150), .ZN(new_n1197));
  AND4_X1   g0997(.A1(new_n1194), .A2(new_n1195), .A3(new_n1196), .A4(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT59), .ZN(new_n1199));
  OR2_X1    g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n779), .A2(G159), .ZN(new_n1202));
  AOI211_X1 g1002(.A(G33), .B(G41), .C1(new_n767), .C2(G124), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1200), .A2(new_n1201), .A3(new_n1202), .A4(new_n1203), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1192), .A2(new_n1193), .A3(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1190), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1205), .B1(KEYINPUT117), .B2(new_n1206), .ZN(new_n1207));
  OAI221_X1 g1007(.A(new_n1179), .B1(new_n742), .B2(new_n1207), .C1(new_n1160), .C2(new_n790), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1178), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1177), .A2(new_n1210), .ZN(G375));
  NAND2_X1  g1011(.A1(new_n916), .A2(new_n835), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1212), .B1(new_n1107), .B2(new_n1094), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1111), .A2(new_n1097), .A3(new_n835), .A4(new_n1088), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n736), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  AND2_X1   g1015(.A1(new_n1215), .A2(KEYINPUT120), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n756), .A2(new_n760), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n751), .A2(new_n351), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n745), .A2(new_n441), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n764), .A2(new_n748), .ZN(new_n1220));
  NOR4_X1   g1020(.A1(new_n1217), .A2(new_n1218), .A3(new_n1219), .A4(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n275), .B1(new_n779), .B2(G77), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n769), .A2(G116), .B1(new_n767), .B2(G303), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1221), .A2(new_n1035), .A3(new_n1222), .A4(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  AND2_X1   g1025(.A1(new_n1225), .A2(KEYINPUT121), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n755), .A2(G132), .B1(new_n767), .B2(G128), .ZN(new_n1227));
  AND3_X1   g1027(.A1(new_n1227), .A2(new_n275), .A3(new_n1185), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n765), .A2(new_n938), .B1(new_n752), .B2(G150), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(G159), .A2(new_n777), .B1(new_n769), .B2(new_n1123), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n785), .A2(G50), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1228), .A2(new_n1229), .A3(new_n1230), .A4(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1232), .B1(new_n1225), .B2(KEYINPUT121), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n741), .B1(new_n1226), .B2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n739), .B1(new_n312), .B2(new_n832), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1234), .B(new_n1235), .C1(new_n1106), .C2(new_n790), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n1215), .B2(KEYINPUT120), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1216), .A2(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1141), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1113), .A2(new_n986), .A3(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1238), .A2(new_n1240), .ZN(G381));
  OAI21_X1  g1041(.A(new_n695), .B1(new_n1170), .B2(new_n1166), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1175), .B1(new_n1242), .B2(new_n1140), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1209), .B1(new_n1243), .B2(new_n1171), .ZN(new_n1244));
  INV_X1    g1044(.A(G378), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1082), .B(new_n951), .C1(new_n987), .C2(new_n1013), .ZN(new_n1246));
  INV_X1    g1046(.A(G396), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1019), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n695), .B1(new_n983), .B2(new_n728), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1051), .B(new_n1247), .C1(new_n1248), .C2(new_n1249), .ZN(new_n1250));
  NOR4_X1   g1050(.A1(new_n1246), .A2(G381), .A3(G384), .A4(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1244), .A2(new_n1245), .A3(new_n1251), .ZN(G407));
  NAND2_X1  g1052(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1253));
  OAI211_X1 g1053(.A(G407), .B(G213), .C1(new_n1253), .C2(G343), .ZN(new_n1254));
  XOR2_X1   g1054(.A(new_n1254), .B(KEYINPUT122), .Z(G409));
  INV_X1    g1055(.A(KEYINPUT61), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(G387), .A2(G390), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT125), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1250), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1247), .B1(new_n1020), .B2(new_n1051), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1258), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(G393), .A2(G396), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1262), .A2(KEYINPUT125), .A3(new_n1250), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1261), .A2(new_n1263), .ZN(new_n1264));
  AND3_X1   g1064(.A1(new_n1257), .A2(new_n1264), .A3(new_n1246), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1263), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1266), .B1(new_n1257), .B2(new_n1246), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1256), .B1(new_n1265), .B2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(KEYINPUT126), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT126), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n1270), .B(new_n1256), .C1(new_n1265), .C2(new_n1267), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1269), .A2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT63), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT60), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1239), .A2(new_n1274), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1141), .A2(KEYINPUT60), .A3(new_n1213), .A4(new_n1214), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1275), .A2(new_n695), .A3(new_n1113), .A4(new_n1276), .ZN(new_n1277));
  AND3_X1   g1077(.A1(new_n1238), .A2(G384), .A3(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(G384), .B1(new_n1238), .B2(new_n1277), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(G213), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1281), .A2(G343), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1209), .A2(G378), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1173), .A2(new_n986), .A3(new_n1174), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1282), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1280), .B(new_n1285), .C1(new_n1244), .C2(new_n1245), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1272), .B1(new_n1273), .B2(new_n1286), .ZN(new_n1287));
  OR2_X1    g1087(.A1(new_n1286), .A2(new_n1273), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1285), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT124), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1282), .A2(G2897), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1291), .B1(new_n1280), .B2(KEYINPUT123), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1279), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1238), .A2(G384), .A3(new_n1277), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1293), .A2(KEYINPUT123), .A3(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT123), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1296), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1295), .A2(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1292), .B1(new_n1291), .B2(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1289), .A2(new_n1290), .A3(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1290), .B1(new_n1289), .B2(new_n1299), .ZN(new_n1302));
  OAI211_X1 g1102(.A(new_n1287), .B(new_n1288), .C1(new_n1301), .C2(new_n1302), .ZN(new_n1303));
  AND3_X1   g1103(.A1(new_n1286), .A2(KEYINPUT127), .A3(KEYINPUT62), .ZN(new_n1304));
  AOI21_X1  g1104(.A(KEYINPUT62), .B1(new_n1286), .B2(KEYINPUT127), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1245), .B1(new_n1177), .B2(new_n1210), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1282), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1299), .B1(new_n1306), .B2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1310), .A2(new_n1256), .ZN(new_n1311));
  NOR3_X1   g1111(.A1(new_n1304), .A2(new_n1305), .A3(new_n1311), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1265), .A2(new_n1267), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1313), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1303), .B1(new_n1312), .B2(new_n1314), .ZN(G405));
  NAND2_X1  g1115(.A1(G375), .A2(G378), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(new_n1253), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(new_n1280), .ZN(new_n1318));
  OAI211_X1 g1118(.A(new_n1316), .B(new_n1253), .C1(new_n1279), .C2(new_n1278), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  XNOR2_X1  g1120(.A(new_n1320), .B(new_n1314), .ZN(G402));
endmodule


