//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 0 0 1 1 1 1 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 0 1 0 1 1 1 1 1 1 0 0 0 1 1 0 1 0 1 1 0 0 0 0 0 0 0 0 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:18 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968;
  XNOR2_X1  g000(.A(G125), .B(G140), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT16), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT16), .ZN(new_n189));
  INV_X1    g003(.A(G140), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(G125), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n188), .A2(G146), .A3(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G146), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n193), .B1(new_n194), .B2(new_n187), .ZN(new_n195));
  XOR2_X1   g009(.A(KEYINPUT24), .B(G110), .Z(new_n196));
  INV_X1    g010(.A(KEYINPUT70), .ZN(new_n197));
  XNOR2_X1  g011(.A(G119), .B(G128), .ZN(new_n198));
  OR3_X1    g012(.A1(new_n196), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n197), .B1(new_n196), .B2(new_n198), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT23), .ZN(new_n201));
  INV_X1    g015(.A(G128), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n201), .B1(G119), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G119), .ZN(new_n204));
  NOR3_X1   g018(.A1(new_n204), .A2(KEYINPUT23), .A3(G128), .ZN(new_n205));
  OAI22_X1  g019(.A1(new_n203), .A2(new_n205), .B1(G119), .B2(new_n202), .ZN(new_n206));
  OAI211_X1 g020(.A(new_n199), .B(new_n200), .C1(G110), .C2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n195), .A2(new_n207), .ZN(new_n208));
  AOI21_X1  g022(.A(G146), .B1(new_n188), .B2(new_n191), .ZN(new_n209));
  OR2_X1    g023(.A1(new_n193), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n206), .A2(G110), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n196), .A2(new_n198), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  AOI21_X1  g028(.A(KEYINPUT69), .B1(new_n210), .B2(new_n214), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n193), .A2(new_n209), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT69), .ZN(new_n217));
  NOR3_X1   g031(.A1(new_n216), .A2(new_n213), .A3(new_n217), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n208), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G953), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(G221), .A3(G234), .ZN(new_n221));
  XNOR2_X1  g035(.A(new_n221), .B(KEYINPUT71), .ZN(new_n222));
  XNOR2_X1  g036(.A(KEYINPUT22), .B(G137), .ZN(new_n223));
  XNOR2_X1  g037(.A(new_n222), .B(new_n223), .ZN(new_n224));
  OR2_X1    g038(.A1(new_n224), .A2(KEYINPUT72), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(KEYINPUT72), .ZN(new_n226));
  AND2_X1   g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n219), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G902), .ZN(new_n229));
  INV_X1    g043(.A(new_n222), .ZN(new_n230));
  AND2_X1   g044(.A1(new_n230), .A2(new_n223), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n230), .A2(new_n223), .ZN(new_n232));
  OAI221_X1 g046(.A(new_n208), .B1(new_n231), .B2(new_n232), .C1(new_n215), .C2(new_n218), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n228), .A2(new_n229), .A3(new_n233), .ZN(new_n234));
  AND2_X1   g048(.A1(KEYINPUT73), .A2(KEYINPUT25), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NOR2_X1   g050(.A1(KEYINPUT73), .A2(KEYINPUT25), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n228), .A2(new_n233), .A3(new_n229), .A4(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G217), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n240), .B1(G234), .B2(new_n229), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n236), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n241), .A2(G902), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n228), .A2(new_n233), .A3(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT74), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  AND2_X1   g060(.A1(new_n228), .A2(new_n233), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n247), .A2(KEYINPUT74), .A3(new_n243), .ZN(new_n248));
  AND3_X1   g062(.A1(new_n242), .A2(new_n246), .A3(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n204), .A2(G116), .ZN(new_n251));
  INV_X1    g065(.A(G116), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G119), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT2), .B(G113), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n254), .B(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G137), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT65), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT65), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G137), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(KEYINPUT11), .A2(G134), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G131), .ZN(new_n265));
  AOI21_X1  g079(.A(KEYINPUT11), .B1(new_n257), .B2(G134), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n257), .A2(G134), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n264), .A2(new_n265), .A3(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n262), .B1(new_n258), .B2(new_n260), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT11), .ZN(new_n271));
  INV_X1    g085(.A(G134), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n271), .B1(new_n272), .B2(G137), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(G137), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g089(.A(G131), .B1(new_n270), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n269), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n194), .A2(G143), .ZN(new_n278));
  INV_X1    g092(.A(G143), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(G146), .ZN(new_n280));
  AND2_X1   g094(.A1(KEYINPUT0), .A2(G128), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n278), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  OR2_X1    g096(.A1(KEYINPUT0), .A2(G128), .ZN(new_n283));
  NAND2_X1  g097(.A1(KEYINPUT0), .A2(G128), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g099(.A(G143), .B(G146), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n282), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n277), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n257), .A2(G134), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n290), .B1(new_n261), .B2(G134), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(G131), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT1), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n293), .B1(G143), .B2(new_n194), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n279), .A2(G146), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n194), .A2(G143), .ZN(new_n296));
  OAI22_X1  g110(.A1(new_n294), .A2(new_n202), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n278), .A2(new_n280), .A3(new_n293), .A4(G128), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n292), .A2(new_n269), .A3(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n289), .A2(new_n300), .A3(KEYINPUT30), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT64), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n282), .B(new_n302), .C1(new_n285), .C2(new_n286), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  OAI211_X1 g118(.A(new_n284), .B(new_n283), .C1(new_n295), .C2(new_n296), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n302), .B1(new_n305), .B2(new_n282), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n270), .A2(new_n275), .ZN(new_n308));
  AOI22_X1  g122(.A1(new_n308), .A2(new_n265), .B1(new_n297), .B2(new_n298), .ZN(new_n309));
  AOI22_X1  g123(.A1(new_n307), .A2(new_n277), .B1(new_n292), .B2(new_n309), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n256), .B(new_n301), .C1(new_n310), .C2(KEYINPUT30), .ZN(new_n311));
  NOR2_X1   g125(.A1(G237), .A2(G953), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G210), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n313), .B(G101), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n314), .B(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n256), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n289), .A2(new_n300), .A3(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n311), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT31), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT28), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n289), .A2(new_n300), .A3(KEYINPUT28), .A4(new_n317), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n322), .B(new_n323), .C1(new_n317), .C2(new_n310), .ZN(new_n324));
  INV_X1    g138(.A(new_n316), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT31), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n311), .A2(new_n327), .A3(new_n316), .A4(new_n318), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n320), .A2(new_n326), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(KEYINPUT66), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT66), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n320), .A2(new_n331), .A3(new_n326), .A4(new_n328), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NOR2_X1   g147(.A1(G472), .A2(G902), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT32), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n334), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n338), .B1(new_n330), .B2(new_n332), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(KEYINPUT32), .ZN(new_n340));
  INV_X1    g154(.A(G472), .ZN(new_n341));
  OR2_X1    g155(.A1(new_n324), .A2(new_n325), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n311), .A2(new_n318), .ZN(new_n343));
  AOI21_X1  g157(.A(KEYINPUT29), .B1(new_n343), .B2(new_n325), .ZN(new_n344));
  AOI21_X1  g158(.A(G902), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT67), .ZN(new_n346));
  INV_X1    g160(.A(new_n318), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n317), .B1(new_n289), .B2(new_n300), .ZN(new_n348));
  OAI21_X1  g162(.A(KEYINPUT28), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n346), .B1(new_n349), .B2(new_n322), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n322), .A2(new_n346), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n351), .A2(KEYINPUT29), .A3(new_n316), .A4(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n341), .B1(new_n345), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n337), .A2(new_n340), .A3(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT68), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(KEYINPUT32), .B1(new_n333), .B2(new_n334), .ZN(new_n359));
  AOI211_X1 g173(.A(new_n336), .B(new_n338), .C1(new_n330), .C2(new_n332), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(KEYINPUT68), .A3(new_n355), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n250), .B1(new_n358), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(G214), .B1(G237), .B2(G902), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(G210), .B1(G237), .B2(G902), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT79), .ZN(new_n368));
  INV_X1    g182(.A(G104), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(G107), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n369), .A2(G107), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT75), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n372), .A2(KEYINPUT3), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n370), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G107), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G104), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT3), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT75), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n372), .A2(KEYINPUT3), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n376), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(G101), .B1(new_n374), .B2(new_n380), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n375), .A2(G104), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n382), .B1(new_n376), .B2(new_n378), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n377), .A2(KEYINPUT75), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n371), .B1(new_n373), .B2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(G101), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n383), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n381), .A2(new_n387), .A3(KEYINPUT4), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT4), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n389), .B(G101), .C1(new_n374), .C2(new_n380), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n388), .A2(new_n256), .A3(new_n390), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n254), .A2(new_n255), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n251), .A2(new_n253), .A3(KEYINPUT5), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n251), .A2(KEYINPUT5), .ZN(new_n394));
  INV_X1    g208(.A(G113), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n392), .B1(new_n393), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(G101), .B1(new_n382), .B2(new_n371), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n397), .A2(new_n398), .A3(new_n387), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n391), .A2(new_n399), .ZN(new_n400));
  XOR2_X1   g214(.A(G110), .B(G122), .Z(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n401), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n391), .A2(new_n399), .A3(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n402), .A2(KEYINPUT6), .A3(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT6), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n400), .A2(new_n406), .A3(new_n401), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n368), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  AND2_X1   g222(.A1(new_n404), .A2(KEYINPUT6), .ZN(new_n409));
  AOI21_X1  g223(.A(KEYINPUT79), .B1(new_n409), .B2(new_n402), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n287), .A2(G125), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n411), .B1(G125), .B2(new_n299), .ZN(new_n412));
  INV_X1    g226(.A(G224), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n413), .A2(G953), .ZN(new_n414));
  XOR2_X1   g228(.A(new_n412), .B(new_n414), .Z(new_n415));
  NOR3_X1   g229(.A1(new_n408), .A2(new_n410), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n387), .A2(new_n398), .ZN(new_n417));
  XOR2_X1   g231(.A(new_n417), .B(new_n397), .Z(new_n418));
  XOR2_X1   g232(.A(new_n401), .B(KEYINPUT8), .Z(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT7), .ZN(new_n421));
  OR3_X1    g235(.A1(new_n412), .A2(new_n421), .A3(new_n414), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n412), .B1(new_n421), .B2(new_n414), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT80), .ZN(new_n424));
  OR2_X1    g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n423), .A2(new_n424), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n420), .A2(new_n422), .A3(new_n425), .A4(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n404), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n229), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n367), .B1(new_n416), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n415), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n405), .A2(new_n368), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n405), .A2(new_n407), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n431), .B(new_n432), .C1(new_n433), .C2(new_n368), .ZN(new_n434));
  INV_X1    g248(.A(new_n429), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n434), .A2(new_n435), .A3(new_n366), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n365), .B1(new_n430), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n312), .A2(G214), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT82), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n438), .A2(new_n439), .A3(new_n279), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n312), .B(G214), .C1(KEYINPUT82), .C2(G143), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT18), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n440), .B(new_n441), .C1(new_n442), .C2(new_n265), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n187), .B(new_n194), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n440), .A2(new_n441), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(G131), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n443), .B(new_n444), .C1(new_n446), .C2(new_n442), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n440), .A2(new_n265), .A3(new_n441), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n265), .B1(new_n440), .B2(new_n441), .ZN(new_n449));
  NOR3_X1   g263(.A1(new_n448), .A2(new_n449), .A3(KEYINPUT17), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n216), .B1(new_n450), .B2(KEYINPUT85), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT17), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n440), .A2(new_n265), .A3(new_n441), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n446), .A2(KEYINPUT85), .A3(new_n452), .A4(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT84), .ZN(new_n455));
  AND3_X1   g269(.A1(new_n449), .A2(new_n455), .A3(KEYINPUT17), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n455), .B1(new_n449), .B2(KEYINPUT17), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n454), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n447), .B1(new_n451), .B2(new_n458), .ZN(new_n459));
  XNOR2_X1  g273(.A(G113), .B(G122), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n460), .B(G104), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n461), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n463), .B(new_n447), .C1(new_n451), .C2(new_n458), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n229), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(G475), .ZN(new_n467));
  XNOR2_X1  g281(.A(KEYINPUT90), .B(G952), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n468), .A2(G953), .ZN(new_n469));
  NAND2_X1  g283(.A1(G234), .A2(G237), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n470), .A2(G902), .A3(G953), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(KEYINPUT21), .B(G898), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT19), .ZN(new_n477));
  OR2_X1    g291(.A1(new_n187), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n187), .A2(new_n477), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n478), .A2(new_n479), .A3(new_n194), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n480), .B(new_n192), .C1(new_n448), .C2(new_n449), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n447), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n461), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(KEYINPUT83), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT83), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n482), .A2(new_n485), .A3(new_n461), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n484), .A2(new_n464), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT20), .ZN(new_n488));
  NOR2_X1   g302(.A1(G475), .A2(G902), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(KEYINPUT81), .B(KEYINPUT20), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n493), .B1(new_n487), .B2(new_n489), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n467), .B(new_n476), .C1(new_n491), .C2(new_n494), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n279), .A2(G128), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n202), .A2(G143), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n498), .B(new_n272), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n252), .A2(G122), .ZN(new_n500));
  INV_X1    g314(.A(G122), .ZN(new_n501));
  OAI21_X1  g315(.A(KEYINPUT86), .B1(new_n501), .B2(G116), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT86), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n503), .A2(new_n252), .A3(G122), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n500), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT14), .ZN(new_n506));
  OAI21_X1  g320(.A(G107), .B1(new_n500), .B2(new_n506), .ZN(new_n507));
  OR2_X1    g321(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n505), .A2(new_n507), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n499), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT87), .ZN(new_n511));
  AOI21_X1  g325(.A(KEYINPUT13), .B1(new_n279), .B2(G128), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n511), .B1(new_n512), .B2(new_n496), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n202), .A2(G143), .ZN(new_n514));
  OAI211_X1 g328(.A(KEYINPUT87), .B(new_n514), .C1(new_n497), .C2(KEYINPUT13), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n497), .A2(KEYINPUT13), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n513), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT88), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n517), .A2(new_n518), .A3(G134), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n505), .B(new_n375), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n498), .A2(new_n272), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n518), .B1(new_n517), .B2(G134), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n510), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  XOR2_X1   g338(.A(KEYINPUT9), .B(G234), .Z(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  NOR3_X1   g340(.A1(new_n526), .A2(new_n240), .A3(G953), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n524), .A2(new_n528), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n527), .B(new_n510), .C1(new_n522), .C2(new_n523), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n529), .A2(KEYINPUT89), .A3(new_n530), .ZN(new_n531));
  OR3_X1    g345(.A1(new_n524), .A2(KEYINPUT89), .A3(new_n528), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n531), .A2(new_n532), .A3(new_n229), .ZN(new_n533));
  INV_X1    g347(.A(G478), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n534), .A2(KEYINPUT15), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n533), .B(new_n535), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n495), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(G221), .B1(new_n526), .B2(G902), .ZN(new_n538));
  AND3_X1   g352(.A1(new_n387), .A2(new_n299), .A3(new_n398), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n299), .B1(new_n398), .B2(new_n387), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n277), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT76), .ZN(new_n542));
  AOI21_X1  g356(.A(KEYINPUT12), .B1(new_n277), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n299), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n417), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n387), .A2(new_n299), .A3(new_n398), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n543), .B1(new_n549), .B2(new_n277), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n545), .A2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT78), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n388), .A2(new_n288), .A3(new_n390), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT10), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n548), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n277), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n387), .A2(new_n299), .A3(KEYINPUT10), .A4(new_n398), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n553), .A2(new_n555), .A3(new_n556), .A4(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(G110), .B(G140), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n220), .A2(G227), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n559), .B(new_n560), .ZN(new_n561));
  AND2_X1   g375(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n551), .A2(new_n552), .A3(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n553), .A2(new_n555), .A3(new_n557), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n277), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n558), .ZN(new_n566));
  INV_X1    g380(.A(new_n561), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n541), .A2(new_n544), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n549), .A2(new_n277), .A3(new_n543), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n558), .A2(new_n561), .ZN(new_n572));
  OAI21_X1  g386(.A(KEYINPUT78), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n563), .A2(new_n568), .A3(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(G469), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n574), .A2(new_n575), .A3(new_n229), .ZN(new_n576));
  NAND2_X1  g390(.A1(G469), .A2(G902), .ZN(new_n577));
  OR2_X1    g391(.A1(new_n572), .A2(KEYINPUT77), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n572), .A2(KEYINPUT77), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n578), .A2(new_n565), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n551), .A2(new_n558), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n567), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n576), .B(new_n577), .C1(new_n575), .C2(new_n583), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n437), .A2(new_n537), .A3(new_n538), .A4(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT91), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n584), .A2(new_n538), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n589), .A2(KEYINPUT91), .A3(new_n437), .A4(new_n537), .ZN(new_n590));
  AND2_X1   g404(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n363), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(KEYINPUT92), .B(G101), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n592), .B(new_n593), .ZN(G3));
  AOI21_X1  g408(.A(new_n341), .B1(new_n333), .B2(new_n229), .ZN(new_n595));
  OR2_X1    g409(.A1(new_n595), .A2(new_n339), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n487), .A2(new_n489), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n492), .ZN(new_n598));
  AOI22_X1  g412(.A1(new_n598), .A2(new_n490), .B1(G475), .B2(new_n466), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT33), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n531), .A2(new_n532), .A3(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n529), .A2(KEYINPUT33), .A3(new_n530), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n534), .A2(G902), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  AOI22_X1  g418(.A1(new_n604), .A2(KEYINPUT93), .B1(new_n534), .B2(new_n533), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT93), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n601), .A2(new_n606), .A3(new_n602), .A4(new_n603), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n599), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n608), .A2(new_n437), .A3(new_n476), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n249), .A2(new_n584), .A3(new_n538), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n596), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(KEYINPUT94), .ZN(new_n612));
  XNOR2_X1  g426(.A(KEYINPUT34), .B(G104), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(G6));
  NOR2_X1   g428(.A1(new_n596), .A2(new_n610), .ZN(new_n615));
  XOR2_X1   g429(.A(new_n476), .B(KEYINPUT95), .Z(new_n616));
  AND2_X1   g430(.A1(new_n437), .A2(new_n616), .ZN(new_n617));
  XOR2_X1   g431(.A(new_n533), .B(new_n535), .Z(new_n618));
  NOR2_X1   g432(.A1(new_n597), .A2(new_n492), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n467), .B1(new_n619), .B2(new_n494), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n615), .A2(new_n617), .A3(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(KEYINPUT35), .B(G107), .Z(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G9));
  INV_X1    g438(.A(KEYINPUT97), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n225), .A2(new_n226), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT96), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT36), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n627), .B1(new_n626), .B2(new_n628), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n219), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n631), .ZN(new_n633));
  INV_X1    g447(.A(new_n219), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n633), .A2(new_n634), .A3(new_n629), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n632), .A2(new_n635), .A3(new_n243), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n242), .A2(new_n625), .A3(new_n636), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n625), .B1(new_n242), .B2(new_n636), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n639), .A2(new_n595), .A3(new_n339), .ZN(new_n640));
  AND3_X1   g454(.A1(new_n640), .A2(new_n587), .A3(new_n590), .ZN(new_n641));
  XNOR2_X1  g455(.A(KEYINPUT37), .B(G110), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G12));
  NAND2_X1  g457(.A1(new_n358), .A2(new_n362), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n471), .B1(G900), .B2(new_n472), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n618), .A2(new_n620), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(KEYINPUT98), .ZN(new_n648));
  INV_X1    g462(.A(new_n437), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n649), .A2(new_n588), .ZN(new_n650));
  INV_X1    g464(.A(new_n639), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n644), .A2(new_n648), .A3(new_n650), .A4(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G128), .ZN(G30));
  XNOR2_X1  g467(.A(new_n645), .B(KEYINPUT39), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n589), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(new_n655), .B(KEYINPUT40), .Z(new_n656));
  OAI21_X1  g470(.A(new_n325), .B1(new_n347), .B2(new_n348), .ZN(new_n657));
  AND3_X1   g471(.A1(new_n319), .A2(KEYINPUT100), .A3(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(KEYINPUT100), .B1(new_n319), .B2(new_n657), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n658), .A2(G902), .A3(new_n659), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n361), .B1(new_n341), .B2(new_n660), .ZN(new_n661));
  NOR3_X1   g475(.A1(new_n618), .A2(new_n599), .A3(new_n365), .ZN(new_n662));
  AND2_X1   g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n430), .A2(new_n436), .ZN(new_n664));
  XNOR2_X1  g478(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n665));
  XOR2_X1   g479(.A(new_n664), .B(new_n665), .Z(new_n666));
  NAND2_X1  g480(.A1(new_n242), .A2(new_n636), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n656), .A2(new_n663), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G143), .ZN(G45));
  NAND3_X1  g484(.A1(new_n608), .A2(new_n437), .A3(new_n645), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT101), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n673), .A2(new_n644), .A3(new_n589), .A4(new_n651), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G146), .ZN(G48));
  NAND2_X1  g489(.A1(new_n574), .A2(new_n229), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(G469), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n677), .A2(new_n538), .A3(new_n576), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT102), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n677), .A2(KEYINPUT102), .A3(new_n538), .A4(new_n576), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n682), .A2(new_n609), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n363), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(KEYINPUT41), .B(G113), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G15));
  NAND3_X1  g500(.A1(new_n621), .A2(new_n437), .A3(new_n616), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n682), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(KEYINPUT68), .B1(new_n361), .B2(new_n355), .ZN(new_n689));
  NOR4_X1   g503(.A1(new_n359), .A2(new_n360), .A3(new_n357), .A4(new_n354), .ZN(new_n690));
  OAI211_X1 g504(.A(new_n688), .B(new_n249), .C1(new_n689), .C2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G116), .ZN(G18));
  AND4_X1   g506(.A1(new_n437), .A2(new_n680), .A3(new_n537), .A4(new_n681), .ZN(new_n693));
  OAI211_X1 g507(.A(new_n651), .B(new_n693), .C1(new_n689), .C2(new_n690), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G119), .ZN(G21));
  INV_X1    g509(.A(new_n352), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n325), .B1(new_n350), .B2(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n697), .A2(new_n320), .A3(new_n328), .ZN(new_n698));
  AND2_X1   g512(.A1(new_n698), .A2(new_n334), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n595), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n700), .A2(new_n249), .A3(new_n680), .A4(new_n681), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n618), .A2(new_n599), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n617), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(new_n501), .ZN(G24));
  NAND2_X1  g519(.A1(new_n700), .A2(new_n667), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n608), .A2(new_n645), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n682), .A2(new_n649), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G125), .ZN(G27));
  INV_X1    g525(.A(KEYINPUT42), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n664), .A2(new_n365), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n581), .A2(KEYINPUT103), .A3(new_n567), .ZN(new_n714));
  AOI21_X1  g528(.A(KEYINPUT103), .B1(new_n581), .B2(new_n567), .ZN(new_n715));
  OAI211_X1 g529(.A(G469), .B(new_n580), .C1(new_n714), .C2(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n716), .A2(new_n576), .A3(new_n577), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n713), .A2(new_n538), .A3(new_n717), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n718), .A2(new_n707), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n250), .B1(new_n361), .B2(new_n355), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n712), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  AOI211_X1 g535(.A(new_n250), .B(new_n718), .C1(new_n358), .C2(new_n362), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n707), .A2(KEYINPUT42), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n721), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G131), .ZN(G33));
  INV_X1    g539(.A(KEYINPUT104), .ZN(new_n726));
  INV_X1    g540(.A(new_n718), .ZN(new_n727));
  OAI211_X1 g541(.A(new_n249), .B(new_n727), .C1(new_n689), .C2(new_n690), .ZN(new_n728));
  INV_X1    g542(.A(new_n648), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n726), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n363), .A2(KEYINPUT104), .A3(new_n648), .A4(new_n727), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G134), .ZN(G36));
  NAND2_X1  g547(.A1(new_n605), .A2(new_n607), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(new_n599), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(KEYINPUT43), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n737), .A2(new_n596), .A3(new_n667), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT44), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n713), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  OR2_X1    g554(.A1(new_n740), .A2(KEYINPUT105), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(KEYINPUT105), .ZN(new_n742));
  OAI211_X1 g556(.A(KEYINPUT45), .B(new_n580), .C1(new_n714), .C2(new_n715), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT45), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n583), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n743), .A2(G469), .A3(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n746), .A2(KEYINPUT46), .A3(new_n577), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(new_n576), .ZN(new_n748));
  AOI21_X1  g562(.A(KEYINPUT46), .B1(new_n746), .B2(new_n577), .ZN(new_n749));
  OR2_X1    g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n750), .A2(new_n538), .A3(new_n654), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n751), .B1(new_n738), .B2(new_n739), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n741), .A2(new_n742), .A3(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G137), .ZN(G39));
  NAND2_X1  g568(.A1(new_n750), .A2(new_n538), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT106), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT47), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n755), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n756), .A2(new_n757), .ZN(new_n760));
  MUX2_X1   g574(.A(new_n759), .B(new_n755), .S(new_n760), .Z(new_n761));
  NAND2_X1  g575(.A1(new_n713), .A2(new_n250), .ZN(new_n762));
  NOR4_X1   g576(.A1(new_n761), .A2(new_n644), .A3(new_n707), .A4(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(new_n190), .ZN(G42));
  INV_X1    g578(.A(new_n682), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n713), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(KEYINPUT114), .ZN(new_n767));
  AND4_X1   g581(.A1(new_n470), .A2(new_n767), .A3(new_n469), .A4(new_n737), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n720), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT116), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n768), .A2(KEYINPUT116), .A3(new_n720), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n771), .A2(KEYINPUT48), .A3(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT48), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n769), .A2(new_n770), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n700), .A2(new_n249), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n736), .A2(new_n471), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n709), .ZN(new_n778));
  OR2_X1    g592(.A1(new_n661), .A2(new_n250), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n779), .A2(new_n471), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n767), .A2(new_n780), .ZN(new_n781));
  AOI211_X1 g595(.A(G953), .B(new_n468), .C1(new_n781), .C2(new_n608), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n773), .A2(new_n775), .A3(new_n778), .A4(new_n782), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n781), .A2(new_n599), .A3(new_n607), .A4(new_n605), .ZN(new_n784));
  OR2_X1    g598(.A1(new_n784), .A2(KEYINPUT115), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n666), .A2(new_n365), .A3(new_n765), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(KEYINPUT113), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n777), .ZN(new_n788));
  XOR2_X1   g602(.A(new_n788), .B(KEYINPUT50), .Z(new_n789));
  INV_X1    g603(.A(new_n706), .ZN(new_n790));
  AOI22_X1  g604(.A1(new_n784), .A2(KEYINPUT115), .B1(new_n768), .B2(new_n790), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n785), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n677), .A2(new_n576), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(KEYINPUT107), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n761), .B1(new_n538), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n796), .A2(new_n713), .A3(new_n777), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n792), .A2(new_n797), .ZN(new_n798));
  AOI21_X1  g612(.A(KEYINPUT51), .B1(new_n792), .B2(KEYINPUT112), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n798), .A2(new_n799), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n783), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n708), .A2(new_n727), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n589), .B(new_n651), .C1(new_n689), .C2(new_n690), .ZN(new_n804));
  INV_X1    g618(.A(new_n620), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n713), .A2(new_n618), .A3(new_n805), .A4(new_n645), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n803), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n732), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT109), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n807), .B1(new_n730), .B2(new_n731), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(KEYINPUT109), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n437), .A2(new_n616), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n599), .A2(new_n536), .ZN(new_n815));
  OR3_X1    g629(.A1(new_n814), .A2(KEYINPUT108), .A3(new_n815), .ZN(new_n816));
  OAI21_X1  g630(.A(KEYINPUT108), .B1(new_n814), .B2(new_n815), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n816), .A2(new_n615), .A3(new_n817), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n691), .A2(new_n694), .A3(new_n818), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n249), .A2(new_n538), .A3(new_n584), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n595), .A2(new_n339), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n617), .A2(new_n820), .A3(new_n608), .A4(new_n821), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n822), .B1(new_n701), .B2(new_n703), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n823), .B1(new_n363), .B2(new_n591), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n641), .B1(new_n363), .B2(new_n683), .ZN(new_n825));
  AND4_X1   g639(.A1(new_n724), .A2(new_n819), .A3(new_n824), .A4(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n811), .A2(new_n813), .A3(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT53), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n667), .A2(new_n646), .ZN(new_n829));
  AND4_X1   g643(.A1(new_n664), .A2(new_n717), .A3(new_n538), .A4(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n661), .A2(new_n830), .A3(new_n662), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n674), .A2(new_n652), .A3(new_n710), .A4(new_n831), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(KEYINPUT52), .ZN(new_n833));
  OR3_X1    g647(.A1(new_n827), .A2(new_n828), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(KEYINPUT52), .B1(new_n832), .B2(KEYINPUT110), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n832), .A2(KEYINPUT110), .A3(KEYINPUT52), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n827), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n834), .B1(KEYINPUT53), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(KEYINPUT54), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n828), .B1(new_n827), .B2(new_n833), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n836), .A2(new_n835), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n724), .A2(new_n819), .A3(new_n824), .A4(new_n825), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n842), .B1(KEYINPUT109), .B2(new_n812), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n841), .A2(new_n843), .A3(KEYINPUT53), .A4(new_n811), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n845), .A2(KEYINPUT54), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT111), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n839), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n839), .A2(new_n847), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(KEYINPUT111), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n802), .A2(new_n849), .A3(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n852), .B1(G952), .B2(G953), .ZN(new_n853));
  INV_X1    g667(.A(new_n779), .ZN(new_n854));
  OR2_X1    g668(.A1(new_n795), .A2(KEYINPUT49), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n735), .B1(new_n795), .B2(KEYINPUT49), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n666), .A2(new_n364), .A3(new_n538), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n854), .A2(new_n855), .A3(new_n856), .A4(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n853), .A2(new_n858), .ZN(G75));
  NOR2_X1   g673(.A1(new_n220), .A2(G952), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT119), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n862), .B1(new_n845), .B2(G902), .ZN(new_n863));
  AOI211_X1 g677(.A(KEYINPUT119), .B(new_n229), .C1(new_n840), .C2(new_n844), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n865), .A2(new_n366), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n415), .B1(new_n408), .B2(new_n410), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n434), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n868), .B(KEYINPUT55), .ZN(new_n869));
  OR2_X1    g683(.A1(new_n869), .A2(KEYINPUT56), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n861), .B1(new_n866), .B2(new_n870), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n845), .A2(G210), .A3(G902), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT117), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT56), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n875), .B1(new_n872), .B2(new_n873), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n869), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT118), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  OAI211_X1 g693(.A(KEYINPUT118), .B(new_n869), .C1(new_n874), .C2(new_n876), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n871), .B1(new_n879), .B2(new_n880), .ZN(G51));
  INV_X1    g695(.A(new_n746), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n882), .B1(new_n863), .B2(new_n864), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(KEYINPUT120), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT120), .ZN(new_n885));
  OAI211_X1 g699(.A(new_n885), .B(new_n882), .C1(new_n863), .C2(new_n864), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n577), .B(KEYINPUT57), .Z(new_n887));
  INV_X1    g701(.A(KEYINPUT54), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n888), .B1(new_n840), .B2(new_n844), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n887), .B1(new_n846), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(new_n574), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n884), .A2(new_n886), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(new_n861), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(KEYINPUT121), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT121), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n892), .A2(new_n895), .A3(new_n861), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n894), .A2(new_n896), .ZN(G54));
  NAND2_X1  g711(.A1(KEYINPUT58), .A2(G475), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n898), .B(KEYINPUT122), .Z(new_n899));
  OAI21_X1  g713(.A(new_n899), .B1(new_n863), .B2(new_n864), .ZN(new_n900));
  INV_X1    g714(.A(new_n487), .ZN(new_n901));
  OR2_X1    g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n860), .B1(new_n900), .B2(new_n901), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n902), .A2(new_n903), .ZN(G60));
  NOR2_X1   g718(.A1(new_n846), .A2(new_n889), .ZN(new_n905));
  NAND2_X1  g719(.A1(G478), .A2(G902), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n906), .B(KEYINPUT59), .Z(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n601), .A2(new_n602), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n861), .B1(new_n905), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n851), .A2(new_n849), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(new_n908), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n601), .A2(new_n602), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n910), .B1(new_n912), .B2(new_n913), .ZN(G63));
  NAND2_X1  g728(.A1(G217), .A2(G902), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT60), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n916), .B1(new_n840), .B2(new_n844), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n632), .A2(new_n635), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n247), .B(KEYINPUT123), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n920), .B(new_n861), .C1(new_n917), .C2(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(KEYINPUT61), .B1(new_n920), .B2(KEYINPUT124), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n922), .B(new_n923), .ZN(G66));
  NAND3_X1  g738(.A1(new_n819), .A2(new_n824), .A3(new_n825), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(new_n220), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT125), .ZN(new_n927));
  OAI21_X1  g741(.A(G953), .B1(new_n474), .B2(new_n413), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI22_X1  g743(.A1(new_n408), .A2(new_n410), .B1(G898), .B2(new_n220), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n929), .B(new_n930), .ZN(G69));
  OAI21_X1  g745(.A(new_n301), .B1(new_n310), .B2(KEYINPUT30), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n478), .A2(new_n479), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n933), .B(KEYINPUT126), .Z(new_n934));
  XNOR2_X1  g748(.A(new_n932), .B(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(G900), .A2(G953), .ZN(new_n936));
  INV_X1    g750(.A(new_n753), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n937), .A2(new_n763), .ZN(new_n938));
  INV_X1    g752(.A(new_n751), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n939), .A2(new_n437), .A3(new_n702), .A4(new_n720), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT127), .ZN(new_n941));
  INV_X1    g755(.A(new_n724), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n674), .A2(new_n652), .A3(new_n710), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n938), .A2(new_n732), .A3(new_n941), .A4(new_n944), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n935), .B(new_n936), .C1(new_n945), .C2(G953), .ZN(new_n946));
  INV_X1    g760(.A(new_n655), .ZN(new_n947));
  INV_X1    g761(.A(new_n608), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n948), .A2(new_n815), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n363), .A2(new_n947), .A3(new_n713), .A4(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n669), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n951), .A2(new_n943), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT62), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n938), .A2(new_n950), .A3(new_n953), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n954), .A2(new_n220), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n946), .B1(new_n955), .B2(new_n935), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n220), .B1(G227), .B2(G900), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n956), .B(new_n957), .ZN(G72));
  NAND2_X1  g772(.A1(G472), .A2(G902), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT63), .Z(new_n960));
  OAI21_X1  g774(.A(new_n960), .B1(new_n945), .B2(new_n925), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n343), .A2(new_n316), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n860), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n343), .A2(new_n325), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n319), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n838), .A2(new_n960), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n960), .B1(new_n954), .B2(new_n925), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n967), .A2(new_n316), .A3(new_n343), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n963), .A2(new_n966), .A3(new_n968), .ZN(G57));
endmodule


