//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 1 0 0 0 1 1 0 0 0 0 0 0 1 1 0 0 0 0 1 0 1 0 1 0 1 0 0 0 1 1 0 0 0 0 0 1 1 1 0 1 0 0 0 0 1 0 0 0 0 1 1 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:52 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1305,
    new_n1306, new_n1307;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n202), .A2(new_n203), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G50), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n208), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT64), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n210), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n213), .B(new_n219), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G250), .B(G257), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G264), .B(G270), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT65), .Z(new_n232));
  XOR2_X1   g0032(.A(G238), .B(G244), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT2), .B(G226), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n232), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n201), .A2(G68), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n203), .A2(G50), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n240), .B(new_n245), .ZN(G351));
  XNOR2_X1  g0046(.A(KEYINPUT3), .B(G33), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n247), .A2(G223), .A3(G1698), .ZN(new_n248));
  INV_X1    g0048(.A(G77), .ZN(new_n249));
  INV_X1    g0049(.A(G222), .ZN(new_n250));
  OR2_X1    g0050(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n251));
  NAND2_X1  g0051(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n252));
  AND2_X1   g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  OAI211_X1 g0054(.A(new_n251), .B(new_n252), .C1(new_n253), .C2(new_n254), .ZN(new_n255));
  OAI221_X1 g0055(.A(new_n248), .B1(new_n249), .B2(new_n247), .C1(new_n250), .C2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(G1), .A3(G13), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G274), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n261), .A2(G1), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(KEYINPUT66), .A2(G41), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(KEYINPUT66), .A2(G41), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G45), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n263), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n270));
  AND2_X1   g0070(.A1(new_n258), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n269), .B1(G226), .B2(new_n271), .ZN(new_n272));
  AND3_X1   g0072(.A1(new_n260), .A2(G190), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G200), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n274), .B1(new_n260), .B2(new_n272), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT9), .ZN(new_n277));
  NAND3_X1  g0077(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n217), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n279), .B1(new_n207), .B2(G20), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G50), .ZN(new_n281));
  INV_X1    g0081(.A(G13), .ZN(new_n282));
  NOR3_X1   g0082(.A1(new_n282), .A2(new_n208), .A3(G1), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(new_n201), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  OR2_X1    g0086(.A1(KEYINPUT8), .A2(G58), .ZN(new_n287));
  NAND2_X1  g0087(.A1(KEYINPUT8), .A2(G58), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n208), .A2(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(KEYINPUT68), .ZN(new_n292));
  INV_X1    g0092(.A(G33), .ZN(new_n293));
  OR3_X1    g0093(.A1(new_n293), .A2(KEYINPUT68), .A3(G20), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n290), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT69), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n296), .A2(new_n208), .A3(new_n293), .ZN(new_n297));
  OAI21_X1  g0097(.A(KEYINPUT69), .B1(G20), .B2(G33), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  AOI22_X1  g0099(.A1(new_n299), .A2(G150), .B1(G20), .B2(new_n204), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n295), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(new_n279), .ZN(new_n302));
  AOI21_X1  g0102(.A(KEYINPUT71), .B1(new_n286), .B2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n279), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n304), .B1(new_n295), .B2(new_n300), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT71), .ZN(new_n306));
  NOR3_X1   g0106(.A1(new_n305), .A2(new_n285), .A3(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n277), .B1(new_n303), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n286), .A2(new_n302), .A3(KEYINPUT71), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n306), .B1(new_n305), .B2(new_n285), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n309), .A2(KEYINPUT9), .A3(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n276), .A2(new_n308), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(KEYINPUT10), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT10), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n276), .A2(new_n308), .A3(new_n314), .A4(new_n311), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  AND2_X1   g0116(.A1(new_n260), .A2(new_n272), .ZN(new_n317));
  OAI22_X1  g0117(.A1(new_n317), .A2(G169), .B1(new_n305), .B2(new_n285), .ZN(new_n318));
  INV_X1    g0118(.A(G179), .ZN(new_n319));
  AND2_X1   g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n280), .A2(G77), .ZN(new_n323));
  INV_X1    g0123(.A(new_n283), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n323), .B1(G77), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n290), .A2(new_n299), .ZN(new_n326));
  XOR2_X1   g0126(.A(KEYINPUT15), .B(G87), .Z(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  OAI221_X1 g0128(.A(new_n326), .B1(new_n208), .B2(new_n249), .C1(new_n291), .C2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n325), .B1(new_n329), .B2(new_n279), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n247), .A2(G238), .A3(G1698), .ZN(new_n332));
  INV_X1    g0132(.A(new_n252), .ZN(new_n333));
  NOR2_X1   g0133(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n335), .A2(G232), .A3(new_n247), .ZN(new_n336));
  INV_X1    g0136(.A(G107), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n332), .B(new_n336), .C1(new_n337), .C2(new_n247), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n259), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n269), .B1(G244), .B2(new_n271), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G190), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n331), .B1(new_n343), .B2(KEYINPUT70), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n274), .B1(new_n339), .B2(new_n340), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT70), .ZN(new_n346));
  OAI22_X1  g0146(.A1(new_n345), .A2(new_n346), .B1(new_n341), .B2(new_n342), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n339), .A2(new_n319), .A3(new_n340), .ZN(new_n348));
  INV_X1    g0148(.A(G169), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n330), .B1(new_n341), .B2(new_n349), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n344), .A2(new_n347), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n316), .A2(KEYINPUT72), .A3(new_n322), .A4(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n247), .A2(G232), .A3(G1698), .ZN(new_n353));
  NAND2_X1  g0153(.A1(G33), .A2(G97), .ZN(new_n354));
  INV_X1    g0154(.A(G226), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n353), .B(new_n354), .C1(new_n355), .C2(new_n255), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(new_n259), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT13), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n269), .B1(G238), .B2(new_n271), .ZN(new_n359));
  AND3_X1   g0159(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n358), .B1(new_n357), .B2(new_n359), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(KEYINPUT14), .B1(new_n362), .B2(new_n349), .ZN(new_n363));
  INV_X1    g0163(.A(new_n361), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT14), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n366), .A2(new_n367), .A3(G169), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n362), .A2(G179), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n363), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n299), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n294), .A2(new_n292), .A3(G77), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n304), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  OR2_X1    g0173(.A1(new_n373), .A2(KEYINPUT11), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(KEYINPUT11), .ZN(new_n375));
  OR3_X1    g0175(.A1(new_n324), .A2(KEYINPUT12), .A3(G68), .ZN(new_n376));
  OAI21_X1  g0176(.A(KEYINPUT12), .B1(new_n324), .B2(G68), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n376), .A2(new_n377), .B1(G68), .B2(new_n280), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n374), .A2(new_n375), .A3(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n364), .A2(G190), .A3(new_n365), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT73), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n362), .A2(KEYINPUT73), .A3(G190), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n379), .B1(new_n366), .B2(G200), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n370), .A2(new_n379), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(KEYINPUT7), .B1(new_n247), .B2(G20), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n253), .A2(new_n254), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT7), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(new_n389), .A3(new_n208), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n387), .A2(new_n390), .A3(G68), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT16), .ZN(new_n392));
  XNOR2_X1  g0192(.A(G58), .B(G68), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n299), .A2(G159), .B1(new_n393), .B2(G20), .ZN(new_n394));
  AND3_X1   g0194(.A1(new_n391), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n392), .B1(new_n391), .B2(new_n394), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n279), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n324), .A2(new_n304), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n289), .B1(new_n207), .B2(G20), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n399), .A2(new_n400), .B1(new_n289), .B2(new_n283), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n251), .A2(G223), .A3(new_n252), .ZN(new_n402));
  NAND2_X1  g0202(.A1(G226), .A2(G1698), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n388), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(G87), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n293), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n259), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  AND3_X1   g0207(.A1(new_n258), .A2(G232), .A3(new_n270), .ZN(new_n408));
  OAI21_X1  g0208(.A(KEYINPUT74), .B1(new_n269), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT66), .ZN(new_n410));
  INV_X1    g0210(.A(G41), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n412), .A2(new_n268), .A3(new_n264), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n262), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT74), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n258), .A2(G232), .A3(new_n270), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n407), .A2(new_n409), .A3(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n418), .A2(G190), .ZN(new_n419));
  AND3_X1   g0219(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n415), .B1(new_n414), .B2(new_n416), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(G200), .B1(new_n422), .B2(new_n407), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n397), .B(new_n401), .C1(new_n419), .C2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT17), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n418), .A2(new_n274), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n427), .B1(G190), .B2(new_n418), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n428), .A2(KEYINPUT17), .A3(new_n397), .A4(new_n401), .ZN(new_n429));
  AND2_X1   g0229(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT75), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n349), .B1(new_n422), .B2(new_n407), .ZN(new_n432));
  AND4_X1   g0232(.A1(G179), .A2(new_n407), .A3(new_n409), .A4(new_n417), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n431), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n397), .A2(new_n401), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n418), .A2(G169), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n422), .A2(G179), .A3(new_n407), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n436), .A2(new_n437), .A3(KEYINPUT75), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n434), .A2(new_n435), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT18), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT18), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n434), .A2(new_n435), .A3(new_n438), .A4(new_n441), .ZN(new_n442));
  AND2_X1   g0242(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n352), .A2(new_n386), .A3(new_n430), .A4(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n321), .B1(new_n313), .B2(new_n315), .ZN(new_n445));
  AOI21_X1  g0245(.A(KEYINPUT72), .B1(new_n445), .B2(new_n351), .ZN(new_n446));
  OAI21_X1  g0246(.A(KEYINPUT76), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n445), .A2(new_n351), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT72), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n370), .A2(new_n379), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n384), .A2(new_n385), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n440), .A2(new_n426), .A3(new_n429), .A4(new_n442), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT76), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n450), .A2(new_n455), .A3(new_n456), .A4(new_n352), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n447), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n207), .A2(G45), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n258), .A2(G250), .A3(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n460), .B1(new_n261), .B2(new_n459), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n247), .A2(G244), .A3(G1698), .ZN(new_n462));
  NAND2_X1  g0262(.A1(G33), .A2(G116), .ZN(new_n463));
  INV_X1    g0263(.A(G238), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n462), .B(new_n463), .C1(new_n464), .C2(new_n255), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n461), .B1(new_n465), .B2(new_n259), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n342), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n467), .B1(G200), .B2(new_n466), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n207), .A2(G33), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n324), .A2(new_n304), .A3(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n470), .A2(new_n405), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT81), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT19), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n208), .B1(new_n354), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(G87), .A2(G97), .ZN(new_n476));
  AND3_X1   g0276(.A1(new_n476), .A2(KEYINPUT79), .A3(new_n337), .ZN(new_n477));
  AOI21_X1  g0277(.A(KEYINPUT79), .B1(new_n476), .B2(new_n337), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(KEYINPUT80), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT80), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n481), .B(new_n475), .C1(new_n477), .C2(new_n478), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n208), .B(G68), .C1(new_n253), .C2(new_n254), .ZN(new_n483));
  INV_X1    g0283(.A(G97), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n474), .B1(new_n291), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n480), .A2(new_n482), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n279), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n324), .A2(new_n327), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n473), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  AOI211_X1 g0292(.A(KEYINPUT81), .B(new_n490), .C1(new_n488), .C2(new_n279), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n468), .B(new_n472), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n489), .A2(new_n473), .A3(new_n491), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n486), .B1(new_n479), .B2(KEYINPUT80), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n304), .B1(new_n496), .B2(new_n482), .ZN(new_n497));
  OAI21_X1  g0297(.A(KEYINPUT81), .B1(new_n497), .B2(new_n490), .ZN(new_n498));
  INV_X1    g0298(.A(new_n470), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n495), .A2(new_n498), .B1(new_n327), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n466), .A2(G169), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n501), .B1(new_n319), .B2(new_n466), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n494), .B1(new_n500), .B2(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(KEYINPUT5), .B1(new_n412), .B2(new_n264), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT5), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n207), .B(G45), .C1(new_n506), .C2(G41), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n217), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n261), .B1(new_n509), .B2(new_n257), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n508), .A2(KEYINPUT78), .A3(new_n510), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n506), .B1(new_n265), .B2(new_n266), .ZN(new_n512));
  INV_X1    g0312(.A(new_n507), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n512), .A2(new_n510), .A3(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT78), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n259), .B1(new_n512), .B2(new_n513), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n511), .A2(new_n516), .B1(G257), .B2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT77), .ZN(new_n519));
  INV_X1    g0319(.A(G244), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n519), .B1(new_n255), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(KEYINPUT4), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT4), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n519), .B(new_n523), .C1(new_n255), .C2(new_n520), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n247), .A2(G250), .A3(G1698), .ZN(new_n525));
  NAND2_X1  g0325(.A1(G33), .A2(G283), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  AND3_X1   g0328(.A1(new_n522), .A2(new_n524), .A3(new_n528), .ZN(new_n529));
  OAI211_X1 g0329(.A(G190), .B(new_n518), .C1(new_n529), .C2(new_n258), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n337), .A2(KEYINPUT6), .A3(G97), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n484), .A2(new_n337), .ZN(new_n532));
  NOR2_X1   g0332(.A1(G97), .A2(G107), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n531), .B1(new_n534), .B2(KEYINPUT6), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n535), .A2(G20), .B1(G77), .B2(new_n299), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n387), .A2(new_n390), .A3(G107), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n304), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n283), .A2(new_n484), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n539), .B1(new_n470), .B2(new_n484), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n527), .B1(KEYINPUT4), .B2(new_n521), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n258), .B1(new_n542), .B2(new_n524), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n511), .A2(new_n516), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n517), .A2(G257), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n530), .B(new_n541), .C1(new_n547), .C2(new_n274), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n349), .B1(new_n543), .B2(new_n546), .ZN(new_n549));
  OR2_X1    g0349(.A1(new_n538), .A2(new_n540), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n319), .B(new_n518), .C1(new_n529), .C2(new_n258), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n504), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(KEYINPUT25), .B1(new_n283), .B2(new_n337), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n283), .A2(KEYINPUT25), .A3(new_n337), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n499), .A2(G107), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT24), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n208), .B(G87), .C1(new_n253), .C2(new_n254), .ZN(new_n561));
  XNOR2_X1  g0361(.A(new_n561), .B(KEYINPUT22), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n463), .A2(G20), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT23), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n564), .B1(new_n208), .B2(G107), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n337), .A2(KEYINPUT23), .A3(G20), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n563), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n560), .B1(new_n562), .B2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n562), .A2(new_n560), .A3(new_n567), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n559), .B1(new_n571), .B2(new_n279), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n247), .A2(G257), .A3(G1698), .ZN(new_n573));
  NAND2_X1  g0373(.A1(G33), .A2(G294), .ZN(new_n574));
  INV_X1    g0374(.A(G250), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n573), .B(new_n574), .C1(new_n255), .C2(new_n575), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n576), .A2(new_n259), .B1(new_n517), .B2(G264), .ZN(new_n577));
  AOI21_X1  g0377(.A(G200), .B1(new_n577), .B2(new_n544), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT85), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n577), .A2(new_n544), .ZN(new_n580));
  OAI22_X1  g0380(.A1(new_n578), .A2(new_n579), .B1(new_n580), .B2(G190), .ZN(new_n581));
  AND2_X1   g0381(.A1(new_n578), .A2(new_n579), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n572), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  AND3_X1   g0383(.A1(new_n577), .A2(G179), .A3(new_n544), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n349), .B1(new_n577), .B2(new_n544), .ZN(new_n585));
  OAI21_X1  g0385(.A(KEYINPUT84), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n580), .A2(G169), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT84), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n577), .A2(G179), .A3(new_n544), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(new_n570), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n279), .B1(new_n591), .B2(new_n568), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n558), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n586), .A2(new_n590), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n583), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n247), .A2(G264), .A3(G1698), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n388), .A2(G303), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT83), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n335), .A2(new_n599), .A3(new_n247), .A4(G257), .ZN(new_n600));
  INV_X1    g0400(.A(G257), .ZN(new_n601));
  OAI21_X1  g0401(.A(KEYINPUT83), .B1(new_n255), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n598), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  OR2_X1    g0403(.A1(new_n603), .A2(new_n258), .ZN(new_n604));
  OAI211_X1 g0404(.A(G270), .B(new_n258), .C1(new_n505), .C2(new_n507), .ZN(new_n605));
  XNOR2_X1  g0405(.A(new_n605), .B(KEYINPUT82), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n604), .A2(G190), .A3(new_n606), .A4(new_n544), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n544), .B1(new_n603), .B2(new_n258), .ZN(new_n608));
  XOR2_X1   g0408(.A(new_n605), .B(KEYINPUT82), .Z(new_n609));
  OAI21_X1  g0409(.A(G200), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n324), .A2(G116), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n611), .B1(new_n499), .B2(G116), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n526), .B(new_n208), .C1(G33), .C2(new_n484), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n613), .B(new_n279), .C1(new_n208), .C2(G116), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT20), .ZN(new_n615));
  XNOR2_X1  g0415(.A(new_n614), .B(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n607), .A2(new_n610), .A3(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n349), .B1(new_n612), .B2(new_n616), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n620), .B1(new_n608), .B2(new_n609), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT21), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n608), .A2(new_n609), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n624), .A2(G179), .A3(new_n617), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n620), .B(KEYINPUT21), .C1(new_n608), .C2(new_n609), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n619), .A2(new_n623), .A3(new_n625), .A4(new_n626), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n595), .A2(new_n627), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n458), .A2(new_n554), .A3(new_n628), .ZN(G372));
  NAND2_X1  g0429(.A1(new_n499), .A2(new_n327), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n630), .B1(new_n492), .B2(new_n493), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n502), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n553), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n471), .B1(new_n495), .B2(new_n498), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n631), .A2(new_n502), .B1(new_n635), .B2(new_n468), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n634), .A2(new_n636), .A3(new_n583), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n587), .A2(new_n589), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n593), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n639), .A2(new_n623), .A3(new_n626), .A4(new_n625), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n633), .B1(new_n637), .B2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n552), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n632), .A2(new_n642), .A3(KEYINPUT26), .A4(new_n494), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(KEYINPUT86), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT86), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n636), .A2(new_n645), .A3(KEYINPUT26), .A4(new_n642), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT26), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n647), .B1(new_n504), .B2(new_n552), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n644), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n641), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n458), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n436), .A2(new_n437), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n435), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(KEYINPUT18), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n435), .A2(new_n441), .A3(new_n652), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n350), .A2(new_n348), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n452), .A2(new_n659), .B1(new_n370), .B2(new_n379), .ZN(new_n660));
  INV_X1    g0460(.A(new_n430), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n657), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n321), .B1(new_n662), .B2(new_n316), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n651), .A2(new_n663), .ZN(G369));
  INV_X1    g0464(.A(new_n595), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(G213), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g0469(.A(new_n669), .B(KEYINPUT87), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(G343), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n665), .B1(new_n572), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n594), .B2(new_n671), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n623), .A2(new_n625), .A3(new_n626), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n618), .A2(new_n671), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n676), .B1(new_n627), .B2(new_n675), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(G330), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n673), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g0480(.A(new_n680), .B(KEYINPUT88), .Z(new_n681));
  AND2_X1   g0481(.A1(new_n674), .A2(new_n671), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(new_n665), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n593), .A2(new_n638), .A3(new_n671), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n681), .A2(new_n685), .ZN(G399));
  INV_X1    g0486(.A(new_n211), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n412), .A2(new_n264), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n477), .A2(new_n478), .ZN(new_n690));
  INV_X1    g0490(.A(G116), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NOR3_X1   g0492(.A1(new_n689), .A2(new_n207), .A3(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT89), .ZN(new_n694));
  AOI22_X1  g0494(.A1(new_n693), .A2(new_n694), .B1(new_n216), .B2(new_n689), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n695), .B1(new_n694), .B2(new_n693), .ZN(new_n696));
  XNOR2_X1  g0496(.A(new_n696), .B(KEYINPUT28), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT29), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n650), .A2(new_n698), .A3(new_n671), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n648), .A2(new_n643), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n594), .A2(new_n623), .A3(new_n626), .A4(new_n625), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n554), .A2(new_n583), .A3(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n700), .A2(new_n702), .A3(new_n632), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n671), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(KEYINPUT29), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n699), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT30), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n624), .A2(new_n547), .A3(G179), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n577), .A2(new_n466), .A3(KEYINPUT90), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(KEYINPUT90), .B1(new_n577), .B2(new_n466), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n707), .B1(new_n708), .B2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n711), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(new_n709), .ZN(new_n715));
  NOR3_X1   g0515(.A1(new_n608), .A2(new_n609), .A3(new_n319), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n715), .A2(new_n716), .A3(KEYINPUT30), .A4(new_n547), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n466), .A2(G179), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(new_n580), .ZN(new_n719));
  OR3_X1    g0519(.A1(new_n624), .A2(new_n547), .A3(new_n719), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n713), .A2(new_n717), .A3(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n671), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT31), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n628), .A2(new_n554), .A3(new_n671), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n721), .A2(KEYINPUT31), .A3(new_n722), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(G330), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n706), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n697), .B1(new_n731), .B2(G1), .ZN(G364));
  NOR2_X1   g0532(.A1(new_n282), .A2(G20), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n207), .B1(new_n733), .B2(G45), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n689), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n679), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n737), .B1(G330), .B2(new_n677), .ZN(new_n738));
  INV_X1    g0538(.A(new_n736), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n217), .B1(G20), .B2(new_n349), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n319), .A2(new_n274), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n208), .A2(G190), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(G317), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(KEYINPUT33), .ZN(new_n747));
  OR2_X1    g0547(.A1(new_n746), .A2(KEYINPUT33), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n745), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(G303), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n208), .A2(new_n342), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n751), .A2(new_n319), .A3(G200), .ZN(new_n752));
  INV_X1    g0552(.A(G322), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n319), .A2(G200), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  OAI221_X1 g0555(.A(new_n749), .B1(new_n750), .B2(new_n752), .C1(new_n753), .C2(new_n755), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n743), .A2(new_n319), .A3(G200), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT91), .ZN(new_n758));
  OR2_X1    g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n757), .A2(new_n758), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n756), .B1(G283), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G179), .A2(G200), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G190), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G20), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G294), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n751), .A2(new_n742), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n247), .B1(new_n769), .B2(G326), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n743), .A2(new_n754), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n743), .A2(new_n764), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  AOI22_X1  g0574(.A1(G311), .A2(new_n772), .B1(new_n774), .B2(G329), .ZN(new_n775));
  NAND4_X1  g0575(.A1(new_n763), .A2(new_n767), .A3(new_n770), .A4(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n766), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(new_n484), .ZN(new_n778));
  INV_X1    g0578(.A(new_n755), .ZN(new_n779));
  AOI211_X1 g0579(.A(new_n388), .B(new_n778), .C1(G58), .C2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(G159), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n773), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g0582(.A(new_n782), .B(KEYINPUT32), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n762), .A2(G107), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n752), .A2(new_n405), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n768), .A2(new_n201), .B1(new_n771), .B2(new_n249), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n785), .B(new_n786), .C1(G68), .C2(new_n745), .ZN(new_n787));
  NAND4_X1  g0587(.A1(new_n780), .A2(new_n783), .A3(new_n784), .A4(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n741), .B1(new_n776), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(G13), .A2(G33), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(G20), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n740), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n687), .A2(new_n388), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n794), .A2(G355), .B1(new_n691), .B2(new_n687), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n687), .A2(new_n247), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(G45), .B2(new_n215), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n245), .A2(new_n268), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n795), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n739), .B(new_n789), .C1(new_n793), .C2(new_n799), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n800), .B(KEYINPUT92), .ZN(new_n801));
  INV_X1    g0601(.A(new_n792), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n801), .B1(new_n677), .B2(new_n802), .ZN(new_n803));
  AND2_X1   g0603(.A1(new_n738), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(G396));
  NOR2_X1   g0605(.A1(new_n740), .A2(new_n790), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n739), .B1(new_n249), .B2(new_n806), .ZN(new_n807));
  AOI22_X1  g0607(.A1(G143), .A2(new_n779), .B1(new_n772), .B2(G159), .ZN(new_n808));
  INV_X1    g0608(.A(G137), .ZN(new_n809));
  INV_X1    g0609(.A(G150), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n808), .B1(new_n809), .B2(new_n768), .C1(new_n810), .C2(new_n744), .ZN(new_n811));
  XOR2_X1   g0611(.A(KEYINPUT93), .B(KEYINPUT34), .Z(new_n812));
  XNOR2_X1  g0612(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n762), .A2(G68), .ZN(new_n814));
  INV_X1    g0614(.A(G132), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n247), .B1(new_n773), .B2(new_n815), .C1(new_n752), .C2(new_n201), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n816), .B1(G58), .B2(new_n766), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n813), .A2(new_n814), .A3(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(G311), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n768), .A2(new_n750), .B1(new_n773), .B2(new_n819), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n247), .B(new_n820), .C1(G116), .C2(new_n772), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n762), .A2(G87), .ZN(new_n822));
  INV_X1    g0622(.A(new_n778), .ZN(new_n823));
  INV_X1    g0623(.A(G294), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n752), .A2(new_n337), .B1(new_n755), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(G283), .B2(new_n745), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n821), .A2(new_n822), .A3(new_n823), .A4(new_n826), .ZN(new_n827));
  AND2_X1   g0627(.A1(new_n818), .A2(new_n827), .ZN(new_n828));
  AND2_X1   g0628(.A1(new_n344), .A2(new_n347), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n671), .A2(new_n330), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n658), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n659), .A2(new_n671), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n807), .B1(new_n741), .B2(new_n828), .C1(new_n834), .C2(new_n791), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n834), .B1(new_n650), .B2(new_n671), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n722), .B(new_n833), .C1(new_n641), .C2(new_n649), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n736), .B1(new_n838), .B2(new_n730), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n729), .B1(new_n836), .B2(new_n837), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT94), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n839), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AND2_X1   g0642(.A1(new_n840), .A2(new_n841), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n835), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n844), .B(KEYINPUT95), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(G384));
  OR2_X1    g0646(.A1(new_n535), .A2(KEYINPUT35), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n535), .A2(KEYINPUT35), .ZN(new_n848));
  NAND4_X1  g0648(.A1(new_n847), .A2(G116), .A3(new_n218), .A4(new_n848), .ZN(new_n849));
  XNOR2_X1  g0649(.A(KEYINPUT96), .B(KEYINPUT36), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n849), .B(new_n850), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n216), .B(G77), .C1(new_n202), .C2(new_n203), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n207), .B(G13), .C1(new_n852), .C2(new_n241), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n451), .A2(new_n722), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT100), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n391), .A2(new_n394), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(KEYINPUT16), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n391), .A2(new_n392), .A3(new_n394), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n304), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n401), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n670), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n862), .B(KEYINPUT97), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n454), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(KEYINPUT98), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT98), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n454), .A2(new_n866), .A3(new_n863), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n653), .A2(new_n424), .ZN(new_n869));
  OAI21_X1  g0669(.A(KEYINPUT37), .B1(new_n863), .B2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT37), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n439), .A2(new_n871), .A3(new_n424), .A4(new_n862), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(KEYINPUT38), .B1(new_n868), .B2(new_n873), .ZN(new_n874));
  AND3_X1   g0674(.A1(new_n454), .A2(new_n866), .A3(new_n863), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n866), .B1(new_n454), .B2(new_n863), .ZN(new_n876));
  OAI211_X1 g0676(.A(KEYINPUT38), .B(new_n873), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n856), .B(KEYINPUT39), .C1(new_n874), .C2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n653), .A2(new_n424), .A3(new_n862), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(KEYINPUT37), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n872), .ZN(new_n882));
  INV_X1    g0682(.A(new_n862), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n654), .A2(new_n426), .A3(new_n429), .A4(new_n655), .ZN(new_n884));
  AOI22_X1  g0684(.A1(new_n882), .A2(KEYINPUT101), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT101), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n881), .A2(new_n872), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(KEYINPUT38), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n865), .A2(new_n867), .B1(new_n870), .B2(new_n872), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n888), .B1(new_n889), .B2(KEYINPUT38), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT39), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n879), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n873), .B1(new_n875), .B2(new_n876), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT38), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n877), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n856), .B1(new_n897), .B2(KEYINPUT39), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n855), .B1(new_n893), .B2(new_n898), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n722), .A2(new_n379), .ZN(new_n900));
  OR2_X1    g0700(.A1(new_n453), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n370), .A2(new_n900), .ZN(new_n902));
  AND2_X1   g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AND3_X1   g0703(.A1(new_n644), .A2(new_n646), .A3(new_n648), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n554), .A2(new_n583), .A3(new_n640), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n632), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n671), .B(new_n834), .C1(new_n904), .C2(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n903), .B1(new_n907), .B2(new_n832), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n897), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n657), .A2(new_n670), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(KEYINPUT99), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT99), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n909), .A2(new_n914), .A3(new_n911), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n899), .A2(new_n913), .A3(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n663), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT102), .B1(new_n706), .B2(new_n458), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  AOI211_X1 g0719(.A(KEYINPUT29), .B(new_n722), .C1(new_n641), .C2(new_n649), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n698), .B1(new_n703), .B2(new_n671), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n458), .B(KEYINPUT102), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n917), .B1(new_n919), .B2(new_n922), .ZN(new_n923));
  XOR2_X1   g0723(.A(new_n916), .B(new_n923), .Z(new_n924));
  NAND2_X1  g0724(.A1(new_n728), .A2(KEYINPUT103), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n833), .B1(new_n901), .B2(new_n902), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT103), .ZN(new_n927));
  NAND4_X1  g0727(.A1(new_n725), .A2(new_n726), .A3(new_n927), .A4(new_n727), .ZN(new_n928));
  AND3_X1   g0728(.A1(new_n925), .A2(new_n926), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(KEYINPUT40), .B1(new_n896), .B2(new_n877), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n925), .A2(new_n926), .A3(new_n928), .ZN(new_n933));
  OAI21_X1  g0733(.A(KEYINPUT40), .B1(new_n933), .B2(new_n890), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n932), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n458), .A2(new_n925), .A3(new_n928), .ZN(new_n937));
  OR2_X1    g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n936), .A2(new_n937), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n938), .A2(G330), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n924), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n207), .B2(new_n733), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n924), .A2(new_n940), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n854), .B1(new_n942), .B2(new_n943), .ZN(G367));
  OAI21_X1  g0744(.A(new_n793), .B1(new_n211), .B2(new_n328), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(new_n796), .B2(new_n231), .ZN(new_n946));
  INV_X1    g0746(.A(new_n752), .ZN(new_n947));
  AOI22_X1  g0747(.A1(new_n947), .A2(G58), .B1(new_n745), .B2(G159), .ZN(new_n948));
  OAI221_X1 g0748(.A(new_n948), .B1(new_n201), .B2(new_n771), .C1(new_n761), .C2(new_n249), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n777), .A2(new_n203), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n247), .B1(new_n755), .B2(new_n810), .ZN(new_n951));
  INV_X1    g0751(.A(G143), .ZN(new_n952));
  OAI22_X1  g0752(.A1(new_n768), .A2(new_n952), .B1(new_n773), .B2(new_n809), .ZN(new_n953));
  NOR4_X1   g0753(.A1(new_n949), .A2(new_n950), .A3(new_n951), .A4(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT108), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n752), .B2(new_n691), .ZN(new_n956));
  AOI22_X1  g0756(.A1(new_n956), .A2(KEYINPUT46), .B1(G294), .B2(new_n745), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(KEYINPUT46), .B2(new_n956), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n958), .B(KEYINPUT109), .Z(new_n959));
  OAI221_X1 g0759(.A(new_n388), .B1(new_n755), .B2(new_n750), .C1(new_n777), .C2(new_n337), .ZN(new_n960));
  AOI22_X1  g0760(.A1(G283), .A2(new_n772), .B1(new_n774), .B2(G317), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n819), .B2(new_n768), .ZN(new_n962));
  AOI211_X1 g0762(.A(new_n960), .B(new_n962), .C1(G97), .C2(new_n762), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n954), .B1(new_n959), .B2(new_n963), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT47), .Z(new_n965));
  AOI211_X1 g0765(.A(new_n739), .B(new_n946), .C1(new_n965), .C2(new_n740), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n635), .A2(new_n671), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n633), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n504), .B2(new_n967), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n966), .B1(new_n969), .B2(new_n802), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n634), .B1(new_n541), .B2(new_n671), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n642), .A2(new_n722), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(new_n685), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT44), .Z(new_n976));
  NOR2_X1   g0776(.A1(new_n974), .A2(new_n685), .ZN(new_n977));
  XNOR2_X1  g0777(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n977), .B(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n976), .A2(new_n979), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(new_n681), .Z(new_n981));
  OAI21_X1  g0781(.A(new_n683), .B1(new_n673), .B2(new_n682), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(new_n679), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n730), .B(new_n706), .C1(new_n981), .C2(new_n983), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n689), .B(KEYINPUT41), .Z(new_n985));
  OAI21_X1  g0785(.A(new_n734), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT107), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n974), .A2(new_n683), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT42), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n552), .B1(new_n971), .B2(new_n594), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n671), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n969), .A2(KEYINPUT43), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT105), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n681), .A2(new_n973), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n995), .B(new_n996), .ZN(new_n997));
  XOR2_X1   g0797(.A(KEYINPUT104), .B(KEYINPUT43), .Z(new_n998));
  OR2_X1    g0798(.A1(new_n969), .A2(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n997), .B(new_n999), .ZN(new_n1000));
  AND3_X1   g0800(.A1(new_n986), .A2(new_n987), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n987), .B1(new_n986), .B2(new_n1000), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n970), .B1(new_n1001), .B2(new_n1002), .ZN(G387));
  OR2_X1    g0803(.A1(new_n673), .A2(new_n802), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n796), .B1(new_n236), .B2(new_n268), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n692), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n794), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1005), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n268), .B1(new_n203), .B2(new_n249), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n290), .A2(new_n201), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1009), .B1(new_n1010), .B2(KEYINPUT50), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n1006), .B(new_n1011), .C1(KEYINPUT50), .C2(new_n1010), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n1008), .A2(new_n1012), .B1(new_n337), .B2(new_n687), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n793), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n736), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n947), .A2(G77), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n289), .B2(new_n744), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n388), .B(new_n1017), .C1(G150), .C2(new_n774), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n762), .A2(G97), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n766), .A2(new_n327), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n755), .A2(new_n201), .B1(new_n771), .B2(new_n203), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(G159), .B2(new_n769), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .A4(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(G283), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n777), .A2(new_n1024), .B1(new_n752), .B2(new_n824), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n768), .A2(new_n753), .B1(new_n744), .B2(new_n819), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n755), .A2(new_n746), .B1(new_n771), .B2(new_n750), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1025), .B1(new_n1028), .B2(KEYINPUT48), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(KEYINPUT48), .B2(new_n1028), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(KEYINPUT110), .B(KEYINPUT49), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1030), .B(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n247), .B1(new_n774), .B2(G326), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n761), .B2(new_n691), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1023), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  OR2_X1    g0835(.A1(new_n1035), .A2(KEYINPUT111), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n741), .B1(new_n1035), .B2(KEYINPUT111), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1015), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n983), .A2(new_n735), .B1(new_n1004), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n731), .A2(new_n983), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n689), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n731), .A2(new_n983), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1039), .B1(new_n1041), .B2(new_n1042), .ZN(G393));
  NAND2_X1  g0843(.A1(new_n974), .A2(new_n792), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n796), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n793), .B1(new_n484), .B2(new_n211), .C1(new_n1045), .C2(new_n240), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(new_n736), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n744), .A2(new_n750), .B1(new_n773), .B2(new_n753), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n388), .B1(new_n771), .B2(new_n824), .C1(new_n777), .C2(new_n691), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n1048), .B(new_n1049), .C1(G283), .C2(new_n947), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n768), .A2(new_n746), .B1(new_n755), .B2(new_n819), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT52), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1050), .A2(new_n784), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n1055), .A2(KEYINPUT112), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(KEYINPUT112), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n771), .A2(new_n289), .B1(new_n773), .B2(new_n952), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n766), .A2(G77), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1059), .B(new_n247), .C1(new_n201), .C2(new_n744), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n1058), .B(new_n1060), .C1(G68), .C2(new_n947), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n768), .A2(new_n810), .B1(new_n755), .B2(new_n781), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT51), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1061), .A2(new_n822), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1056), .A2(new_n1057), .A3(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1047), .B1(new_n1067), .B2(new_n740), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n981), .A2(new_n735), .B1(new_n1044), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n981), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n689), .B1(new_n1070), .B2(new_n1040), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n981), .B1(new_n731), .B2(new_n983), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1069), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT113), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(G390));
  NAND2_X1  g0875(.A1(new_n907), .A2(new_n832), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n903), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n855), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n891), .B1(new_n896), .B2(new_n877), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n1080), .A2(new_n856), .B1(new_n891), .B2(new_n890), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n897), .A2(KEYINPUT39), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(KEYINPUT100), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1079), .A2(new_n1081), .A3(new_n1083), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n728), .A2(G330), .A3(new_n834), .ZN(new_n1085));
  OR2_X1    g0885(.A1(new_n1085), .A2(new_n903), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n855), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n703), .A2(new_n671), .A3(new_n831), .ZN(new_n1088));
  AND2_X1   g0888(.A1(new_n1088), .A2(new_n832), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n1087), .B1(new_n878), .B2(new_n888), .C1(new_n1089), .C2(new_n903), .ZN(new_n1090));
  AND3_X1   g0890(.A1(new_n1084), .A2(new_n1086), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(G330), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n933), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(new_n1084), .B2(new_n1090), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n1091), .A2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n458), .A2(G330), .A3(new_n925), .A4(new_n928), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n922), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n663), .B(new_n1097), .C1(new_n1098), .C2(new_n918), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n925), .A2(G330), .A3(new_n928), .ZN(new_n1100));
  AND2_X1   g0900(.A1(new_n1100), .A2(KEYINPUT114), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT114), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n925), .A2(new_n1102), .A3(G330), .A4(new_n928), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n834), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n903), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1105));
  AND2_X1   g0905(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1085), .A2(new_n903), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1094), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n1076), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1099), .B1(new_n1107), .B2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(KEYINPUT115), .B1(new_n1096), .B2(new_n1111), .ZN(new_n1112));
  NOR3_X1   g0912(.A1(new_n893), .A2(new_n898), .A3(new_n1078), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1090), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1093), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1084), .A2(new_n1086), .A3(new_n1090), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT115), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1107), .A2(new_n1110), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1117), .B(new_n1118), .C1(new_n1120), .C2(new_n1099), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1096), .A2(new_n1111), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1112), .A2(new_n689), .A3(new_n1121), .A4(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1115), .A2(new_n735), .A3(new_n1116), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT116), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1115), .A2(KEYINPUT116), .A3(new_n1116), .A4(new_n735), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1129), .A2(new_n791), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(G107), .A2(new_n745), .B1(new_n772), .B2(G97), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n814), .B(new_n1131), .C1(new_n691), .C2(new_n755), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n785), .A2(new_n247), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n769), .A2(G283), .B1(new_n774), .B2(G294), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1133), .A2(new_n1134), .A3(new_n1059), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n752), .A2(new_n810), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n1136), .B(KEYINPUT53), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(KEYINPUT54), .B(G143), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT117), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(new_n772), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1137), .B(new_n1140), .C1(new_n201), .C2(new_n761), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n769), .A2(G128), .B1(new_n774), .B2(G125), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n388), .B1(new_n745), .B2(G137), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n779), .A2(G132), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n766), .A2(G159), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1142), .A2(new_n1143), .A3(new_n1144), .A4(new_n1145), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n1132), .A2(new_n1135), .B1(new_n1141), .B2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n741), .B1(new_n1147), .B2(KEYINPUT118), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1148), .B1(KEYINPUT118), .B2(new_n1147), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n806), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1149), .B(new_n736), .C1(new_n290), .C2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1130), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(KEYINPUT119), .B1(new_n1128), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT119), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n1155), .B(new_n1152), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1123), .B1(new_n1154), .B2(new_n1156), .ZN(G378));
  INV_X1    g0957(.A(new_n1099), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n1117), .B2(new_n1120), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n670), .B1(new_n303), .B2(new_n307), .ZN(new_n1160));
  XOR2_X1   g0960(.A(new_n1160), .B(KEYINPUT55), .Z(new_n1161));
  XNOR2_X1  g0961(.A(new_n445), .B(new_n1161), .ZN(new_n1162));
  XOR2_X1   g0962(.A(KEYINPUT122), .B(KEYINPUT56), .Z(new_n1163));
  XOR2_X1   g0963(.A(new_n1162), .B(new_n1163), .Z(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1092), .B1(new_n931), .B2(new_n934), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  AOI211_X1 g0967(.A(KEYINPUT99), .B(new_n910), .C1(new_n908), .C2(new_n897), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(new_n1129), .B2(new_n855), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1167), .B1(new_n1169), .B2(new_n913), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1087), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n914), .B1(new_n909), .B2(new_n911), .ZN(new_n1172));
  NOR4_X1   g0972(.A1(new_n1171), .A2(new_n1166), .A3(new_n1172), .A4(new_n1168), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1165), .B1(new_n1170), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n916), .A2(new_n1166), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1169), .A2(new_n913), .A3(new_n1167), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1175), .A2(new_n1176), .A3(new_n1164), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1159), .A2(new_n1174), .A3(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT57), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1159), .A2(new_n1174), .A3(KEYINPUT57), .A4(new_n1177), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1180), .A2(new_n689), .A3(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n736), .B1(G50), .B2(new_n1150), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n745), .A2(G97), .B1(new_n774), .B2(G283), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n1184), .B1(new_n337), .B2(new_n755), .C1(new_n761), .C2(new_n202), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n769), .A2(G116), .B1(new_n772), .B2(new_n327), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n688), .A2(new_n247), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1186), .A2(new_n1016), .A3(new_n1187), .ZN(new_n1188));
  NOR3_X1   g0988(.A1(new_n1185), .A2(new_n950), .A3(new_n1188), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1187), .ZN(new_n1191));
  AOI21_X1  g0991(.A(G50), .B1(new_n293), .B2(new_n411), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n1189), .A2(new_n1190), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(G125), .A2(new_n769), .B1(new_n779), .B2(G128), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(G132), .A2(new_n745), .B1(new_n772), .B2(G137), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n766), .A2(G150), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1194), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(new_n947), .B2(new_n1139), .ZN(new_n1198));
  XOR2_X1   g0998(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n1199));
  XNOR2_X1  g0999(.A(new_n1198), .B(new_n1199), .ZN(new_n1200));
  AOI211_X1 g1000(.A(G33), .B(G41), .C1(new_n774), .C2(G124), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(new_n761), .B2(new_n781), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1193), .B1(new_n1190), .B2(new_n1189), .C1(new_n1200), .C2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1183), .B1(new_n1203), .B2(new_n740), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n1164), .B2(new_n791), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  AND3_X1   g1006(.A1(new_n1175), .A2(new_n1176), .A3(new_n1164), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1164), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1206), .B1(new_n1209), .B2(new_n735), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1182), .A2(new_n1210), .ZN(G375));
  NAND2_X1  g1011(.A1(new_n903), .A2(new_n790), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n736), .B1(G68), .B2(new_n1150), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1213), .B(KEYINPUT123), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n947), .A2(G97), .B1(new_n779), .B2(G283), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n824), .B2(new_n768), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(G77), .B2(new_n762), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n388), .B1(new_n773), .B2(new_n750), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n744), .A2(new_n691), .B1(new_n771), .B2(new_n337), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n1219), .B(new_n1220), .C1(new_n327), .C2(new_n766), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n388), .B1(new_n774), .B2(G128), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n201), .B2(new_n777), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n768), .A2(new_n815), .B1(new_n771), .B2(new_n810), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n752), .A2(new_n781), .B1(new_n755), .B2(new_n809), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(new_n1223), .A2(new_n1224), .A3(new_n1225), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n762), .A2(G58), .B1(new_n1139), .B2(new_n745), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n1218), .A2(new_n1221), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1215), .B1(new_n1229), .B2(new_n740), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n1119), .A2(new_n735), .B1(new_n1212), .B2(new_n1230), .ZN(new_n1231));
  OR2_X1    g1031(.A1(new_n1111), .A2(new_n985), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1119), .A2(new_n1158), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1231), .B1(new_n1232), .B2(new_n1233), .ZN(G381));
  OR4_X1    g1034(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1152), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1236));
  AND2_X1   g1036(.A1(new_n1123), .A2(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1182), .A2(new_n1237), .A3(new_n1210), .ZN(new_n1238));
  OR4_X1    g1038(.A1(G387), .A2(new_n1235), .A3(G381), .A4(new_n1238), .ZN(G407));
  OAI211_X1 g1039(.A(G407), .B(G213), .C1(G343), .C2(new_n1238), .ZN(G409));
  INV_X1    g1040(.A(KEYINPUT61), .ZN(new_n1241));
  INV_X1    g1041(.A(G213), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1242), .A2(G343), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(G378), .A2(new_n1182), .A3(new_n1210), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT124), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1245), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1174), .A2(KEYINPUT124), .A3(new_n1177), .ZN(new_n1247));
  AND3_X1   g1047(.A1(new_n1246), .A2(new_n735), .A3(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1205), .B1(new_n1178), .B2(new_n985), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1237), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1243), .B1(new_n1244), .B2(new_n1250), .ZN(new_n1251));
  OAI21_X1  g1051(.A(KEYINPUT60), .B1(new_n1120), .B2(new_n1099), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1233), .ZN(new_n1253));
  AND2_X1   g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1107), .A2(new_n1110), .A3(new_n1099), .A4(KEYINPUT60), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n689), .ZN(new_n1256));
  OAI211_X1 g1056(.A(G384), .B(new_n1231), .C1(new_n1254), .C2(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1256), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1231), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n845), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1243), .A2(KEYINPUT125), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1257), .A2(new_n1260), .A3(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1243), .A2(G2897), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1262), .A2(new_n1264), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1257), .A2(new_n1260), .A3(new_n1261), .A4(new_n1263), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1241), .B1(new_n1251), .B2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT63), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1244), .A2(new_n1250), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1243), .ZN(new_n1271));
  AND2_X1   g1071(.A1(new_n1257), .A2(new_n1260), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1270), .A2(new_n1271), .A3(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1268), .B1(new_n1269), .B2(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1251), .A2(KEYINPUT63), .A3(new_n1272), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(G387), .A2(new_n1074), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(G387), .A2(new_n1074), .ZN(new_n1278));
  XNOR2_X1  g1078(.A(G393), .B(new_n804), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  NOR3_X1   g1080(.A1(new_n1277), .A2(new_n1278), .A3(new_n1280), .ZN(new_n1281));
  OR2_X1    g1081(.A1(G387), .A2(new_n1074), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1279), .B1(new_n1282), .B2(new_n1276), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1281), .A2(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1274), .A2(new_n1275), .A3(new_n1284), .ZN(new_n1285));
  OR2_X1    g1085(.A1(new_n1281), .A2(new_n1283), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT62), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1273), .A2(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1251), .A2(KEYINPUT62), .A3(new_n1272), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1268), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT126), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1286), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1293));
  AND2_X1   g1093(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1294));
  AOI21_X1  g1094(.A(KEYINPUT61), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1289), .ZN(new_n1296));
  AOI21_X1  g1096(.A(KEYINPUT62), .B1(new_n1251), .B2(new_n1272), .ZN(new_n1297));
  OAI211_X1 g1097(.A(new_n1295), .B(new_n1291), .C1(new_n1296), .C2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1285), .B1(new_n1292), .B2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT127), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  OAI211_X1 g1102(.A(KEYINPUT127), .B(new_n1285), .C1(new_n1292), .C2(new_n1299), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(G405));
  NAND2_X1  g1104(.A1(G375), .A2(new_n1237), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n1244), .ZN(new_n1306));
  XOR2_X1   g1106(.A(new_n1306), .B(new_n1272), .Z(new_n1307));
  XNOR2_X1  g1107(.A(new_n1307), .B(new_n1284), .ZN(G402));
endmodule


