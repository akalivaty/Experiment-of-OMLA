//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 1 0 1 0 1 1 1 1 1 1 0 0 0 0 1 0 0 0 0 1 1 1 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:08 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n905,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(G110), .B(G122), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT82), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT84), .B(KEYINPUT8), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G107), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(KEYINPUT76), .A3(G104), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT3), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n192), .A2(G104), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G101), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT3), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n198), .A2(new_n192), .A3(KEYINPUT76), .A4(G104), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n194), .A2(new_n196), .A3(new_n197), .A4(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G104), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n201), .A2(G107), .ZN(new_n202));
  OAI21_X1  g016(.A(G101), .B1(new_n195), .B2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n200), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G119), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G116), .ZN(new_n207));
  OR2_X1    g021(.A1(new_n207), .A2(KEYINPUT5), .ZN(new_n208));
  INV_X1    g022(.A(G116), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G119), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n207), .A2(new_n210), .A3(KEYINPUT5), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n208), .A2(G113), .A3(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT81), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n208), .A2(KEYINPUT81), .A3(new_n211), .A4(G113), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G113), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(KEYINPUT2), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT2), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G113), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(G116), .B(G119), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT68), .ZN(new_n223));
  AND3_X1   g037(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n223), .B1(new_n221), .B2(new_n222), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n205), .B1(new_n216), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n212), .ZN(new_n229));
  NOR3_X1   g043(.A1(new_n226), .A2(new_n229), .A3(new_n204), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n191), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n216), .A2(new_n227), .A3(new_n205), .ZN(new_n232));
  INV_X1    g046(.A(new_n189), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n194), .A2(new_n196), .A3(new_n199), .ZN(new_n234));
  AND2_X1   g048(.A1(KEYINPUT77), .A2(KEYINPUT4), .ZN(new_n235));
  AND3_X1   g049(.A1(new_n234), .A2(G101), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n234), .A2(G101), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n200), .A2(new_n235), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n236), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  OAI22_X1  g053(.A1(new_n224), .A2(new_n225), .B1(new_n222), .B2(new_n221), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  OAI211_X1 g055(.A(new_n232), .B(new_n233), .C1(new_n239), .C2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G146), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G143), .ZN(new_n244));
  INV_X1    g058(.A(G143), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G146), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT1), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n244), .A2(new_n246), .A3(new_n247), .A4(G128), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT65), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g064(.A(G143), .B(G146), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n251), .A2(KEYINPUT65), .A3(new_n247), .A4(G128), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n244), .A2(new_n246), .ZN(new_n254));
  INV_X1    g068(.A(G128), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(KEYINPUT66), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT66), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G128), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n247), .B1(G143), .B2(new_n243), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n254), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT67), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G125), .ZN(new_n264));
  OAI21_X1  g078(.A(KEYINPUT1), .B1(new_n245), .B2(G146), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n265), .A2(new_n256), .A3(new_n258), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(KEYINPUT67), .A3(new_n254), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n253), .A2(new_n263), .A3(new_n264), .A4(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT83), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  AND3_X1   g084(.A1(new_n266), .A2(KEYINPUT67), .A3(new_n254), .ZN(new_n271));
  AOI21_X1  g085(.A(KEYINPUT67), .B1(new_n266), .B2(new_n254), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n273), .A2(KEYINPUT83), .A3(new_n264), .A4(new_n253), .ZN(new_n274));
  INV_X1    g088(.A(G224), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n275), .A2(G953), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(KEYINPUT0), .A2(G128), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  NOR2_X1   g093(.A1(KEYINPUT0), .A2(G128), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n254), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n251), .A2(new_n278), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(G125), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n270), .A2(new_n274), .A3(new_n277), .A4(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT7), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n231), .B(new_n242), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  AND2_X1   g102(.A1(new_n270), .A2(new_n274), .ZN(new_n289));
  AOI22_X1  g103(.A1(new_n289), .A2(new_n285), .B1(KEYINPUT7), .B2(new_n277), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n187), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT85), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n289), .A2(new_n285), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(new_n276), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n286), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n232), .B1(new_n239), .B2(new_n241), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT6), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n297), .A2(new_n298), .A3(new_n189), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n297), .A2(new_n189), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n300), .A2(KEYINPUT6), .A3(new_n242), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n296), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  OAI211_X1 g116(.A(KEYINPUT85), .B(new_n187), .C1(new_n288), .C2(new_n290), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n293), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(G210), .B1(G237), .B2(G902), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n293), .A2(new_n302), .A3(new_n305), .A4(new_n303), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(G214), .B1(G237), .B2(G902), .ZN(new_n310));
  XOR2_X1   g124(.A(new_n310), .B(KEYINPUT80), .Z(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n245), .B1(new_n256), .B2(new_n258), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n255), .A2(G143), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT90), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G134), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT90), .ZN(new_n317));
  INV_X1    g131(.A(new_n314), .ZN(new_n318));
  XNOR2_X1  g132(.A(KEYINPUT66), .B(G128), .ZN(new_n319));
  OAI211_X1 g133(.A(new_n317), .B(new_n318), .C1(new_n319), .C2(new_n245), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n315), .A2(new_n316), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n314), .A2(KEYINPUT13), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n322), .B1(new_n319), .B2(new_n245), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n314), .A2(KEYINPUT13), .ZN(new_n324));
  OAI21_X1  g138(.A(G134), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  XOR2_X1   g139(.A(G116), .B(G122), .Z(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G107), .ZN(new_n327));
  XNOR2_X1  g141(.A(G116), .B(G122), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n192), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n321), .A2(new_n325), .A3(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT91), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n315), .A2(new_n320), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G134), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(new_n321), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n209), .A2(KEYINPUT14), .A3(G122), .ZN(new_n336));
  OAI211_X1 g150(.A(G107), .B(new_n336), .C1(new_n326), .C2(KEYINPUT14), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n329), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n332), .B1(new_n335), .B2(new_n339), .ZN(new_n340));
  AND3_X1   g154(.A1(new_n315), .A2(new_n316), .A3(new_n320), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n316), .B1(new_n315), .B2(new_n320), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n339), .B(new_n332), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n331), .B1(new_n340), .B2(new_n344), .ZN(new_n345));
  XOR2_X1   g159(.A(KEYINPUT9), .B(G234), .Z(new_n346));
  INV_X1    g160(.A(G953), .ZN(new_n347));
  XNOR2_X1  g161(.A(KEYINPUT71), .B(G217), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n345), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT92), .ZN(new_n351));
  INV_X1    g165(.A(new_n331), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n339), .B1(new_n341), .B2(new_n342), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(KEYINPUT91), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n352), .B1(new_n354), .B2(new_n343), .ZN(new_n355));
  INV_X1    g169(.A(new_n349), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n350), .A2(new_n351), .A3(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n355), .A2(KEYINPUT92), .A3(new_n356), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT15), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(G478), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n361), .B(KEYINPUT93), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n358), .A2(new_n187), .A3(new_n359), .A4(new_n362), .ZN(new_n363));
  OR2_X1    g177(.A1(new_n363), .A2(KEYINPUT94), .ZN(new_n364));
  NAND2_X1  g178(.A1(G234), .A2(G237), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n365), .A2(G952), .A3(new_n347), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  XOR2_X1   g181(.A(KEYINPUT21), .B(G898), .Z(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n365), .A2(G902), .A3(G953), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n367), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  NOR3_X1   g186(.A1(new_n264), .A2(KEYINPUT16), .A3(G140), .ZN(new_n373));
  INV_X1    g187(.A(G140), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n264), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(G125), .A2(G140), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n373), .B1(new_n377), .B2(KEYINPUT16), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n378), .A2(G146), .ZN(new_n379));
  AOI211_X1 g193(.A(new_n243), .B(new_n373), .C1(new_n377), .C2(KEYINPUT16), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NOR2_X1   g195(.A1(G237), .A2(G953), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(G143), .A3(G214), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(G143), .B1(new_n382), .B2(G214), .ZN(new_n385));
  OAI211_X1 g199(.A(KEYINPUT17), .B(G131), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(G237), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n387), .A2(new_n347), .A3(G214), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n245), .ZN(new_n389));
  INV_X1    g203(.A(G131), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(new_n390), .A3(new_n383), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(KEYINPUT87), .ZN(new_n392));
  OAI21_X1  g206(.A(G131), .B1(new_n384), .B2(new_n385), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT87), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n389), .A2(new_n394), .A3(new_n390), .A4(new_n383), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n392), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n381), .B(new_n386), .C1(new_n396), .C2(KEYINPUT17), .ZN(new_n397));
  XNOR2_X1  g211(.A(G113), .B(G122), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n398), .B(new_n201), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n384), .A2(new_n385), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT86), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT18), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n400), .B(new_n401), .C1(new_n402), .C2(new_n390), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n377), .B(new_n243), .ZN(new_n404));
  OAI211_X1 g218(.A(KEYINPUT18), .B(G131), .C1(new_n384), .C2(new_n385), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n389), .B(new_n383), .C1(new_n402), .C2(new_n390), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(KEYINPUT86), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n403), .A2(new_n404), .A3(new_n405), .A4(new_n407), .ZN(new_n408));
  AND3_X1   g222(.A1(new_n397), .A2(new_n399), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n399), .B1(new_n397), .B2(new_n408), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n187), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  AND2_X1   g225(.A1(new_n411), .A2(G475), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n378), .A2(G146), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT19), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n377), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n375), .A2(KEYINPUT19), .A3(new_n376), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n415), .A2(new_n243), .A3(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n396), .A2(new_n413), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n408), .ZN(new_n419));
  INV_X1    g233(.A(new_n399), .ZN(new_n420));
  AOI21_X1  g234(.A(KEYINPUT88), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT88), .ZN(new_n422));
  AOI211_X1 g236(.A(new_n422), .B(new_n399), .C1(new_n418), .C2(new_n408), .ZN(new_n423));
  NOR3_X1   g237(.A1(new_n421), .A2(new_n423), .A3(new_n409), .ZN(new_n424));
  NOR2_X1   g238(.A1(G475), .A2(G902), .ZN(new_n425));
  XOR2_X1   g239(.A(new_n425), .B(KEYINPUT89), .Z(new_n426));
  OAI21_X1  g240(.A(KEYINPUT20), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n421), .ZN(new_n428));
  INV_X1    g242(.A(new_n409), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n419), .A2(KEYINPUT88), .A3(new_n420), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT20), .ZN(new_n432));
  INV_X1    g246(.A(new_n426), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n431), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  AOI211_X1 g248(.A(new_n372), .B(new_n412), .C1(new_n427), .C2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n358), .A2(new_n187), .A3(new_n359), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n436), .A2(new_n360), .A3(G478), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n363), .A2(KEYINPUT94), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n364), .A2(new_n435), .A3(new_n437), .A4(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(KEYINPUT95), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT94), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n363), .B(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT95), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n442), .A2(new_n443), .A3(new_n437), .A4(new_n435), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n312), .B1(new_n440), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(G472), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT11), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n447), .B1(new_n316), .B2(G137), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n316), .A2(G137), .ZN(new_n449));
  INV_X1    g263(.A(G137), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n450), .A2(KEYINPUT11), .A3(G134), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n448), .A2(new_n449), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(G131), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n448), .A2(new_n451), .A3(new_n390), .A4(new_n449), .ZN(new_n454));
  AOI22_X1  g268(.A1(new_n453), .A2(new_n454), .B1(new_n281), .B2(new_n282), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n253), .A2(new_n263), .A3(new_n267), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n450), .A2(G134), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n316), .A2(G137), .ZN(new_n458));
  OAI21_X1  g272(.A(G131), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n454), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  AOI211_X1 g275(.A(new_n455), .B(new_n240), .C1(new_n456), .C2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT28), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n455), .B1(new_n456), .B2(new_n461), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n241), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT28), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT64), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n460), .B(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n455), .B1(new_n470), .B2(new_n456), .ZN(new_n471));
  OR2_X1    g285(.A1(new_n471), .A2(new_n241), .ZN(new_n472));
  XNOR2_X1  g286(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n473), .B(G101), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n382), .A2(G210), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n474), .B(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n468), .A2(new_n472), .A3(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT29), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n456), .A2(new_n461), .ZN(new_n479));
  INV_X1    g293(.A(new_n455), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n479), .A2(KEYINPUT30), .A3(new_n480), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n481), .B(new_n240), .C1(new_n471), .C2(KEYINPUT30), .ZN(new_n482));
  AND2_X1   g296(.A1(new_n482), .A2(new_n466), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n477), .B(new_n478), .C1(new_n483), .C2(new_n476), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n465), .A2(new_n241), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n485), .B1(new_n464), .B2(new_n467), .ZN(new_n486));
  INV_X1    g300(.A(new_n476), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n487), .A2(new_n478), .ZN(new_n488));
  AOI21_X1  g302(.A(G902), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n446), .B1(new_n484), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(KEYINPUT69), .B1(new_n462), .B2(new_n487), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT69), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n466), .A2(new_n492), .A3(new_n476), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n491), .A2(new_n482), .A3(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT31), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n491), .A2(new_n482), .A3(KEYINPUT31), .A4(new_n493), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n468), .A2(new_n472), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n487), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT32), .ZN(new_n502));
  NOR2_X1   g316(.A1(G472), .A2(G902), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n503), .B(KEYINPUT70), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n501), .A2(new_n502), .A3(new_n505), .ZN(new_n506));
  AOI22_X1  g320(.A1(new_n496), .A2(new_n497), .B1(new_n499), .B2(new_n487), .ZN(new_n507));
  OAI21_X1  g321(.A(KEYINPUT32), .B1(new_n507), .B2(new_n504), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n490), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n347), .A2(G221), .A3(G234), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n510), .B(KEYINPUT22), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n511), .B(new_n450), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n255), .A2(G119), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n514), .B1(new_n319), .B2(new_n206), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  XOR2_X1   g330(.A(KEYINPUT24), .B(G110), .Z(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n518), .B1(new_n379), .B2(new_n380), .ZN(new_n519));
  AOI21_X1  g333(.A(KEYINPUT23), .B1(new_n255), .B2(G119), .ZN(new_n520));
  AOI211_X1 g334(.A(KEYINPUT72), .B(new_n520), .C1(new_n515), .C2(KEYINPUT23), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT72), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n206), .B1(new_n256), .B2(new_n258), .ZN(new_n523));
  OAI21_X1  g337(.A(KEYINPUT23), .B1(new_n523), .B2(new_n513), .ZN(new_n524));
  INV_X1    g338(.A(new_n520), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n522), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n521), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n519), .B1(new_n527), .B2(G110), .ZN(new_n528));
  INV_X1    g342(.A(G110), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n524), .A2(new_n529), .A3(new_n525), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n530), .B1(new_n516), .B2(new_n517), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n380), .B1(new_n243), .B2(new_n377), .ZN(new_n532));
  AND2_X1   g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n512), .B1(new_n528), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n531), .A2(new_n532), .ZN(new_n535));
  INV_X1    g349(.A(new_n512), .ZN(new_n536));
  NOR3_X1   g350(.A1(new_n521), .A2(new_n526), .A3(new_n529), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n535), .B(new_n536), .C1(new_n537), .C2(new_n519), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n534), .A2(new_n187), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(KEYINPUT25), .ZN(new_n540));
  INV_X1    g354(.A(new_n348), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n541), .B1(G234), .B2(new_n187), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT25), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n534), .A2(new_n543), .A3(new_n187), .A4(new_n538), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n540), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT73), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n534), .A2(new_n538), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n542), .A2(G902), .ZN(new_n550));
  AOI21_X1  g364(.A(KEYINPUT74), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  AND4_X1   g365(.A1(KEYINPUT74), .A2(new_n534), .A3(new_n538), .A4(new_n550), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n540), .A2(KEYINPUT73), .A3(new_n542), .A4(new_n544), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n547), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n509), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(G469), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n251), .B1(G128), .B2(new_n265), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n253), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(new_n205), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n204), .A2(new_n253), .A3(new_n263), .A4(new_n267), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n453), .A2(new_n454), .ZN(new_n564));
  AOI21_X1  g378(.A(KEYINPUT12), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT12), .ZN(new_n566));
  INV_X1    g380(.A(new_n564), .ZN(new_n567));
  AOI211_X1 g381(.A(new_n566), .B(new_n567), .C1(new_n561), .C2(new_n562), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n238), .A2(new_n237), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n234), .A2(G101), .A3(new_n235), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n283), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT10), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n558), .B1(new_n250), .B2(new_n252), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n574), .B1(new_n575), .B2(new_n204), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n456), .A2(KEYINPUT10), .A3(new_n205), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT78), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n564), .B(new_n578), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n573), .A2(new_n576), .A3(new_n577), .A4(new_n579), .ZN(new_n580));
  XNOR2_X1  g394(.A(G110), .B(G140), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n581), .B(KEYINPUT75), .ZN(new_n582));
  AND2_X1   g396(.A1(new_n347), .A2(G227), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n582), .B(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n580), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n569), .A2(new_n586), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n577), .B(new_n576), .C1(new_n239), .C2(new_n284), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n564), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n585), .B1(new_n589), .B2(new_n580), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n557), .B(new_n187), .C1(new_n587), .C2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(G469), .A2(G902), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n580), .B1(new_n565), .B2(new_n568), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n584), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n589), .A2(new_n580), .A3(new_n585), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n594), .A2(G469), .A3(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n591), .A2(new_n592), .A3(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(G221), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n598), .B1(new_n346), .B2(new_n187), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n597), .A2(KEYINPUT79), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(KEYINPUT79), .B1(new_n597), .B2(new_n600), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n445), .A2(new_n556), .A3(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(G101), .ZN(G3));
  INV_X1    g419(.A(KEYINPUT33), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n358), .A2(new_n606), .A3(new_n359), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n350), .A2(KEYINPUT33), .A3(new_n357), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n607), .A2(new_n187), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(G478), .ZN(new_n610));
  OR2_X1    g424(.A1(new_n436), .A2(G478), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(KEYINPUT96), .ZN(new_n613));
  INV_X1    g427(.A(new_n372), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n427), .A2(new_n434), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n411), .A2(G475), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT96), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n610), .A2(new_n618), .A3(new_n611), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n613), .A2(new_n614), .A3(new_n617), .A4(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n309), .A2(new_n310), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g436(.A(G472), .B1(new_n507), .B2(G902), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n501), .A2(new_n505), .ZN(new_n624));
  AND2_X1   g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n555), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n597), .A2(new_n600), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT79), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n597), .A2(KEYINPUT79), .A3(new_n600), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n625), .A2(new_n626), .A3(new_n629), .A4(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n622), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT34), .B(G104), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G6));
  NAND3_X1  g449(.A1(new_n364), .A2(new_n437), .A3(new_n438), .ZN(new_n636));
  INV_X1    g450(.A(new_n310), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n637), .B1(new_n307), .B2(new_n308), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n616), .B(KEYINPUT97), .ZN(new_n639));
  AND2_X1   g453(.A1(new_n639), .A2(new_n615), .ZN(new_n640));
  XOR2_X1   g454(.A(new_n372), .B(KEYINPUT98), .Z(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  AND4_X1   g456(.A1(new_n636), .A2(new_n638), .A3(new_n640), .A4(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n632), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT99), .B(KEYINPUT35), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(new_n192), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n644), .B(new_n646), .ZN(G9));
  NOR2_X1   g461(.A1(new_n512), .A2(KEYINPUT36), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(KEYINPUT100), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n528), .A2(new_n533), .ZN(new_n650));
  XOR2_X1   g464(.A(new_n649), .B(new_n650), .Z(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n550), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n547), .A2(new_n554), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(KEYINPUT101), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT101), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n547), .A2(new_n652), .A3(new_n655), .A4(new_n554), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  AND2_X1   g471(.A1(new_n657), .A2(new_n603), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n445), .A2(new_n658), .A3(new_n625), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(KEYINPUT37), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(new_n529), .ZN(G12));
  AND3_X1   g475(.A1(new_n364), .A2(new_n437), .A3(new_n438), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n366), .B1(new_n370), .B2(G900), .ZN(new_n663));
  AND3_X1   g477(.A1(new_n639), .A2(new_n615), .A3(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n621), .A2(new_n509), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n658), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G128), .ZN(G30));
  XOR2_X1   g483(.A(new_n663), .B(KEYINPUT39), .Z(new_n670));
  NOR3_X1   g484(.A1(new_n601), .A2(new_n602), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(new_n671), .B(KEYINPUT40), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n309), .B(KEYINPUT38), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n506), .A2(new_n508), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n487), .B1(new_n485), .B2(new_n462), .ZN(new_n675));
  AND2_X1   g489(.A1(new_n494), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g490(.A(G472), .B1(new_n676), .B2(G902), .ZN(new_n677));
  AND2_X1   g491(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n617), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n662), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n673), .A2(new_n679), .A3(new_n310), .A4(new_n681), .ZN(new_n682));
  OR3_X1    g496(.A1(new_n672), .A2(new_n653), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G143), .ZN(G45));
  AND3_X1   g498(.A1(new_n610), .A2(new_n618), .A3(new_n611), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n618), .B1(new_n610), .B2(new_n611), .ZN(new_n686));
  NOR3_X1   g500(.A1(new_n685), .A2(new_n686), .A3(new_n680), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n687), .A2(new_n658), .A3(new_n663), .A4(new_n667), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G146), .ZN(G48));
  OAI21_X1  g503(.A(new_n187), .B1(new_n587), .B2(new_n590), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(G469), .ZN(new_n691));
  AND3_X1   g505(.A1(new_n691), .A2(KEYINPUT102), .A3(new_n591), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT102), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n690), .A2(new_n693), .A3(G469), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n600), .B1(new_n692), .B2(new_n695), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n696), .A2(new_n509), .A3(new_n555), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n687), .A2(new_n614), .A3(new_n697), .A4(new_n638), .ZN(new_n698));
  XNOR2_X1  g512(.A(KEYINPUT41), .B(G113), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G15));
  NAND2_X1  g514(.A1(new_n643), .A2(new_n697), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G116), .ZN(G18));
  NAND2_X1  g516(.A1(new_n440), .A2(new_n444), .ZN(new_n703));
  INV_X1    g517(.A(new_n490), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n674), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n621), .A2(new_n696), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n703), .A2(new_n705), .A3(new_n706), .A4(new_n657), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G119), .ZN(G21));
  NAND3_X1  g522(.A1(new_n691), .A2(KEYINPUT102), .A3(new_n591), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n599), .B1(new_n709), .B2(new_n694), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n638), .A2(new_n636), .A3(new_n710), .A4(new_n617), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n498), .B1(new_n476), .B2(new_n486), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n505), .ZN(new_n713));
  AND2_X1   g527(.A1(new_n713), .A2(new_n623), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n714), .A2(new_n626), .A3(new_n642), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  XOR2_X1   g530(.A(new_n716), .B(G122), .Z(G24));
  AND2_X1   g531(.A1(new_n714), .A2(new_n653), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n687), .A2(new_n663), .A3(new_n706), .A4(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G125), .ZN(G27));
  INV_X1    g534(.A(KEYINPUT42), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n307), .A2(new_n308), .A3(new_n310), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT103), .ZN(new_n723));
  AND3_X1   g537(.A1(new_n597), .A2(new_n723), .A3(new_n600), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n723), .B1(new_n597), .B2(new_n600), .ZN(new_n725));
  NOR3_X1   g539(.A1(new_n722), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n556), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n613), .A2(new_n617), .A3(new_n619), .A4(new_n663), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n721), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n687), .A2(new_n663), .A3(new_n726), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT104), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n502), .B1(new_n501), .B2(new_n505), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n507), .A2(KEYINPUT32), .A3(new_n504), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n731), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n506), .A2(new_n508), .A3(KEYINPUT104), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n734), .A2(new_n704), .A3(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n736), .A2(KEYINPUT42), .A3(new_n626), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n729), .B1(new_n730), .B2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G131), .ZN(G33));
  NAND3_X1  g553(.A1(new_n666), .A2(new_n726), .A3(new_n556), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G134), .ZN(G36));
  XNOR2_X1  g555(.A(new_n722), .B(KEYINPUT107), .ZN(new_n742));
  INV_X1    g556(.A(new_n625), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n613), .A2(new_n619), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT106), .ZN(new_n745));
  AOI21_X1  g559(.A(KEYINPUT43), .B1(new_n680), .B2(new_n745), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n744), .A2(new_n617), .A3(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n746), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n685), .A2(new_n686), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n748), .B1(new_n749), .B2(new_n680), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n743), .B(new_n653), .C1(new_n747), .C2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT44), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n742), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(KEYINPUT108), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n594), .A2(new_n595), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(KEYINPUT45), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(G469), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n757), .A2(KEYINPUT46), .A3(new_n592), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(KEYINPUT105), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT46), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n760), .B(G469), .C1(new_n756), .C2(G902), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT105), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n757), .A2(new_n762), .A3(KEYINPUT46), .A4(new_n592), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n759), .A2(new_n761), .A3(new_n591), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(new_n600), .ZN(new_n765));
  AOI211_X1 g579(.A(new_n670), .B(new_n765), .C1(new_n751), .C2(new_n752), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT108), .ZN(new_n767));
  OAI211_X1 g581(.A(new_n767), .B(new_n742), .C1(new_n751), .C2(new_n752), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n754), .A2(new_n766), .A3(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G137), .ZN(G39));
  INV_X1    g584(.A(KEYINPUT47), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n765), .B(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n728), .A2(new_n722), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n773), .A2(new_n509), .A3(new_n555), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n774), .A2(KEYINPUT109), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n774), .A2(KEYINPUT109), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n772), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT110), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n772), .B(KEYINPUT110), .C1(new_n775), .C2(new_n776), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G140), .ZN(G42));
  NOR2_X1   g596(.A1(new_n747), .A2(new_n750), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n783), .A2(new_n366), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n784), .A2(new_n626), .A3(new_n714), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n673), .A2(new_n310), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n785), .A2(new_n710), .A3(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(KEYINPUT50), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n692), .A2(new_n695), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n790), .A2(new_n600), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n785), .B(new_n742), .C1(new_n772), .C2(new_n791), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n696), .A2(new_n722), .ZN(new_n793));
  AND4_X1   g607(.A1(new_n626), .A2(new_n793), .A3(new_n367), .A4(new_n678), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n794), .A2(new_n680), .A3(new_n744), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n784), .A2(new_n718), .A3(new_n793), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n792), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n789), .A2(KEYINPUT51), .A3(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT51), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n800), .B1(new_n788), .B2(new_n797), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n678), .A2(new_n653), .ZN(new_n804));
  INV_X1    g618(.A(new_n627), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n638), .A2(new_n636), .A3(new_n617), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n804), .A2(new_n805), .A3(new_n806), .A4(new_n663), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n688), .A2(new_n719), .A3(new_n807), .A4(new_n668), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(KEYINPUT52), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT114), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n604), .A2(new_n659), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n666), .A2(new_n556), .A3(new_n726), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n657), .A2(new_n603), .A3(new_n662), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n665), .A2(new_n509), .A3(new_n722), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n813), .A2(KEYINPUT113), .A3(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT113), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n657), .A2(new_n603), .A3(new_n662), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n307), .A2(new_n308), .A3(new_n310), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n705), .A2(new_n818), .A3(new_n664), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n816), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n812), .B1(new_n815), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n309), .A2(new_n311), .A3(new_n642), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n631), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n613), .A2(KEYINPUT112), .A3(new_n617), .A4(new_n619), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT112), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n825), .B1(new_n662), .B2(new_n617), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n823), .B(new_n824), .C1(new_n687), .C2(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n687), .A2(new_n663), .A3(new_n718), .A4(new_n726), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n811), .A2(new_n821), .A3(new_n827), .A4(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n716), .B1(new_n622), .B2(new_n697), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n707), .A2(new_n701), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n738), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n810), .B1(new_n829), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(KEYINPUT113), .B1(new_n813), .B2(new_n814), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n817), .A2(new_n819), .A3(new_n816), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n740), .B(new_n828), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n827), .A2(new_n604), .A3(new_n659), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n687), .A2(new_n556), .A3(new_n663), .A4(new_n726), .ZN(new_n839));
  OR3_X1    g653(.A1(new_n722), .A2(new_n724), .A3(new_n725), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n728), .A2(new_n840), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n736), .A2(KEYINPUT42), .A3(new_n626), .ZN(new_n842));
  AOI22_X1  g656(.A1(new_n839), .A2(new_n721), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n716), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n698), .A2(new_n707), .A3(new_n844), .A4(new_n701), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n838), .A2(new_n846), .A3(KEYINPUT114), .ZN(new_n847));
  AOI211_X1 g661(.A(new_n803), .B(new_n809), .C1(new_n833), .C2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n833), .A2(new_n847), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT52), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n808), .B(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(KEYINPUT53), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(KEYINPUT54), .B1(new_n848), .B2(new_n852), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n736), .A2(new_n626), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n784), .A2(new_n854), .A3(new_n793), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT48), .ZN(new_n856));
  OR2_X1    g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT54), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT115), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n832), .B1(new_n829), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n838), .A2(KEYINPUT115), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n860), .A2(KEYINPUT53), .A3(new_n851), .A4(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n809), .B1(new_n833), .B2(new_n847), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n858), .B(new_n862), .C1(new_n863), .C2(KEYINPUT53), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n855), .A2(new_n856), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n853), .A2(new_n857), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n785), .A2(new_n706), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n794), .A2(new_n687), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n867), .A2(G952), .A3(new_n347), .A4(new_n868), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n869), .B(KEYINPUT116), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n802), .A2(new_n866), .A3(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(G952), .A2(G953), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n600), .A2(new_n311), .ZN(new_n873));
  NOR4_X1   g687(.A1(new_n744), .A2(new_n555), .A3(new_n617), .A4(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n874), .A2(KEYINPUT111), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n673), .B1(new_n874), .B2(KEYINPUT111), .ZN(new_n876));
  XOR2_X1   g690(.A(new_n790), .B(KEYINPUT49), .Z(new_n877));
  NAND3_X1  g691(.A1(new_n876), .A2(new_n678), .A3(new_n877), .ZN(new_n878));
  OAI22_X1  g692(.A1(new_n871), .A2(new_n872), .B1(new_n875), .B2(new_n878), .ZN(G75));
  NOR3_X1   g693(.A1(new_n829), .A2(new_n832), .A3(new_n810), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT114), .B1(new_n838), .B2(new_n846), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n851), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(new_n803), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n187), .B1(new_n883), .B2(new_n862), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(G210), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT56), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n301), .A2(new_n299), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT117), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT55), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n889), .B(new_n296), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n885), .A2(new_n886), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n890), .B1(new_n885), .B2(new_n886), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n347), .A2(G952), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT118), .Z(new_n894));
  NOR3_X1   g708(.A1(new_n891), .A2(new_n892), .A3(new_n894), .ZN(G51));
  NAND2_X1  g709(.A1(new_n592), .A2(KEYINPUT57), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n858), .B1(new_n883), .B2(new_n862), .ZN(new_n897));
  INV_X1    g711(.A(new_n864), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n592), .A2(KEYINPUT57), .ZN(new_n900));
  OAI22_X1  g714(.A1(new_n899), .A2(new_n900), .B1(new_n590), .B2(new_n587), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n757), .B(KEYINPUT119), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n884), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n893), .B1(new_n901), .B2(new_n903), .ZN(G54));
  NAND3_X1  g718(.A1(new_n884), .A2(KEYINPUT58), .A3(G475), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n905), .A2(new_n424), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n905), .A2(new_n424), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n906), .A2(new_n907), .A3(new_n893), .ZN(G60));
  NAND2_X1  g722(.A1(new_n607), .A2(new_n608), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT120), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(G478), .A2(G902), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(KEYINPUT59), .Z(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  OAI211_X1 g728(.A(new_n911), .B(new_n914), .C1(new_n897), .C2(new_n898), .ZN(new_n915));
  INV_X1    g729(.A(new_n894), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n913), .B1(new_n853), .B2(new_n864), .ZN(new_n917));
  OAI211_X1 g731(.A(new_n915), .B(new_n916), .C1(new_n917), .C2(new_n911), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT121), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n863), .A2(KEYINPUT53), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n858), .B1(new_n883), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n914), .B1(new_n922), .B2(new_n898), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n894), .B1(new_n923), .B2(new_n910), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n924), .A2(KEYINPUT121), .A3(new_n915), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n920), .A2(new_n925), .ZN(G63));
  NAND2_X1  g740(.A1(new_n883), .A2(new_n862), .ZN(new_n927));
  NAND2_X1  g741(.A1(G217), .A2(G902), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT60), .Z(new_n929));
  NAND3_X1  g743(.A1(new_n927), .A2(new_n651), .A3(new_n929), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n927), .A2(new_n929), .ZN(new_n931));
  OAI211_X1 g745(.A(new_n916), .B(new_n930), .C1(new_n931), .C2(new_n549), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT61), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n932), .B(new_n933), .ZN(G66));
  OR2_X1    g748(.A1(new_n837), .A2(new_n845), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(new_n347), .ZN(new_n936));
  OAI21_X1  g750(.A(G953), .B1(new_n369), .B2(new_n275), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n888), .B1(G898), .B2(new_n347), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n938), .B(new_n939), .ZN(G69));
  AOI21_X1  g754(.A(new_n347), .B1(G227), .B2(G900), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n481), .B1(new_n471), .B2(KEYINPUT30), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n415), .A2(new_n416), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT122), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n942), .B(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(G900), .A2(G953), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n765), .A2(new_n670), .ZN(new_n947));
  AND3_X1   g761(.A1(new_n947), .A2(new_n854), .A3(new_n806), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT127), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n843), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OR2_X1    g764(.A1(new_n948), .A2(new_n949), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n769), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT124), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n719), .A2(new_n668), .ZN(new_n954));
  INV_X1    g768(.A(new_n688), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n953), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n688), .A2(new_n719), .A3(KEYINPUT124), .A4(new_n668), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n958), .B1(new_n779), .B2(new_n780), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n952), .A2(new_n740), .A3(new_n959), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n945), .B(new_n946), .C1(new_n960), .C2(G953), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT126), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n941), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n956), .A2(new_n683), .A3(new_n957), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT62), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n964), .B(new_n965), .ZN(new_n966));
  OR2_X1    g780(.A1(new_n687), .A2(new_n826), .ZN(new_n967));
  AOI21_X1  g781(.A(KEYINPUT125), .B1(new_n967), .B2(new_n824), .ZN(new_n968));
  INV_X1    g782(.A(new_n556), .ZN(new_n969));
  NOR3_X1   g783(.A1(new_n968), .A2(new_n969), .A3(new_n722), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n967), .A2(KEYINPUT125), .A3(new_n824), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n970), .A2(new_n671), .A3(new_n971), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n966), .A2(new_n769), .A3(new_n781), .A4(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n347), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n945), .B(KEYINPUT123), .Z(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n961), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n963), .A2(new_n977), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n961), .B(new_n976), .C1(new_n962), .C2(new_n941), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n978), .A2(new_n979), .ZN(G72));
  INV_X1    g794(.A(new_n893), .ZN(new_n981));
  NAND2_X1  g795(.A1(G472), .A2(G902), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n982), .B(KEYINPUT63), .Z(new_n983));
  OAI21_X1  g797(.A(new_n983), .B1(new_n960), .B2(new_n935), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n984), .A2(new_n487), .A3(new_n483), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n494), .B1(new_n483), .B2(new_n476), .ZN(new_n986));
  OAI211_X1 g800(.A(new_n983), .B(new_n986), .C1(new_n848), .C2(new_n852), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n983), .B1(new_n973), .B2(new_n935), .ZN(new_n988));
  INV_X1    g802(.A(new_n483), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n988), .A2(new_n476), .A3(new_n989), .ZN(new_n990));
  AND4_X1   g804(.A1(new_n981), .A2(new_n985), .A3(new_n987), .A4(new_n990), .ZN(G57));
endmodule


