//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 0 1 0 0 1 1 1 1 0 1 1 0 0 1 1 1 0 1 0 1 0 0 0 0 0 0 1 1 1 1 1 0 0 0 0 0 1 1 0 0 0 0 0 0 1 0 0 1 0 0 1 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:42 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1298, new_n1299, new_n1300, new_n1302, new_n1303,
    new_n1304, new_n1305, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370, new_n1371,
    new_n1372, new_n1373, new_n1374, new_n1375, new_n1376, new_n1377,
    new_n1378, new_n1379, new_n1380, new_n1381, new_n1382;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G107), .A2(G264), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n212));
  AND4_X1   g0012(.A1(new_n209), .A2(new_n210), .A3(new_n211), .A4(new_n212), .ZN(new_n213));
  XNOR2_X1  g0013(.A(KEYINPUT65), .B(G238), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G68), .ZN(new_n216));
  AOI21_X1  g0016(.A(new_n208), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(KEYINPUT1), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT66), .Z(new_n220));
  INV_X1    g0020(.A(G13), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n208), .A2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT0), .ZN(new_n225));
  INV_X1    g0025(.A(new_n202), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(G50), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n229), .A2(new_n207), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n225), .B(new_n231), .C1(new_n218), .C2(new_n217), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n220), .A2(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G264), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G50), .B(G58), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT67), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G68), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(G41), .ZN(new_n250));
  OAI211_X1 g0050(.A(new_n206), .B(G45), .C1(new_n250), .C2(KEYINPUT5), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(KEYINPUT78), .ZN(new_n252));
  INV_X1    g0052(.A(G45), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n253), .A2(G1), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT78), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT5), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G41), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n254), .A2(new_n255), .A3(new_n257), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n256), .A2(G41), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G274), .ZN(new_n261));
  AND2_X1   g0061(.A1(G1), .A2(G13), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G33), .A2(G41), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n261), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND4_X1  g0064(.A1(new_n252), .A2(new_n258), .A3(new_n260), .A4(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n262), .A2(new_n263), .ZN(new_n266));
  OAI211_X1 g0066(.A(new_n266), .B(G270), .C1(new_n251), .C2(new_n259), .ZN(new_n267));
  AND2_X1   g0067(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT84), .ZN(new_n269));
  AND2_X1   g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  NOR2_X1   g0070(.A1(KEYINPUT3), .A2(G33), .ZN(new_n271));
  OAI211_X1 g0071(.A(G264), .B(G1698), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G1698), .ZN(new_n273));
  OAI211_X1 g0073(.A(G257), .B(new_n273), .C1(new_n270), .C2(new_n271), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT3), .ZN(new_n275));
  INV_X1    g0075(.A(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(KEYINPUT3), .A2(G33), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n277), .A2(G303), .A3(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n272), .A2(new_n274), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(KEYINPUT83), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT83), .ZN(new_n282));
  NAND4_X1  g0082(.A1(new_n272), .A2(new_n274), .A3(new_n282), .A4(new_n279), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT69), .ZN(new_n285));
  AND2_X1   g0085(.A1(G33), .A2(G41), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n285), .B1(new_n286), .B2(new_n229), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n262), .A2(KEYINPUT69), .A3(new_n263), .ZN(new_n288));
  AND2_X1   g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n269), .B1(new_n284), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n287), .A2(new_n288), .ZN(new_n291));
  AOI211_X1 g0091(.A(KEYINPUT84), .B(new_n291), .C1(new_n281), .C2(new_n283), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n268), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT21), .ZN(new_n294));
  INV_X1    g0094(.A(G169), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n221), .A2(G1), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G116), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G20), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(G33), .A2(G283), .ZN(new_n301));
  INV_X1    g0101(.A(G97), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n301), .B(new_n207), .C1(G33), .C2(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(new_n229), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n303), .A2(new_n305), .A3(new_n299), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT20), .ZN(new_n307));
  OR2_X1    g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n306), .A2(new_n307), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n300), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n276), .A2(G1), .ZN(new_n311));
  XNOR2_X1  g0111(.A(new_n311), .B(KEYINPUT77), .ZN(new_n312));
  AND2_X1   g0112(.A1(new_n312), .A2(G116), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT71), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n314), .B1(new_n316), .B2(new_n305), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n315), .A2(KEYINPUT71), .A3(new_n229), .A4(new_n304), .ZN(new_n318));
  AND2_X1   g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n313), .A2(new_n319), .ZN(new_n320));
  AOI211_X1 g0120(.A(new_n294), .B(new_n295), .C1(new_n310), .C2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n293), .A2(new_n321), .ZN(new_n322));
  AND3_X1   g0122(.A1(new_n265), .A2(G179), .A3(new_n267), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n324), .B1(new_n310), .B2(new_n320), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n325), .B1(new_n292), .B2(new_n290), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n322), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n295), .B1(new_n310), .B2(new_n320), .ZN(new_n328));
  AOI21_X1  g0128(.A(KEYINPUT21), .B1(new_n293), .B2(new_n328), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(G1698), .B1(new_n277), .B2(new_n278), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G222), .ZN(new_n332));
  INV_X1    g0132(.A(G77), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n277), .A2(new_n278), .ZN(new_n334));
  INV_X1    g0134(.A(G223), .ZN(new_n335));
  OAI21_X1  g0135(.A(G1698), .B1(new_n270), .B2(new_n271), .ZN(new_n336));
  OAI221_X1 g0136(.A(new_n332), .B1(new_n333), .B2(new_n334), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n289), .ZN(new_n338));
  AOI21_X1  g0138(.A(G1), .B1(new_n250), .B2(new_n253), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n266), .A2(G274), .A3(new_n339), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n266), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(G226), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n340), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT68), .ZN(new_n345));
  OR2_X1    g0145(.A1(new_n344), .A2(KEYINPUT68), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n338), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  OR2_X1    g0147(.A1(new_n347), .A2(G179), .ZN(new_n348));
  INV_X1    g0148(.A(new_n305), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n203), .A2(G20), .ZN(new_n350));
  XNOR2_X1  g0150(.A(KEYINPUT8), .B(G58), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n207), .A2(G33), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  NOR2_X1   g0154(.A1(G20), .A2(G33), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n352), .A2(new_n354), .B1(G150), .B2(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n349), .B1(new_n350), .B2(new_n356), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n316), .A2(new_n305), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n206), .A2(G20), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n358), .A2(G50), .A3(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n360), .B1(G50), .B2(new_n315), .ZN(new_n361));
  OR2_X1    g0161(.A1(new_n357), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n347), .A2(new_n295), .ZN(new_n363));
  AND3_X1   g0163(.A1(new_n348), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT9), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  OR3_X1    g0166(.A1(new_n357), .A2(new_n361), .A3(new_n365), .ZN(new_n367));
  AND2_X1   g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT10), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n338), .A2(G190), .A3(new_n346), .A4(new_n345), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n347), .A2(G200), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n368), .A2(new_n369), .A3(new_n370), .A4(new_n371), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n371), .A2(new_n366), .A3(new_n370), .A4(new_n367), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(KEYINPUT10), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n364), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n319), .A2(G68), .A3(new_n359), .ZN(new_n376));
  INV_X1    g0176(.A(G68), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n355), .A2(G50), .B1(G20), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n378), .B1(new_n333), .B2(new_n353), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n305), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT11), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n316), .A2(new_n377), .ZN(new_n383));
  XNOR2_X1  g0183(.A(new_n383), .B(KEYINPUT12), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n379), .A2(KEYINPUT11), .A3(new_n305), .ZN(new_n385));
  AND4_X1   g0185(.A1(new_n376), .A2(new_n382), .A3(new_n384), .A4(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n343), .A2(new_n273), .ZN(new_n387));
  INV_X1    g0187(.A(G232), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(G1698), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n387), .B(new_n389), .C1(new_n270), .C2(new_n271), .ZN(new_n390));
  NAND2_X1  g0190(.A1(G33), .A2(G97), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n289), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT13), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n250), .A2(new_n253), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n206), .A2(new_n395), .B1(new_n262), .B2(new_n263), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n396), .A2(G238), .B1(new_n264), .B2(new_n339), .ZN(new_n397));
  AND3_X1   g0197(.A1(new_n393), .A2(new_n394), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n394), .B1(new_n393), .B2(new_n397), .ZN(new_n399));
  OAI21_X1  g0199(.A(G200), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n291), .B1(new_n391), .B2(new_n390), .ZN(new_n401));
  INV_X1    g0201(.A(G238), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n340), .B1(new_n342), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(KEYINPUT13), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n393), .A2(new_n394), .A3(new_n397), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n404), .A2(G190), .A3(new_n405), .ZN(new_n406));
  AND3_X1   g0206(.A1(new_n386), .A2(new_n400), .A3(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(G169), .B1(new_n398), .B2(new_n399), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(KEYINPUT14), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n404), .A2(G179), .A3(new_n405), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT14), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n411), .B(G169), .C1(new_n398), .C2(new_n399), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n409), .A2(new_n410), .A3(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n386), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n407), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  OAI211_X1 g0215(.A(G232), .B(new_n273), .C1(new_n270), .C2(new_n271), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(KEYINPUT70), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT70), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n334), .A2(new_n418), .A3(G232), .A4(new_n273), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n277), .A2(G107), .A3(new_n278), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n421), .B1(new_n336), .B2(new_n214), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n291), .B1(new_n420), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(G244), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n340), .B1(new_n342), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g0226(.A(G200), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(G20), .A2(G77), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n207), .A2(new_n276), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n428), .B1(new_n351), .B2(new_n429), .ZN(new_n430));
  XNOR2_X1  g0230(.A(KEYINPUT15), .B(G87), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n431), .A2(new_n353), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n305), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n316), .A2(new_n333), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n333), .B1(new_n206), .B2(G20), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n317), .A2(new_n318), .A3(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT72), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n317), .A2(KEYINPUT72), .A3(new_n318), .A4(new_n436), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n435), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n426), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n422), .B1(new_n419), .B2(new_n417), .ZN(new_n443));
  OAI211_X1 g0243(.A(G190), .B(new_n442), .C1(new_n443), .C2(new_n291), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n427), .A2(new_n441), .A3(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n442), .B1(new_n443), .B2(new_n291), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n439), .A2(new_n440), .ZN(new_n447));
  AND2_X1   g0247(.A1(new_n433), .A2(new_n434), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n446), .A2(new_n295), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(G179), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n450), .B(new_n442), .C1(new_n443), .C2(new_n291), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n375), .A2(new_n415), .A3(new_n445), .A4(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT75), .ZN(new_n454));
  NAND2_X1  g0254(.A1(G33), .A2(G87), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n335), .A2(new_n273), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n343), .A2(G1698), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n270), .A2(new_n271), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n455), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n289), .A2(new_n460), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n396), .A2(G232), .B1(new_n264), .B2(new_n339), .ZN(new_n462));
  AND3_X1   g0262(.A1(new_n461), .A2(G179), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n295), .B1(new_n461), .B2(new_n462), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n454), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n461), .A2(G179), .A3(new_n462), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n266), .A2(G232), .A3(new_n341), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n340), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n468), .B1(new_n289), .B2(new_n460), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n466), .B(KEYINPUT75), .C1(new_n469), .C2(new_n295), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n351), .B1(new_n206), .B2(G20), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n472), .A2(new_n358), .B1(new_n316), .B2(new_n351), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT74), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n459), .A2(new_n475), .A3(KEYINPUT7), .A4(new_n207), .ZN(new_n476));
  XNOR2_X1  g0276(.A(KEYINPUT73), .B(KEYINPUT7), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n477), .B1(new_n207), .B2(new_n459), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n277), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n278), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(KEYINPUT74), .ZN(new_n480));
  OAI211_X1 g0280(.A(G68), .B(new_n476), .C1(new_n478), .C2(new_n480), .ZN(new_n481));
  XNOR2_X1  g0281(.A(G58), .B(G68), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n482), .A2(G20), .B1(G159), .B2(new_n355), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT16), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n482), .A2(G20), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n355), .A2(G159), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n277), .A2(new_n207), .A3(new_n278), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n377), .B1(new_n490), .B2(KEYINPUT7), .ZN(new_n491));
  OR2_X1    g0291(.A1(new_n490), .A2(new_n477), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n489), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n349), .B1(new_n493), .B2(KEYINPUT16), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n474), .B1(new_n486), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(KEYINPUT18), .B1(new_n471), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(G190), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n461), .A2(new_n497), .A3(new_n462), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n498), .B1(new_n469), .B2(G200), .ZN(new_n499));
  AOI21_X1  g0299(.A(KEYINPUT16), .B1(new_n481), .B2(new_n483), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n490), .A2(KEYINPUT7), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(G68), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n490), .A2(new_n477), .ZN(new_n503));
  OAI211_X1 g0303(.A(KEYINPUT16), .B(new_n483), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n305), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n499), .B(new_n473), .C1(new_n500), .C2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT17), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n495), .A2(KEYINPUT17), .A3(new_n499), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n473), .B1(new_n505), .B2(new_n500), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT18), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n510), .A2(new_n511), .A3(new_n465), .A4(new_n470), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n496), .A2(new_n508), .A3(new_n509), .A4(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n453), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n293), .A2(G200), .ZN(new_n515));
  AND2_X1   g0315(.A1(new_n310), .A2(new_n320), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n515), .B(new_n516), .C1(new_n497), .C2(new_n293), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT79), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n266), .B(G257), .C1(new_n251), .C2(new_n259), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n265), .A2(new_n519), .ZN(new_n520));
  OAI211_X1 g0320(.A(G244), .B(new_n273), .C1(new_n270), .C2(new_n271), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT4), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n334), .A2(KEYINPUT4), .A3(G244), .A4(new_n273), .ZN(new_n524));
  OAI211_X1 g0324(.A(G250), .B(G1698), .C1(new_n270), .C2(new_n271), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n523), .A2(new_n524), .A3(new_n301), .A4(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n520), .B1(new_n289), .B2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(G200), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n518), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n316), .A2(new_n302), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n312), .A2(new_n358), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n530), .B1(new_n531), .B2(new_n302), .ZN(new_n532));
  INV_X1    g0332(.A(G107), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n533), .A2(KEYINPUT6), .A3(G97), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n302), .A2(new_n533), .ZN(new_n535));
  NOR2_X1   g0335(.A1(G97), .A2(G107), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n534), .B1(new_n537), .B2(KEYINPUT6), .ZN(new_n538));
  OAI21_X1  g0338(.A(KEYINPUT76), .B1(new_n429), .B2(new_n333), .ZN(new_n539));
  OR3_X1    g0339(.A1(new_n429), .A2(KEYINPUT76), .A3(new_n333), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n538), .A2(G20), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OAI211_X1 g0341(.A(G107), .B(new_n476), .C1(new_n478), .C2(new_n480), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n532), .B1(new_n543), .B2(new_n305), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n301), .B(new_n525), .C1(new_n521), .C2(new_n522), .ZN(new_n545));
  AOI21_X1  g0345(.A(KEYINPUT4), .B1(new_n331), .B2(G244), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n289), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AND2_X1   g0347(.A1(new_n265), .A2(new_n519), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n549), .A2(KEYINPUT79), .A3(G200), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n527), .A2(G190), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n529), .A2(new_n544), .A3(new_n550), .A4(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(G20), .B1(new_n277), .B2(new_n278), .ZN(new_n553));
  XNOR2_X1  g0353(.A(KEYINPUT85), .B(KEYINPUT22), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n553), .A2(G87), .A3(new_n554), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n207), .B(G87), .C1(new_n270), .C2(new_n271), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT22), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(KEYINPUT85), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT85), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(KEYINPUT22), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n556), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n555), .A2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT24), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT23), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(new_n207), .B2(G107), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n533), .A2(KEYINPUT23), .A3(G20), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n276), .A2(new_n298), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n566), .A2(new_n567), .B1(new_n568), .B2(new_n207), .ZN(new_n569));
  AND3_X1   g0369(.A1(new_n563), .A2(new_n564), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n564), .B1(new_n563), .B2(new_n569), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n305), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n531), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(G107), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n315), .A2(G107), .ZN(new_n575));
  XNOR2_X1  g0375(.A(new_n575), .B(KEYINPUT25), .ZN(new_n576));
  AND2_X1   g0376(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  OAI211_X1 g0377(.A(G257), .B(G1698), .C1(new_n270), .C2(new_n271), .ZN(new_n578));
  OAI211_X1 g0378(.A(G250), .B(new_n273), .C1(new_n270), .C2(new_n271), .ZN(new_n579));
  NAND2_X1  g0379(.A1(G33), .A2(G294), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n289), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n286), .A2(new_n229), .ZN(new_n583));
  INV_X1    g0383(.A(new_n251), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n583), .B1(new_n584), .B2(new_n260), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(G264), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n582), .A2(new_n586), .A3(new_n265), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n587), .A2(G190), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n289), .A2(new_n581), .B1(new_n585), .B2(G264), .ZN(new_n589));
  AOI21_X1  g0389(.A(G200), .B1(new_n589), .B2(new_n265), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n572), .B(new_n577), .C1(new_n588), .C2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n547), .A2(new_n548), .A3(new_n450), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n349), .B1(new_n541), .B2(new_n542), .ZN(new_n593));
  OAI221_X1 g0393(.A(new_n592), .B1(new_n527), .B2(G169), .C1(new_n593), .C2(new_n532), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n552), .A2(new_n591), .A3(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n589), .A2(new_n450), .A3(new_n265), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n587), .A2(new_n295), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n554), .B1(new_n553), .B2(G87), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n556), .A2(new_n561), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n569), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(KEYINPUT24), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n563), .A2(new_n564), .A3(new_n569), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n349), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n574), .A2(new_n576), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n596), .B(new_n597), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT19), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n207), .A2(G33), .A3(G97), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n553), .A2(G68), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(G87), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n609), .A2(new_n302), .A3(new_n533), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT81), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g0412(.A1(G87), .A2(G97), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n613), .A2(KEYINPUT81), .A3(new_n533), .ZN(new_n614));
  NAND3_X1  g0414(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n612), .A2(new_n614), .B1(new_n207), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n608), .B1(new_n616), .B2(KEYINPUT82), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n615), .A2(new_n207), .ZN(new_n618));
  INV_X1    g0418(.A(new_n614), .ZN(new_n619));
  AOI21_X1  g0419(.A(KEYINPUT81), .B1(new_n613), .B2(new_n533), .ZN(new_n620));
  OAI211_X1 g0420(.A(KEYINPUT82), .B(new_n618), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n305), .B1(new_n617), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n431), .A2(new_n316), .ZN(new_n624));
  OR2_X1    g0424(.A1(new_n531), .A2(new_n431), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT80), .ZN(new_n627));
  OAI21_X1  g0427(.A(G274), .B1(new_n286), .B2(new_n229), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n206), .A2(G45), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n627), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n264), .A2(KEYINPUT80), .A3(new_n254), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n629), .A2(G250), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n583), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n568), .B1(new_n331), .B2(G238), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n273), .B1(new_n277), .B2(new_n278), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(G244), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n291), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n450), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n295), .B1(new_n636), .B2(new_n640), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n626), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT82), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n647), .A2(new_n621), .A3(new_n608), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n648), .A2(new_n305), .B1(new_n316), .B2(new_n431), .ZN(new_n649));
  OAI21_X1  g0449(.A(G200), .B1(new_n636), .B2(new_n640), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n573), .A2(G87), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n634), .B1(new_n630), .B2(new_n631), .ZN(new_n652));
  OAI211_X1 g0452(.A(G238), .B(new_n273), .C1(new_n270), .C2(new_n271), .ZN(new_n653));
  INV_X1    g0453(.A(new_n568), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n653), .B(new_n654), .C1(new_n336), .C2(new_n425), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n289), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n652), .A2(new_n656), .A3(G190), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n649), .A2(new_n650), .A3(new_n651), .A4(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n605), .A2(new_n644), .A3(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n595), .A2(new_n659), .ZN(new_n660));
  AND4_X1   g0460(.A1(new_n330), .A2(new_n514), .A3(new_n517), .A4(new_n660), .ZN(G372));
  INV_X1    g0461(.A(KEYINPUT86), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n636), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n652), .A2(KEYINPUT86), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n640), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  OAI211_X1 g0465(.A(new_n626), .B(new_n642), .C1(new_n665), .C2(G169), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n293), .A2(new_n328), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(new_n294), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n284), .A2(new_n289), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(KEYINPUT84), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n284), .A2(new_n269), .A3(new_n289), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AOI22_X1  g0473(.A1(new_n293), .A2(new_n321), .B1(new_n673), .B2(new_n325), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n669), .A2(new_n674), .A3(new_n605), .ZN(new_n675));
  AND4_X1   g0475(.A1(new_n623), .A2(new_n624), .A3(new_n651), .A4(new_n657), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n652), .A2(KEYINPUT86), .ZN(new_n677));
  AOI211_X1 g0477(.A(new_n662), .B(new_n634), .C1(new_n630), .C2(new_n631), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n656), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(G200), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n676), .A2(new_n680), .ZN(new_n681));
  AND4_X1   g0481(.A1(new_n552), .A2(new_n681), .A3(new_n594), .A4(new_n591), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n667), .B1(new_n675), .B2(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n592), .B1(new_n527), .B2(G169), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(new_n544), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n681), .A2(new_n666), .A3(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT26), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n685), .A2(new_n644), .A3(new_n658), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n688), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n683), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n514), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g0492(.A(new_n692), .B(KEYINPUT87), .Z(new_n693));
  NOR2_X1   g0493(.A1(new_n463), .A2(new_n464), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n510), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(KEYINPUT18), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n510), .A2(new_n695), .A3(new_n511), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n446), .A2(new_n295), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n447), .A2(new_n448), .ZN(new_n701));
  AND3_X1   g0501(.A1(new_n700), .A2(new_n701), .A3(new_n451), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n386), .A2(new_n400), .A3(new_n406), .ZN(new_n703));
  AOI22_X1  g0503(.A1(new_n413), .A2(new_n414), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  OAI211_X1 g0504(.A(new_n508), .B(new_n509), .C1(new_n704), .C2(KEYINPUT88), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n704), .A2(KEYINPUT88), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n699), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n372), .A2(new_n374), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n364), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n693), .A2(new_n709), .ZN(G369));
  OR3_X1    g0510(.A1(new_n297), .A2(KEYINPUT27), .A3(G20), .ZN(new_n711));
  OAI21_X1  g0511(.A(KEYINPUT27), .B1(new_n297), .B2(G20), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n711), .A2(G213), .A3(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(G343), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n716), .B1(new_n669), .B2(new_n674), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n605), .A2(new_n716), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n716), .B1(new_n603), .B2(new_n604), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n591), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(new_n605), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n717), .A2(new_n719), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(new_n719), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(KEYINPUT89), .ZN(new_n725));
  AOI211_X1 g0525(.A(KEYINPUT89), .B(new_n718), .C1(new_n717), .C2(new_n722), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(G330), .ZN(new_n729));
  OAI211_X1 g0529(.A(new_n330), .B(new_n517), .C1(new_n516), .C2(new_n715), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n669), .A2(new_n674), .ZN(new_n731));
  INV_X1    g0531(.A(new_n516), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n731), .A2(new_n732), .A3(new_n716), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n729), .B1(new_n730), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n719), .A2(new_n722), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n728), .A2(new_n737), .ZN(G399));
  NOR2_X1   g0538(.A1(new_n222), .A2(G41), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR3_X1   g0540(.A1(new_n619), .A2(G116), .A3(new_n620), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n740), .A2(new_n741), .A3(G1), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n742), .B1(new_n227), .B2(new_n740), .ZN(new_n743));
  XOR2_X1   g0543(.A(KEYINPUT90), .B(KEYINPUT28), .Z(new_n744));
  XNOR2_X1  g0544(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n675), .A2(new_n682), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n689), .A2(new_n687), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n747), .B1(new_n687), .B2(new_n686), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n746), .A2(new_n748), .A3(new_n666), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n749), .A2(KEYINPUT29), .A3(new_n715), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n716), .B1(new_n683), .B2(new_n690), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n750), .B1(KEYINPUT29), .B2(new_n751), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n660), .A2(new_n330), .A3(new_n517), .A4(new_n715), .ZN(new_n753));
  AND3_X1   g0553(.A1(new_n549), .A2(new_n450), .A3(new_n587), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n293), .A2(new_n679), .A3(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT30), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n290), .A2(new_n292), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n641), .A2(new_n527), .A3(new_n323), .A4(new_n589), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n756), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n323), .A2(new_n589), .A3(new_n656), .A4(new_n652), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(new_n549), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n673), .A2(new_n761), .A3(KEYINPUT30), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n755), .A2(new_n759), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(new_n716), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT31), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n763), .A2(KEYINPUT31), .A3(new_n716), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n753), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G330), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n752), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n745), .B1(new_n771), .B2(G1), .ZN(G364));
  INV_X1    g0572(.A(new_n734), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n730), .A2(new_n729), .A3(new_n733), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n221), .A2(G20), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n206), .B1(new_n775), .B2(G45), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n739), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n773), .A2(new_n774), .A3(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(G13), .A2(G33), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(G20), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n730), .A2(new_n733), .A3(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n222), .A2(new_n459), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT91), .ZN(new_n786));
  INV_X1    g0586(.A(G355), .ZN(new_n787));
  OAI22_X1  g0587(.A1(new_n786), .A2(new_n787), .B1(G116), .B2(new_n223), .ZN(new_n788));
  OR2_X1    g0588(.A1(new_n245), .A2(new_n253), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n222), .A2(new_n334), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n790), .B1(G45), .B2(new_n227), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT92), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n788), .B1(new_n789), .B2(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n229), .B1(G20), .B2(new_n295), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n783), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n778), .B1(new_n793), .B2(new_n796), .ZN(new_n797));
  NOR3_X1   g0597(.A1(new_n207), .A2(new_n450), .A3(new_n528), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(G190), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n799), .A2(KEYINPUT93), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n799), .A2(KEYINPUT93), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  XNOR2_X1  g0603(.A(KEYINPUT96), .B(G326), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n207), .A2(G190), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n528), .A2(G179), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(G283), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n207), .A2(new_n497), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(new_n807), .ZN(new_n812));
  INV_X1    g0612(.A(G303), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n450), .A2(G200), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(new_n806), .ZN(new_n815));
  INV_X1    g0615(.A(G311), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n812), .A2(new_n813), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(G179), .A2(G200), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n806), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n810), .B(new_n817), .C1(G329), .C2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n798), .A2(new_n497), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(G317), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(KEYINPUT33), .ZN(new_n825));
  OR2_X1    g0625(.A1(new_n824), .A2(KEYINPUT33), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n823), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n811), .A2(new_n814), .ZN(new_n828));
  INV_X1    g0628(.A(G322), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n459), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n207), .B1(new_n818), .B2(G190), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n830), .B1(G294), .B2(new_n832), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n805), .A2(new_n821), .A3(new_n827), .A4(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(G58), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n828), .A2(new_n835), .B1(new_n815), .B2(new_n333), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(new_n803), .B2(G50), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT94), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n831), .A2(new_n302), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n820), .A2(G159), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n840), .B(KEYINPUT32), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n839), .B(new_n841), .C1(G68), .C2(new_n823), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n334), .B1(new_n808), .B2(new_n533), .C1(new_n609), .C2(new_n812), .ZN(new_n843));
  XOR2_X1   g0643(.A(new_n843), .B(KEYINPUT95), .Z(new_n844));
  NAND2_X1  g0644(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n834), .B1(new_n838), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n797), .B1(new_n846), .B2(new_n794), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n784), .A2(new_n847), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n780), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(G396));
  NAND2_X1  g0650(.A1(new_n716), .A2(new_n701), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n445), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n452), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n702), .A2(new_n715), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT99), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  AOI22_X1  g0656(.A1(new_n445), .A2(new_n851), .B1(new_n449), .B2(new_n451), .ZN(new_n857));
  AND3_X1   g0657(.A1(new_n449), .A2(new_n451), .A3(new_n715), .ZN(new_n858));
  OAI21_X1  g0658(.A(KEYINPUT99), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n751), .B(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n778), .B1(new_n862), .B2(new_n769), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n863), .B1(new_n769), .B2(new_n862), .ZN(new_n864));
  INV_X1    g0664(.A(new_n828), .ZN(new_n865));
  INV_X1    g0665(.A(new_n815), .ZN(new_n866));
  AOI22_X1  g0666(.A1(G143), .A2(new_n865), .B1(new_n866), .B2(G159), .ZN(new_n867));
  INV_X1    g0667(.A(G150), .ZN(new_n868));
  INV_X1    g0668(.A(G137), .ZN(new_n869));
  OAI221_X1 g0669(.A(new_n867), .B1(new_n868), .B2(new_n822), .C1(new_n802), .C2(new_n869), .ZN(new_n870));
  XOR2_X1   g0670(.A(new_n870), .B(KEYINPUT34), .Z(new_n871));
  NOR2_X1   g0671(.A1(new_n831), .A2(new_n835), .ZN(new_n872));
  INV_X1    g0672(.A(G50), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n334), .B1(new_n812), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(G132), .ZN(new_n875));
  OAI22_X1  g0675(.A1(new_n808), .A2(new_n377), .B1(new_n819), .B2(new_n875), .ZN(new_n876));
  NOR4_X1   g0676(.A1(new_n871), .A2(new_n872), .A3(new_n874), .A4(new_n876), .ZN(new_n877));
  XOR2_X1   g0677(.A(KEYINPUT97), .B(G283), .Z(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n823), .A2(new_n879), .B1(G116), .B2(new_n866), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT98), .ZN(new_n881));
  OAI22_X1  g0681(.A1(new_n802), .A2(new_n813), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n812), .ZN(new_n883));
  AOI22_X1  g0683(.A1(G107), .A2(new_n883), .B1(new_n865), .B2(G294), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n884), .B1(new_n816), .B2(new_n819), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n459), .B1(new_n808), .B2(new_n609), .ZN(new_n886));
  OR3_X1    g0686(.A1(new_n885), .A2(new_n839), .A3(new_n886), .ZN(new_n887));
  AOI211_X1 g0687(.A(new_n882), .B(new_n887), .C1(new_n881), .C2(new_n880), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n794), .B1(new_n877), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n794), .A2(new_n781), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n779), .B1(new_n333), .B2(new_n890), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n889), .B(new_n891), .C1(new_n861), .C2(new_n782), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n864), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(G384));
  OR2_X1    g0694(.A1(new_n538), .A2(KEYINPUT35), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n538), .A2(KEYINPUT35), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n895), .A2(G116), .A3(new_n230), .A4(new_n896), .ZN(new_n897));
  XNOR2_X1  g0697(.A(KEYINPUT100), .B(KEYINPUT36), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n897), .B(new_n898), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n228), .B(G77), .C1(new_n835), .C2(new_n377), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n201), .A2(G68), .ZN(new_n901));
  AOI211_X1 g0701(.A(new_n206), .B(G13), .C1(new_n900), .C2(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n414), .B(new_n716), .C1(new_n413), .C2(new_n407), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n414), .A2(new_n716), .ZN(new_n905));
  AOI21_X1  g0705(.A(KEYINPUT101), .B1(new_n415), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n412), .A2(new_n410), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n404), .A2(new_n405), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n411), .B1(new_n908), .B2(G169), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n414), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n910), .A2(KEYINPUT101), .A3(new_n703), .A4(new_n905), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n904), .B1(new_n906), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n494), .B1(KEYINPUT16), .B2(new_n493), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n713), .B1(new_n914), .B2(new_n473), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n513), .A2(new_n915), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n914), .A2(new_n473), .B1(new_n694), .B2(new_n713), .ZN(new_n917));
  INV_X1    g0717(.A(new_n506), .ZN(new_n918));
  OAI21_X1  g0718(.A(KEYINPUT37), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n510), .A2(new_n465), .A3(new_n470), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n510), .A2(new_n714), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT37), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n920), .A2(new_n921), .A3(new_n922), .A4(new_n506), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n919), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n916), .A2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT38), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n916), .A2(KEYINPUT38), .A3(new_n924), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI211_X1 g0729(.A(new_n716), .B(new_n860), .C1(new_n683), .C2(new_n690), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n913), .B(new_n929), .C1(new_n930), .C2(new_n858), .ZN(new_n931));
  OR2_X1    g0731(.A1(new_n699), .A2(new_n714), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n923), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n506), .B1(new_n495), .B2(new_n694), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT102), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n696), .A2(KEYINPUT102), .A3(new_n506), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n937), .A2(new_n921), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n934), .B1(new_n939), .B2(KEYINPUT37), .ZN(new_n940));
  NAND4_X1  g0740(.A1(new_n697), .A2(new_n508), .A3(new_n509), .A4(new_n698), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n495), .A2(new_n713), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n926), .B1(new_n940), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(KEYINPUT39), .B1(new_n944), .B2(new_n928), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n413), .A2(new_n414), .A3(new_n715), .ZN(new_n946));
  AND3_X1   g0746(.A1(new_n916), .A2(KEYINPUT38), .A3(new_n924), .ZN(new_n947));
  AOI21_X1  g0747(.A(KEYINPUT38), .B1(new_n916), .B2(new_n924), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT39), .ZN(new_n949));
  NOR3_X1   g0749(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NOR3_X1   g0750(.A1(new_n945), .A2(new_n946), .A3(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(KEYINPUT103), .B1(new_n933), .B2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n946), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n927), .A2(KEYINPUT39), .A3(new_n928), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n941), .A2(new_n942), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n942), .B1(new_n935), .B2(new_n936), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n922), .B1(new_n956), .B2(new_n938), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n955), .B1(new_n957), .B2(new_n934), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n947), .B1(new_n926), .B2(new_n958), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n953), .B(new_n954), .C1(new_n959), .C2(KEYINPUT39), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT103), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n960), .A2(new_n961), .A3(new_n931), .A4(new_n932), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n952), .A2(new_n962), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n514), .B(new_n750), .C1(KEYINPUT29), .C2(new_n751), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n709), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n963), .B(new_n965), .Z(new_n966));
  NOR3_X1   g0766(.A1(new_n947), .A2(new_n948), .A3(KEYINPUT40), .ZN(new_n967));
  NOR2_X1   g0767(.A1(KEYINPUT104), .A2(KEYINPUT31), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n763), .A2(new_n716), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n764), .A2(new_n968), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n753), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(KEYINPUT105), .A2(KEYINPUT40), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n972), .A2(new_n861), .A3(new_n913), .A4(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n967), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n972), .A2(new_n861), .A3(new_n913), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(KEYINPUT105), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n944), .A2(new_n928), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n975), .B1(new_n979), .B2(KEYINPUT40), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n514), .A2(new_n972), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT105), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n910), .A2(new_n703), .A3(new_n905), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT101), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n911), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n860), .B1(new_n987), .B2(new_n904), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n983), .B1(new_n988), .B2(new_n972), .ZN(new_n989));
  OAI21_X1  g0789(.A(KEYINPUT40), .B1(new_n989), .B2(new_n959), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT40), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n927), .A2(new_n991), .A3(new_n928), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n992), .A2(new_n972), .A3(new_n988), .A4(new_n973), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n994), .A2(new_n514), .A3(new_n972), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n982), .A2(new_n995), .A3(G330), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n966), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(new_n206), .B2(new_n775), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n966), .A2(new_n996), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n903), .B1(new_n998), .B2(new_n999), .ZN(G367));
  NAND2_X1  g0800(.A1(new_n552), .A2(new_n594), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n544), .A2(new_n715), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n1001), .A2(new_n1002), .B1(new_n594), .B2(new_n715), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1003), .B(KEYINPUT106), .Z(new_n1004));
  NOR2_X1   g0804(.A1(new_n737), .A2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT107), .ZN(new_n1006));
  AND2_X1   g0806(.A1(new_n649), .A2(new_n651), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n1007), .A2(new_n715), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1008), .A2(new_n666), .A3(new_n681), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n666), .B2(new_n1008), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1010), .A2(KEYINPUT43), .ZN(new_n1011));
  AND2_X1   g0811(.A1(new_n1006), .A2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1006), .A2(new_n1011), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1004), .A2(new_n723), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT42), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n594), .B1(new_n1004), .B2(new_n605), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n715), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1010), .A2(KEYINPUT43), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  OR3_X1    g0820(.A1(new_n1012), .A2(new_n1013), .A3(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1020), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(KEYINPUT108), .B(KEYINPUT41), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n739), .B(new_n1023), .Z(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n725), .A2(new_n727), .A3(new_n1004), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT44), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n725), .A2(new_n727), .A3(new_n1004), .A4(KEYINPUT44), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1003), .B(KEYINPUT106), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n728), .A2(KEYINPUT45), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT89), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(new_n723), .B2(new_n719), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1031), .B1(new_n1034), .B2(new_n726), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT45), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1032), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1030), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n737), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n735), .B1(new_n330), .B2(new_n716), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n723), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n734), .B(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n771), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1030), .A2(new_n1038), .A3(new_n737), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1041), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1025), .B1(new_n1048), .B2(new_n771), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1021), .B(new_n1022), .C1(new_n1049), .C2(new_n777), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n790), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n795), .B1(new_n223), .B2(new_n431), .C1(new_n240), .C2(new_n1051), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n831), .A2(new_n377), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(G58), .A2(new_n883), .B1(new_n820), .B2(G137), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1054), .B1(new_n868), .B2(new_n828), .C1(new_n201), .C2(new_n815), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n1053), .B(new_n1055), .C1(G159), .C2(new_n823), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n803), .A2(G143), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n808), .A2(new_n333), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1058), .A2(new_n459), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT109), .Z(new_n1060));
  NAND3_X1  g0860(.A1(new_n1056), .A2(new_n1057), .A3(new_n1060), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n808), .A2(new_n302), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(G317), .B2(new_n820), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(new_n813), .B2(new_n828), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n883), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT46), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(new_n812), .B2(new_n298), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1065), .B(new_n1067), .C1(new_n533), .C2(new_n831), .ZN(new_n1068));
  INV_X1    g0868(.A(G294), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n459), .B1(new_n878), .B2(new_n815), .C1(new_n822), .C2(new_n1069), .ZN(new_n1070));
  NOR3_X1   g0870(.A1(new_n1064), .A2(new_n1068), .A3(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n816), .B2(new_n802), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1061), .A2(new_n1072), .ZN(new_n1073));
  XOR2_X1   g0873(.A(new_n1073), .B(KEYINPUT47), .Z(new_n1074));
  INV_X1    g0874(.A(new_n794), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n778), .B(new_n1052), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT110), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n783), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1077), .B1(new_n1078), .B2(new_n1010), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1050), .A2(new_n1079), .ZN(G387));
  INV_X1    g0880(.A(new_n1044), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(new_n770), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1045), .A2(new_n739), .A3(new_n1082), .ZN(new_n1083));
  OR3_X1    g0883(.A1(new_n351), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1084));
  OAI21_X1  g0884(.A(KEYINPUT50), .B1(new_n351), .B2(G50), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n741), .B(new_n253), .C1(new_n377), .C2(new_n333), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT111), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1084), .B(new_n1085), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1088));
  AND2_X1   g0888(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n790), .B1(new_n237), .B2(new_n253), .C1(new_n1088), .C2(new_n1089), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n1090), .B1(G107), .B2(new_n223), .C1(new_n741), .C2(new_n786), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n779), .B1(new_n1091), .B2(new_n795), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n736), .B2(new_n1078), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n802), .A2(new_n829), .B1(new_n816), .B2(new_n822), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT112), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  OAI221_X1 g0896(.A(KEYINPUT112), .B1(new_n816), .B2(new_n822), .C1(new_n802), .C2(new_n829), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(G317), .A2(new_n865), .B1(new_n866), .B2(G303), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT48), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n832), .A2(new_n879), .B1(new_n883), .B2(G294), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1102), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT113), .ZN(new_n1104));
  AND2_X1   g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1101), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT49), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  OAI211_X1 g0909(.A(KEYINPUT49), .B(new_n1101), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n459), .B1(new_n808), .B2(new_n298), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(new_n820), .B2(new_n804), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1109), .A2(new_n1110), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(G159), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n802), .A2(new_n1114), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n459), .B(new_n1062), .C1(new_n352), .C2(new_n823), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n812), .A2(new_n333), .B1(new_n815), .B2(new_n377), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n828), .A2(new_n873), .B1(new_n819), .B2(new_n868), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n831), .A2(new_n431), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1116), .A2(new_n1119), .A3(new_n1121), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1113), .B1(new_n1115), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1093), .B1(new_n1123), .B2(new_n794), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(new_n777), .B2(new_n1044), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1083), .A2(new_n1125), .ZN(G393));
  INV_X1    g0926(.A(KEYINPUT114), .ZN(new_n1127));
  AND3_X1   g0927(.A1(new_n1030), .A2(new_n1038), .A3(new_n737), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n737), .B1(new_n1030), .B2(new_n1038), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1127), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1041), .A2(KEYINPUT114), .A3(new_n1047), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1130), .A2(new_n1131), .A3(new_n777), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1045), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1133), .A2(new_n1048), .A3(new_n739), .ZN(new_n1134));
  OAI221_X1 g0934(.A(new_n795), .B1(new_n302), .B2(new_n223), .C1(new_n248), .C2(new_n1051), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n778), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n1136), .B(KEYINPUT115), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(G68), .A2(new_n883), .B1(new_n820), .B2(G143), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1138), .B(new_n334), .C1(new_n609), .C2(new_n808), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT116), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n831), .A2(new_n333), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(new_n352), .B2(new_n866), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1142), .B1(new_n201), .B2(new_n822), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n802), .A2(new_n868), .B1(new_n1114), .B2(new_n828), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT51), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n802), .A2(new_n824), .B1(new_n816), .B2(new_n828), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1147), .B(KEYINPUT52), .ZN(new_n1148));
  OAI221_X1 g0948(.A(new_n459), .B1(new_n533), .B2(new_n808), .C1(new_n822), .C2(new_n813), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n883), .A2(new_n879), .B1(new_n866), .B2(G294), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n829), .B2(new_n819), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n1149), .B(new_n1151), .C1(G116), .C2(new_n832), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n1144), .A2(new_n1146), .B1(new_n1148), .B2(new_n1152), .ZN(new_n1153));
  OAI221_X1 g0953(.A(new_n1137), .B1(new_n1075), .B2(new_n1153), .C1(new_n1031), .C2(new_n1078), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1132), .A2(new_n1134), .A3(new_n1154), .ZN(G390));
  NAND4_X1  g0955(.A1(new_n768), .A2(G330), .A3(new_n913), .A4(new_n861), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n858), .B1(new_n751), .B2(new_n861), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n913), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n946), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n954), .B1(new_n959), .B2(KEYINPUT39), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT117), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n978), .A2(new_n946), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n749), .A2(new_n861), .A3(new_n715), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1159), .B1(new_n1164), .B2(new_n854), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1162), .B1(new_n1163), .B2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n953), .B1(new_n944), .B2(new_n928), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n716), .B1(new_n683), .B2(new_n748), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n858), .B1(new_n1168), .B2(new_n861), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1167), .B(KEYINPUT117), .C1(new_n1169), .C2(new_n1159), .ZN(new_n1170));
  AOI221_X4 g0970(.A(new_n1157), .B1(new_n1160), .B2(new_n1161), .C1(new_n1166), .C2(new_n1170), .ZN(new_n1171));
  AND3_X1   g0971(.A1(new_n763), .A2(new_n716), .A3(new_n969), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n969), .B1(new_n763), .B2(new_n716), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n729), .B1(new_n1174), .B2(new_n753), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(new_n988), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1166), .A2(new_n1170), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1176), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1171), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n768), .A2(G330), .A3(new_n861), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n1159), .A2(new_n1181), .B1(new_n1175), .B2(new_n988), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1169), .A2(new_n1156), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n913), .B1(new_n1175), .B2(new_n861), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n1182), .A2(new_n1158), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1175), .A2(new_n514), .ZN(new_n1186));
  AND3_X1   g0986(.A1(new_n964), .A2(new_n709), .A3(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(KEYINPUT118), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT118), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1185), .A2(new_n1190), .A3(new_n1187), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1189), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1180), .A2(new_n1192), .ZN(new_n1193));
  AND3_X1   g0993(.A1(new_n1185), .A2(new_n1190), .A3(new_n1187), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1190), .B1(new_n1185), .B2(new_n1187), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1177), .A2(new_n1178), .A3(new_n1156), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n1166), .A2(new_n1170), .B1(new_n1161), .B2(new_n1160), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1197), .B1(new_n1198), .B2(new_n1176), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1196), .A2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1193), .A2(new_n1200), .A3(new_n739), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1161), .A2(new_n781), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n459), .B1(new_n812), .B2(new_n609), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1141), .B(new_n1203), .C1(G107), .C2(new_n823), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n828), .A2(new_n298), .B1(new_n808), .B2(new_n377), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n815), .A2(new_n302), .B1(new_n819), .B2(new_n1069), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1204), .B(new_n1207), .C1(new_n809), .C2(new_n802), .ZN(new_n1208));
  INV_X1    g1008(.A(G125), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n334), .B1(new_n1209), .B2(new_n819), .C1(new_n822), .C2(new_n869), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(G159), .B2(new_n832), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n812), .A2(new_n868), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(KEYINPUT119), .B(KEYINPUT53), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1212), .B(new_n1213), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(KEYINPUT54), .B(G143), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n201), .A2(new_n808), .B1(new_n815), .B2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(G132), .B2(new_n865), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1211), .A2(new_n1214), .A3(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(G128), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n802), .A2(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1208), .B1(new_n1218), .B2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(new_n794), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n779), .B1(new_n351), .B2(new_n890), .ZN(new_n1223));
  AND2_X1   g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n1180), .A2(new_n777), .B1(new_n1202), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1201), .A2(new_n1225), .ZN(G378));
  NAND2_X1  g1026(.A1(new_n362), .A2(new_n714), .ZN(new_n1227));
  XNOR2_X1  g1027(.A(new_n1227), .B(KEYINPUT121), .ZN(new_n1228));
  OR2_X1    g1028(.A1(new_n375), .A2(new_n1228), .ZN(new_n1229));
  XOR2_X1   g1029(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1230));
  NAND2_X1  g1030(.A1(new_n375), .A2(new_n1228), .ZN(new_n1231));
  AND3_X1   g1031(.A1(new_n1229), .A2(new_n1230), .A3(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1230), .B1(new_n1229), .B2(new_n1231), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(new_n994), .B2(G330), .ZN(new_n1236));
  AOI211_X1 g1036(.A(new_n729), .B(new_n1234), .C1(new_n990), .C2(new_n993), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n962), .B(new_n952), .C1(new_n1236), .C2(new_n1237), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1234), .B1(new_n980), .B2(new_n729), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n994), .A2(G330), .A3(new_n1235), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n963), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1238), .A2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1234), .A2(new_n781), .ZN(new_n1243));
  AND2_X1   g1043(.A1(new_n890), .A2(new_n201), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(G33), .A2(G41), .ZN(new_n1245));
  AOI211_X1 g1045(.A(G50), .B(new_n1245), .C1(new_n459), .C2(new_n250), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n812), .A2(new_n333), .B1(new_n808), .B2(new_n835), .ZN(new_n1247));
  AOI211_X1 g1047(.A(new_n1053), .B(new_n1247), .C1(G97), .C2(new_n823), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n828), .A2(new_n533), .B1(new_n819), .B2(new_n809), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n250), .B(new_n459), .C1(new_n815), .C2(new_n431), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1248), .B(new_n1251), .C1(new_n298), .C2(new_n802), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT58), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1246), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n822), .A2(new_n875), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n812), .A2(new_n1215), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT120), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  AOI211_X1 g1058(.A(new_n1255), .B(new_n1258), .C1(G150), .C2(new_n832), .ZN(new_n1259));
  OAI22_X1  g1059(.A1(new_n828), .A2(new_n1219), .B1(new_n815), .B2(new_n869), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(new_n1257), .B2(new_n1256), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n1259), .B(new_n1261), .C1(new_n1209), .C2(new_n802), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(KEYINPUT59), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1245), .B1(new_n808), .B2(new_n1114), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1264), .B1(G124), .B2(new_n820), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1263), .A2(new_n1265), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1262), .A2(KEYINPUT59), .ZN(new_n1267));
  OAI221_X1 g1067(.A(new_n1254), .B1(new_n1253), .B2(new_n1252), .C1(new_n1266), .C2(new_n1267), .ZN(new_n1268));
  AOI211_X1 g1068(.A(new_n779), .B(new_n1244), .C1(new_n1268), .C2(new_n794), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(new_n1242), .A2(new_n777), .B1(new_n1243), .B2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1242), .A2(KEYINPUT57), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1187), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1272), .B1(new_n1180), .B2(new_n1192), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n739), .B1(new_n1271), .B2(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1187), .B1(new_n1196), .B2(new_n1199), .ZN(new_n1275));
  AOI21_X1  g1075(.A(KEYINPUT57), .B1(new_n1275), .B2(new_n1242), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1270), .B1(new_n1274), .B2(new_n1276), .ZN(G375));
  AOI21_X1  g1077(.A(new_n779), .B1(new_n377), .B2(new_n890), .ZN(new_n1278));
  OAI221_X1 g1078(.A(new_n334), .B1(new_n835), .B2(new_n808), .C1(new_n822), .C2(new_n1215), .ZN(new_n1279));
  AOI22_X1  g1079(.A1(G159), .A2(new_n883), .B1(new_n820), .B2(G128), .ZN(new_n1280));
  OAI221_X1 g1080(.A(new_n1280), .B1(new_n869), .B2(new_n828), .C1(new_n868), .C2(new_n815), .ZN(new_n1281));
  AOI211_X1 g1081(.A(new_n1279), .B(new_n1281), .C1(G50), .C2(new_n832), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n803), .A2(G132), .ZN(new_n1283));
  AOI22_X1  g1083(.A1(new_n823), .A2(G116), .B1(G107), .B2(new_n866), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1284), .B1(new_n802), .B2(new_n1069), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(new_n1285), .B(KEYINPUT123), .ZN(new_n1286));
  AOI22_X1  g1086(.A1(G97), .A2(new_n883), .B1(new_n865), .B2(G283), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1287), .B1(new_n813), .B2(new_n819), .ZN(new_n1288));
  NOR4_X1   g1088(.A1(new_n1288), .A2(new_n334), .A3(new_n1058), .A4(new_n1120), .ZN(new_n1289));
  AOI22_X1  g1089(.A1(new_n1282), .A2(new_n1283), .B1(new_n1286), .B2(new_n1289), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1278), .B1(new_n1290), .B2(new_n1075), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1291), .B1(new_n1159), .B2(new_n781), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1292), .B1(new_n1185), .B2(new_n777), .ZN(new_n1293));
  OR2_X1    g1093(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1189), .A2(new_n1191), .A3(new_n1294), .ZN(new_n1295));
  XNOR2_X1  g1095(.A(new_n1024), .B(KEYINPUT122), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1293), .B1(new_n1295), .B2(new_n1296), .ZN(G381));
  XNOR2_X1  g1097(.A(G375), .B(KEYINPUT124), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1083), .A2(new_n1125), .A3(new_n849), .ZN(new_n1299));
  OR4_X1    g1099(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1299), .ZN(new_n1300));
  OR4_X1    g1100(.A1(G387), .A2(new_n1298), .A3(G378), .A4(new_n1300), .ZN(G407));
  INV_X1    g1101(.A(G213), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1302), .A2(G343), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1303), .ZN(new_n1304));
  OR3_X1    g1104(.A1(new_n1298), .A2(G378), .A3(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(G407), .A2(new_n1305), .A3(G213), .ZN(G409));
  OAI211_X1 g1106(.A(G378), .B(new_n1270), .C1(new_n1274), .C2(new_n1276), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1275), .A2(new_n1242), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1270), .B1(new_n1308), .B2(new_n1296), .ZN(new_n1309));
  AND2_X1   g1109(.A1(new_n1201), .A2(new_n1225), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1307), .A2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(new_n1304), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1295), .A2(KEYINPUT60), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT60), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1315), .B1(new_n1185), .B2(new_n1187), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(new_n739), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(KEYINPUT125), .B1(new_n1314), .B2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT125), .ZN(new_n1320));
  AOI211_X1 g1120(.A(new_n1320), .B(new_n1317), .C1(new_n1295), .C2(KEYINPUT60), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1293), .B1(new_n1319), .B2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1322), .A2(new_n893), .ZN(new_n1323));
  OAI211_X1 g1123(.A(G384), .B(new_n1293), .C1(new_n1319), .C2(new_n1321), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  OAI21_X1  g1125(.A(KEYINPUT62), .B1(new_n1313), .B2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1303), .A2(G2897), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1323), .A2(new_n1324), .A3(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1327), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1330));
  NOR3_X1   g1130(.A1(new_n1194), .A2(new_n1195), .A3(new_n1330), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1318), .B1(new_n1331), .B2(new_n1315), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1332), .A2(new_n1320), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1314), .A2(KEYINPUT125), .A3(new_n1318), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  AOI21_X1  g1135(.A(G384), .B1(new_n1335), .B2(new_n1293), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1324), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1329), .B1(new_n1336), .B2(new_n1337), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1313), .A2(new_n1328), .A3(new_n1338), .ZN(new_n1339));
  INV_X1    g1139(.A(KEYINPUT61), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1303), .B1(new_n1307), .B2(new_n1311), .ZN(new_n1341));
  NOR2_X1   g1141(.A1(new_n1336), .A2(new_n1337), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT62), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1341), .A2(new_n1342), .A3(new_n1343), .ZN(new_n1344));
  NAND4_X1  g1144(.A1(new_n1326), .A2(new_n1339), .A3(new_n1340), .A4(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(G393), .A2(G396), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1346), .A2(new_n1299), .ZN(new_n1347));
  INV_X1    g1147(.A(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(G390), .A2(new_n1348), .ZN(new_n1349));
  NAND4_X1  g1149(.A1(new_n1347), .A2(new_n1132), .A3(new_n1134), .A4(new_n1154), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1349), .A2(new_n1350), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1351), .A2(G387), .ZN(new_n1352));
  NAND4_X1  g1152(.A1(new_n1349), .A2(new_n1050), .A3(new_n1079), .A4(new_n1350), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1352), .A2(new_n1353), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1345), .A2(new_n1354), .ZN(new_n1355));
  AND3_X1   g1155(.A1(new_n1341), .A2(new_n1342), .A3(KEYINPUT63), .ZN(new_n1356));
  AOI21_X1  g1156(.A(KEYINPUT63), .B1(new_n1341), .B2(new_n1342), .ZN(new_n1357));
  NOR2_X1   g1157(.A1(new_n1356), .A2(new_n1357), .ZN(new_n1358));
  AND3_X1   g1158(.A1(new_n1323), .A2(new_n1324), .A3(new_n1327), .ZN(new_n1359));
  AOI21_X1  g1159(.A(new_n1327), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1360));
  NOR2_X1   g1160(.A1(new_n1359), .A2(new_n1360), .ZN(new_n1361));
  AOI21_X1  g1161(.A(KEYINPUT61), .B1(new_n1361), .B2(new_n1313), .ZN(new_n1362));
  INV_X1    g1162(.A(new_n1354), .ZN(new_n1363));
  NAND3_X1  g1163(.A1(new_n1358), .A2(new_n1362), .A3(new_n1363), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1355), .A2(new_n1364), .ZN(G405));
  AND3_X1   g1165(.A1(new_n1352), .A2(KEYINPUT127), .A3(new_n1353), .ZN(new_n1366));
  INV_X1    g1166(.A(new_n1307), .ZN(new_n1367));
  NAND3_X1  g1167(.A1(new_n1275), .A2(KEYINPUT57), .A3(new_n1242), .ZN(new_n1368));
  AOI22_X1  g1168(.A1(new_n1193), .A2(new_n1187), .B1(new_n1241), .B2(new_n1238), .ZN(new_n1369));
  OAI211_X1 g1169(.A(new_n739), .B(new_n1368), .C1(new_n1369), .C2(KEYINPUT57), .ZN(new_n1370));
  AOI21_X1  g1170(.A(G378), .B1(new_n1370), .B2(new_n1270), .ZN(new_n1371));
  NOR2_X1   g1171(.A1(new_n1367), .A2(new_n1371), .ZN(new_n1372));
  AOI21_X1  g1172(.A(new_n1366), .B1(new_n1372), .B2(new_n1325), .ZN(new_n1373));
  NAND2_X1  g1173(.A1(G375), .A2(new_n1310), .ZN(new_n1374));
  NAND2_X1  g1174(.A1(new_n1374), .A2(new_n1307), .ZN(new_n1375));
  INV_X1    g1175(.A(KEYINPUT126), .ZN(new_n1376));
  AND3_X1   g1176(.A1(new_n1375), .A2(new_n1376), .A3(new_n1342), .ZN(new_n1377));
  AOI21_X1  g1177(.A(new_n1376), .B1(new_n1375), .B2(new_n1342), .ZN(new_n1378));
  OAI21_X1  g1178(.A(new_n1373), .B1(new_n1377), .B2(new_n1378), .ZN(new_n1379));
  NOR2_X1   g1179(.A1(new_n1363), .A2(KEYINPUT127), .ZN(new_n1380));
  NAND2_X1  g1180(.A1(new_n1379), .A2(new_n1380), .ZN(new_n1381));
  OAI221_X1 g1181(.A(new_n1373), .B1(KEYINPUT127), .B2(new_n1363), .C1(new_n1377), .C2(new_n1378), .ZN(new_n1382));
  NAND2_X1  g1182(.A1(new_n1381), .A2(new_n1382), .ZN(G402));
endmodule


