

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U555 ( .A(G2104), .ZN(n536) );
  NOR2_X1 U556 ( .A1(n697), .A2(n963), .ZN(n705) );
  INV_X1 U557 ( .A(n699), .ZN(n735) );
  AND2_X1 U558 ( .A1(n539), .A2(n538), .ZN(G164) );
  AND2_X2 U559 ( .A1(n693), .A2(n778), .ZN(n699) );
  NOR2_X2 U560 ( .A1(n537), .A2(n536), .ZN(n887) );
  NOR2_X2 U561 ( .A1(n650), .A2(n544), .ZN(n654) );
  NOR2_X1 U562 ( .A1(n764), .A2(n765), .ZN(n766) );
  XNOR2_X1 U563 ( .A(n563), .B(n562), .ZN(n564) );
  NAND2_X1 U564 ( .A1(n699), .A2(G1996), .ZN(n694) );
  INV_X1 U565 ( .A(KEYINPUT103), .ZN(n761) );
  INV_X1 U566 ( .A(n947), .ZN(n765) );
  INV_X1 U567 ( .A(G2105), .ZN(n530) );
  NAND2_X1 U568 ( .A1(n814), .A2(n813), .ZN(n815) );
  NOR2_X1 U569 ( .A1(n812), .A2(n525), .ZN(n813) );
  XNOR2_X1 U570 ( .A(n567), .B(n566), .ZN(n963) );
  INV_X1 U571 ( .A(KEYINPUT68), .ZN(n566) );
  NOR2_X1 U572 ( .A1(n565), .A2(n564), .ZN(n567) );
  XNOR2_X1 U573 ( .A(KEYINPUT26), .B(KEYINPUT96), .ZN(n523) );
  AND2_X1 U574 ( .A1(G114), .A2(n887), .ZN(n524) );
  AND2_X1 U575 ( .A1(n827), .A2(n960), .ZN(n525) );
  OR2_X1 U576 ( .A1(n774), .A2(n773), .ZN(n526) );
  AND2_X1 U577 ( .A1(n775), .A2(n526), .ZN(n527) );
  NOR2_X1 U578 ( .A1(n774), .A2(n757), .ZN(n528) );
  XNOR2_X1 U579 ( .A(n694), .B(n523), .ZN(n696) );
  INV_X1 U580 ( .A(KEYINPUT32), .ZN(n743) );
  INV_X1 U581 ( .A(G2104), .ZN(n529) );
  NOR2_X2 U582 ( .A1(G164), .A2(G1384), .ZN(n778) );
  NAND2_X1 U583 ( .A1(n657), .A2(G56), .ZN(n556) );
  XNOR2_X1 U584 ( .A(n531), .B(KEYINPUT17), .ZN(n549) );
  NOR2_X1 U585 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U586 ( .A(KEYINPUT67), .B(KEYINPUT13), .ZN(n562) );
  INV_X1 U587 ( .A(KEYINPUT1), .ZN(n540) );
  NOR2_X2 U588 ( .A1(G2104), .A2(n537), .ZN(n888) );
  XNOR2_X1 U589 ( .A(n815), .B(KEYINPUT104), .ZN(n830) );
  NOR2_X1 U590 ( .A1(n535), .A2(n524), .ZN(n539) );
  NAND2_X1 U591 ( .A1(n530), .A2(n529), .ZN(n531) );
  NAND2_X1 U592 ( .A1(G138), .A2(n549), .ZN(n533) );
  NOR2_X4 U593 ( .A1(G2105), .A2(n536), .ZN(n895) );
  NAND2_X1 U594 ( .A1(G102), .A2(n895), .ZN(n532) );
  NAND2_X1 U595 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U596 ( .A(n534), .B(KEYINPUT84), .ZN(n535) );
  INV_X1 U597 ( .A(G2105), .ZN(n537) );
  NAND2_X1 U598 ( .A1(G126), .A2(n888), .ZN(n538) );
  INV_X1 U599 ( .A(G651), .ZN(n544) );
  NOR2_X1 U600 ( .A1(G543), .A2(n544), .ZN(n541) );
  XNOR2_X2 U601 ( .A(n541), .B(n540), .ZN(n657) );
  NAND2_X1 U602 ( .A1(G60), .A2(n657), .ZN(n543) );
  XOR2_X1 U603 ( .A(KEYINPUT0), .B(G543), .Z(n650) );
  NOR2_X2 U604 ( .A1(G651), .A2(n650), .ZN(n658) );
  NAND2_X1 U605 ( .A1(G47), .A2(n658), .ZN(n542) );
  NAND2_X1 U606 ( .A1(n543), .A2(n542), .ZN(n548) );
  NOR2_X2 U607 ( .A1(G651), .A2(G543), .ZN(n653) );
  NAND2_X1 U608 ( .A1(G85), .A2(n653), .ZN(n546) );
  NAND2_X1 U609 ( .A1(G72), .A2(n654), .ZN(n545) );
  NAND2_X1 U610 ( .A1(n546), .A2(n545), .ZN(n547) );
  OR2_X1 U611 ( .A1(n548), .A2(n547), .ZN(G290) );
  INV_X1 U612 ( .A(n549), .ZN(n550) );
  INV_X1 U613 ( .A(n550), .ZN(n892) );
  NAND2_X1 U614 ( .A1(n892), .A2(G137), .ZN(n553) );
  NAND2_X1 U615 ( .A1(G101), .A2(n895), .ZN(n551) );
  XOR2_X1 U616 ( .A(KEYINPUT23), .B(n551), .Z(n552) );
  AND2_X1 U617 ( .A1(n553), .A2(n552), .ZN(n690) );
  NAND2_X1 U618 ( .A1(G113), .A2(n887), .ZN(n555) );
  NAND2_X1 U619 ( .A1(G125), .A2(n888), .ZN(n554) );
  AND2_X1 U620 ( .A1(n555), .A2(n554), .ZN(n689) );
  AND2_X1 U621 ( .A1(n690), .A2(n689), .ZN(G160) );
  AND2_X1 U622 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U623 ( .A(G860), .ZN(n614) );
  XNOR2_X1 U624 ( .A(n556), .B(KEYINPUT14), .ZN(n558) );
  NAND2_X1 U625 ( .A1(G43), .A2(n658), .ZN(n557) );
  NAND2_X1 U626 ( .A1(n558), .A2(n557), .ZN(n565) );
  NAND2_X1 U627 ( .A1(n653), .A2(G81), .ZN(n559) );
  XNOR2_X1 U628 ( .A(n559), .B(KEYINPUT12), .ZN(n561) );
  NAND2_X1 U629 ( .A1(G68), .A2(n654), .ZN(n560) );
  NAND2_X1 U630 ( .A1(n561), .A2(n560), .ZN(n563) );
  OR2_X1 U631 ( .A1(n614), .A2(n963), .ZN(G153) );
  INV_X1 U632 ( .A(G57), .ZN(G237) );
  INV_X1 U633 ( .A(G132), .ZN(G219) );
  INV_X1 U634 ( .A(G82), .ZN(G220) );
  NAND2_X1 U635 ( .A1(G65), .A2(n657), .ZN(n569) );
  NAND2_X1 U636 ( .A1(G53), .A2(n658), .ZN(n568) );
  NAND2_X1 U637 ( .A1(n569), .A2(n568), .ZN(n573) );
  NAND2_X1 U638 ( .A1(G91), .A2(n653), .ZN(n571) );
  NAND2_X1 U639 ( .A1(G78), .A2(n654), .ZN(n570) );
  NAND2_X1 U640 ( .A1(n571), .A2(n570), .ZN(n572) );
  NOR2_X1 U641 ( .A1(n573), .A2(n572), .ZN(n714) );
  INV_X1 U642 ( .A(n714), .ZN(G299) );
  NAND2_X1 U643 ( .A1(G64), .A2(n657), .ZN(n575) );
  NAND2_X1 U644 ( .A1(G52), .A2(n658), .ZN(n574) );
  NAND2_X1 U645 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U646 ( .A(KEYINPUT64), .B(n576), .ZN(n582) );
  NAND2_X1 U647 ( .A1(n653), .A2(G90), .ZN(n577) );
  XOR2_X1 U648 ( .A(KEYINPUT65), .B(n577), .Z(n579) );
  NAND2_X1 U649 ( .A1(n654), .A2(G77), .ZN(n578) );
  NAND2_X1 U650 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U651 ( .A(KEYINPUT9), .B(n580), .Z(n581) );
  NOR2_X1 U652 ( .A1(n582), .A2(n581), .ZN(G171) );
  NAND2_X1 U653 ( .A1(G63), .A2(n657), .ZN(n584) );
  NAND2_X1 U654 ( .A1(G51), .A2(n658), .ZN(n583) );
  NAND2_X1 U655 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U656 ( .A(KEYINPUT6), .B(n585), .ZN(n594) );
  NAND2_X1 U657 ( .A1(G76), .A2(n654), .ZN(n590) );
  XOR2_X1 U658 ( .A(KEYINPUT4), .B(KEYINPUT74), .Z(n587) );
  NAND2_X1 U659 ( .A1(G89), .A2(n653), .ZN(n586) );
  XNOR2_X1 U660 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U661 ( .A(KEYINPUT73), .B(n588), .ZN(n589) );
  NAND2_X1 U662 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U663 ( .A(n591), .B(KEYINPUT75), .ZN(n592) );
  XNOR2_X1 U664 ( .A(n592), .B(KEYINPUT5), .ZN(n593) );
  NOR2_X1 U665 ( .A1(n594), .A2(n593), .ZN(n595) );
  XOR2_X1 U666 ( .A(KEYINPUT7), .B(n595), .Z(G168) );
  XOR2_X1 U667 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U668 ( .A1(G7), .A2(G661), .ZN(n596) );
  XNOR2_X1 U669 ( .A(n596), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U670 ( .A(G223), .B(KEYINPUT66), .Z(n832) );
  NAND2_X1 U671 ( .A1(n832), .A2(G567), .ZN(n597) );
  XOR2_X1 U672 ( .A(KEYINPUT11), .B(n597), .Z(G234) );
  INV_X1 U673 ( .A(G171), .ZN(G301) );
  NAND2_X1 U674 ( .A1(G66), .A2(n657), .ZN(n599) );
  NAND2_X1 U675 ( .A1(G92), .A2(n653), .ZN(n598) );
  NAND2_X1 U676 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U677 ( .A(KEYINPUT69), .B(n600), .ZN(n606) );
  NAND2_X1 U678 ( .A1(G54), .A2(n658), .ZN(n601) );
  XNOR2_X1 U679 ( .A(n601), .B(KEYINPUT71), .ZN(n604) );
  NAND2_X1 U680 ( .A1(G79), .A2(n654), .ZN(n602) );
  XOR2_X1 U681 ( .A(KEYINPUT70), .B(n602), .Z(n603) );
  NAND2_X1 U682 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X2 U683 ( .A(KEYINPUT15), .B(n607), .ZN(n858) );
  INV_X1 U684 ( .A(n858), .ZN(n966) );
  INV_X1 U685 ( .A(G868), .ZN(n611) );
  NAND2_X1 U686 ( .A1(n966), .A2(n611), .ZN(n608) );
  XNOR2_X1 U687 ( .A(n608), .B(KEYINPUT72), .ZN(n610) );
  NAND2_X1 U688 ( .A1(G868), .A2(G301), .ZN(n609) );
  NAND2_X1 U689 ( .A1(n610), .A2(n609), .ZN(G284) );
  NOR2_X1 U690 ( .A1(G286), .A2(n611), .ZN(n613) );
  NOR2_X1 U691 ( .A1(G868), .A2(G299), .ZN(n612) );
  NOR2_X1 U692 ( .A1(n613), .A2(n612), .ZN(G297) );
  NAND2_X1 U693 ( .A1(n614), .A2(G559), .ZN(n615) );
  NAND2_X1 U694 ( .A1(n615), .A2(n858), .ZN(n616) );
  XNOR2_X1 U695 ( .A(n616), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U696 ( .A1(n858), .A2(G868), .ZN(n617) );
  NOR2_X1 U697 ( .A1(G559), .A2(n617), .ZN(n618) );
  XNOR2_X1 U698 ( .A(n618), .B(KEYINPUT76), .ZN(n620) );
  NOR2_X1 U699 ( .A1(n963), .A2(G868), .ZN(n619) );
  NOR2_X1 U700 ( .A1(n620), .A2(n619), .ZN(G282) );
  NAND2_X1 U701 ( .A1(G135), .A2(n892), .ZN(n622) );
  NAND2_X1 U702 ( .A1(G111), .A2(n887), .ZN(n621) );
  NAND2_X1 U703 ( .A1(n622), .A2(n621), .ZN(n625) );
  NAND2_X1 U704 ( .A1(n888), .A2(G123), .ZN(n623) );
  XOR2_X1 U705 ( .A(KEYINPUT18), .B(n623), .Z(n624) );
  NOR2_X1 U706 ( .A1(n625), .A2(n624), .ZN(n627) );
  NAND2_X1 U707 ( .A1(n895), .A2(G99), .ZN(n626) );
  NAND2_X1 U708 ( .A1(n627), .A2(n626), .ZN(n1008) );
  XOR2_X1 U709 ( .A(G2096), .B(KEYINPUT77), .Z(n628) );
  XNOR2_X1 U710 ( .A(n1008), .B(n628), .ZN(n629) );
  NOR2_X1 U711 ( .A1(G2100), .A2(n629), .ZN(n630) );
  XOR2_X1 U712 ( .A(KEYINPUT78), .B(n630), .Z(G156) );
  NAND2_X1 U713 ( .A1(G559), .A2(n858), .ZN(n631) );
  XNOR2_X1 U714 ( .A(n631), .B(n963), .ZN(n669) );
  NOR2_X1 U715 ( .A1(G860), .A2(n669), .ZN(n639) );
  NAND2_X1 U716 ( .A1(G67), .A2(n657), .ZN(n633) );
  NAND2_X1 U717 ( .A1(G55), .A2(n658), .ZN(n632) );
  NAND2_X1 U718 ( .A1(n633), .A2(n632), .ZN(n636) );
  NAND2_X1 U719 ( .A1(G80), .A2(n654), .ZN(n634) );
  XNOR2_X1 U720 ( .A(KEYINPUT79), .B(n634), .ZN(n635) );
  NOR2_X1 U721 ( .A1(n636), .A2(n635), .ZN(n638) );
  NAND2_X1 U722 ( .A1(n653), .A2(G93), .ZN(n637) );
  NAND2_X1 U723 ( .A1(n638), .A2(n637), .ZN(n668) );
  XOR2_X1 U724 ( .A(n639), .B(n668), .Z(G145) );
  NAND2_X1 U725 ( .A1(G61), .A2(n657), .ZN(n641) );
  NAND2_X1 U726 ( .A1(G48), .A2(n658), .ZN(n640) );
  NAND2_X1 U727 ( .A1(n641), .A2(n640), .ZN(n644) );
  NAND2_X1 U728 ( .A1(n654), .A2(G73), .ZN(n642) );
  XOR2_X1 U729 ( .A(KEYINPUT2), .B(n642), .Z(n643) );
  NOR2_X1 U730 ( .A1(n644), .A2(n643), .ZN(n646) );
  NAND2_X1 U731 ( .A1(n653), .A2(G86), .ZN(n645) );
  NAND2_X1 U732 ( .A1(n646), .A2(n645), .ZN(G305) );
  NAND2_X1 U733 ( .A1(G49), .A2(n658), .ZN(n648) );
  NAND2_X1 U734 ( .A1(G74), .A2(G651), .ZN(n647) );
  NAND2_X1 U735 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U736 ( .A1(n657), .A2(n649), .ZN(n652) );
  NAND2_X1 U737 ( .A1(n650), .A2(G87), .ZN(n651) );
  NAND2_X1 U738 ( .A1(n652), .A2(n651), .ZN(G288) );
  NAND2_X1 U739 ( .A1(G88), .A2(n653), .ZN(n656) );
  NAND2_X1 U740 ( .A1(G75), .A2(n654), .ZN(n655) );
  NAND2_X1 U741 ( .A1(n656), .A2(n655), .ZN(n662) );
  NAND2_X1 U742 ( .A1(G62), .A2(n657), .ZN(n660) );
  NAND2_X1 U743 ( .A1(G50), .A2(n658), .ZN(n659) );
  NAND2_X1 U744 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U745 ( .A1(n662), .A2(n661), .ZN(G166) );
  OR2_X1 U746 ( .A1(G868), .A2(n668), .ZN(n673) );
  XNOR2_X1 U747 ( .A(G288), .B(KEYINPUT19), .ZN(n664) );
  XNOR2_X1 U748 ( .A(G166), .B(n714), .ZN(n663) );
  XNOR2_X1 U749 ( .A(n664), .B(n663), .ZN(n665) );
  XOR2_X1 U750 ( .A(n665), .B(G290), .Z(n666) );
  XNOR2_X1 U751 ( .A(G305), .B(n666), .ZN(n667) );
  XOR2_X1 U752 ( .A(n668), .B(n667), .Z(n857) );
  XNOR2_X1 U753 ( .A(n669), .B(n857), .ZN(n670) );
  XNOR2_X1 U754 ( .A(n670), .B(KEYINPUT80), .ZN(n671) );
  NAND2_X1 U755 ( .A1(n671), .A2(G868), .ZN(n672) );
  NAND2_X1 U756 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U757 ( .A(n674), .B(KEYINPUT81), .ZN(G295) );
  NAND2_X1 U758 ( .A1(G2078), .A2(G2084), .ZN(n675) );
  XOR2_X1 U759 ( .A(KEYINPUT20), .B(n675), .Z(n676) );
  NAND2_X1 U760 ( .A1(G2090), .A2(n676), .ZN(n677) );
  XNOR2_X1 U761 ( .A(KEYINPUT21), .B(n677), .ZN(n678) );
  NAND2_X1 U762 ( .A1(n678), .A2(G2072), .ZN(n679) );
  XNOR2_X1 U763 ( .A(KEYINPUT82), .B(n679), .ZN(G158) );
  XNOR2_X1 U764 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U765 ( .A1(G220), .A2(G219), .ZN(n680) );
  XNOR2_X1 U766 ( .A(KEYINPUT22), .B(n680), .ZN(n681) );
  NAND2_X1 U767 ( .A1(n681), .A2(G96), .ZN(n682) );
  NOR2_X1 U768 ( .A1(n682), .A2(G218), .ZN(n683) );
  XNOR2_X1 U769 ( .A(n683), .B(KEYINPUT83), .ZN(n836) );
  NAND2_X1 U770 ( .A1(n836), .A2(G2106), .ZN(n687) );
  NAND2_X1 U771 ( .A1(G69), .A2(G120), .ZN(n684) );
  NOR2_X1 U772 ( .A1(G237), .A2(n684), .ZN(n685) );
  NAND2_X1 U773 ( .A1(G108), .A2(n685), .ZN(n837) );
  NAND2_X1 U774 ( .A1(n837), .A2(G567), .ZN(n686) );
  NAND2_X1 U775 ( .A1(n687), .A2(n686), .ZN(n838) );
  NAND2_X1 U776 ( .A1(G483), .A2(G661), .ZN(n688) );
  NOR2_X1 U777 ( .A1(n838), .A2(n688), .ZN(n835) );
  NAND2_X1 U778 ( .A1(n835), .A2(G36), .ZN(G176) );
  INV_X1 U779 ( .A(G166), .ZN(G303) );
  AND2_X1 U780 ( .A1(G40), .A2(n689), .ZN(n691) );
  NAND2_X1 U781 ( .A1(n691), .A2(n690), .ZN(n777) );
  INV_X1 U782 ( .A(n777), .ZN(n693) );
  NAND2_X1 U783 ( .A1(n735), .A2(G1341), .ZN(n695) );
  NAND2_X1 U784 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U785 ( .A1(n705), .A2(n858), .ZN(n703) );
  AND2_X1 U786 ( .A1(n735), .A2(G1348), .ZN(n698) );
  XNOR2_X1 U787 ( .A(n698), .B(KEYINPUT97), .ZN(n701) );
  NAND2_X1 U788 ( .A1(n699), .A2(G2067), .ZN(n700) );
  NAND2_X1 U789 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U790 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U791 ( .A(n704), .B(KEYINPUT98), .ZN(n707) );
  OR2_X1 U792 ( .A1(n858), .A2(n705), .ZN(n706) );
  NAND2_X1 U793 ( .A1(n707), .A2(n706), .ZN(n712) );
  NAND2_X1 U794 ( .A1(n699), .A2(G2072), .ZN(n708) );
  XNOR2_X1 U795 ( .A(n708), .B(KEYINPUT27), .ZN(n710) );
  XNOR2_X1 U796 ( .A(G1956), .B(KEYINPUT95), .ZN(n988) );
  NOR2_X1 U797 ( .A1(n988), .A2(n699), .ZN(n709) );
  NOR2_X1 U798 ( .A1(n710), .A2(n709), .ZN(n713) );
  NAND2_X1 U799 ( .A1(n714), .A2(n713), .ZN(n711) );
  NAND2_X1 U800 ( .A1(n712), .A2(n711), .ZN(n717) );
  NOR2_X1 U801 ( .A1(n714), .A2(n713), .ZN(n715) );
  XOR2_X1 U802 ( .A(n715), .B(KEYINPUT28), .Z(n716) );
  NAND2_X1 U803 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U804 ( .A(KEYINPUT29), .B(n718), .ZN(n724) );
  XNOR2_X1 U805 ( .A(G2078), .B(KEYINPUT93), .ZN(n719) );
  XNOR2_X1 U806 ( .A(n719), .B(KEYINPUT25), .ZN(n931) );
  NOR2_X1 U807 ( .A1(n931), .A2(n735), .ZN(n721) );
  NOR2_X1 U808 ( .A1(n699), .A2(G1961), .ZN(n720) );
  NOR2_X1 U809 ( .A1(n721), .A2(n720), .ZN(n728) );
  NOR2_X1 U810 ( .A1(n728), .A2(G301), .ZN(n722) );
  XNOR2_X1 U811 ( .A(n722), .B(KEYINPUT94), .ZN(n723) );
  NOR2_X1 U812 ( .A1(n724), .A2(n723), .ZN(n733) );
  NAND2_X1 U813 ( .A1(G8), .A2(n735), .ZN(n774) );
  NOR2_X1 U814 ( .A1(G1966), .A2(n774), .ZN(n748) );
  NOR2_X1 U815 ( .A1(G2084), .A2(n735), .ZN(n745) );
  NOR2_X1 U816 ( .A1(n748), .A2(n745), .ZN(n725) );
  NAND2_X1 U817 ( .A1(G8), .A2(n725), .ZN(n726) );
  XNOR2_X1 U818 ( .A(KEYINPUT30), .B(n726), .ZN(n727) );
  NOR2_X1 U819 ( .A1(G168), .A2(n727), .ZN(n730) );
  AND2_X1 U820 ( .A1(G301), .A2(n728), .ZN(n729) );
  NOR2_X1 U821 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U822 ( .A(n731), .B(KEYINPUT31), .ZN(n732) );
  NOR2_X1 U823 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U824 ( .A(n734), .B(KEYINPUT99), .ZN(n746) );
  NAND2_X1 U825 ( .A1(n746), .A2(G286), .ZN(n742) );
  INV_X1 U826 ( .A(G8), .ZN(n740) );
  NOR2_X1 U827 ( .A1(G1971), .A2(n774), .ZN(n737) );
  NOR2_X1 U828 ( .A1(G2090), .A2(n735), .ZN(n736) );
  NOR2_X1 U829 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U830 ( .A1(n738), .A2(G303), .ZN(n739) );
  OR2_X1 U831 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U832 ( .A1(n742), .A2(n741), .ZN(n744) );
  XNOR2_X1 U833 ( .A(n744), .B(n743), .ZN(n752) );
  NAND2_X1 U834 ( .A1(G8), .A2(n745), .ZN(n750) );
  INV_X1 U835 ( .A(n746), .ZN(n747) );
  NOR2_X1 U836 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U837 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U838 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U839 ( .A(n753), .B(KEYINPUT100), .ZN(n769) );
  NOR2_X1 U840 ( .A1(G1976), .A2(G288), .ZN(n958) );
  NOR2_X1 U841 ( .A1(G1971), .A2(G303), .ZN(n950) );
  NOR2_X1 U842 ( .A1(n958), .A2(n950), .ZN(n754) );
  XOR2_X1 U843 ( .A(KEYINPUT101), .B(n754), .Z(n755) );
  NAND2_X1 U844 ( .A1(n769), .A2(n755), .ZN(n756) );
  XNOR2_X1 U845 ( .A(n756), .B(KEYINPUT102), .ZN(n758) );
  NAND2_X1 U846 ( .A1(G1976), .A2(G288), .ZN(n952) );
  INV_X1 U847 ( .A(n952), .ZN(n757) );
  NAND2_X1 U848 ( .A1(n758), .A2(n528), .ZN(n760) );
  INV_X1 U849 ( .A(KEYINPUT33), .ZN(n759) );
  NAND2_X1 U850 ( .A1(n760), .A2(n759), .ZN(n762) );
  XNOR2_X1 U851 ( .A(n762), .B(n761), .ZN(n767) );
  NAND2_X1 U852 ( .A1(n958), .A2(KEYINPUT33), .ZN(n763) );
  NOR2_X1 U853 ( .A1(n763), .A2(n774), .ZN(n764) );
  XOR2_X1 U854 ( .A(G1981), .B(G305), .Z(n947) );
  NAND2_X1 U855 ( .A1(n767), .A2(n766), .ZN(n776) );
  NOR2_X1 U856 ( .A1(G2090), .A2(G303), .ZN(n768) );
  NAND2_X1 U857 ( .A1(G8), .A2(n768), .ZN(n770) );
  NAND2_X1 U858 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U859 ( .A1(n771), .A2(n774), .ZN(n775) );
  NOR2_X1 U860 ( .A1(G1981), .A2(G305), .ZN(n772) );
  XOR2_X1 U861 ( .A(n772), .B(KEYINPUT24), .Z(n773) );
  NAND2_X1 U862 ( .A1(n776), .A2(n527), .ZN(n814) );
  NOR2_X1 U863 ( .A1(n778), .A2(n777), .ZN(n779) );
  XOR2_X1 U864 ( .A(KEYINPUT85), .B(n779), .Z(n827) );
  NAND2_X1 U865 ( .A1(G140), .A2(n892), .ZN(n781) );
  NAND2_X1 U866 ( .A1(G104), .A2(n895), .ZN(n780) );
  NAND2_X1 U867 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U868 ( .A(KEYINPUT34), .B(n782), .ZN(n787) );
  NAND2_X1 U869 ( .A1(G116), .A2(n887), .ZN(n784) );
  NAND2_X1 U870 ( .A1(G128), .A2(n888), .ZN(n783) );
  NAND2_X1 U871 ( .A1(n784), .A2(n783), .ZN(n785) );
  XOR2_X1 U872 ( .A(KEYINPUT35), .B(n785), .Z(n786) );
  NOR2_X1 U873 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U874 ( .A(KEYINPUT36), .B(n788), .ZN(n881) );
  XNOR2_X1 U875 ( .A(KEYINPUT37), .B(G2067), .ZN(n825) );
  NOR2_X1 U876 ( .A1(n881), .A2(n825), .ZN(n1015) );
  NAND2_X1 U877 ( .A1(n827), .A2(n1015), .ZN(n823) );
  INV_X1 U878 ( .A(n823), .ZN(n810) );
  XNOR2_X1 U879 ( .A(n827), .B(KEYINPUT90), .ZN(n808) );
  NAND2_X1 U880 ( .A1(G131), .A2(n892), .ZN(n790) );
  NAND2_X1 U881 ( .A1(G107), .A2(n887), .ZN(n789) );
  NAND2_X1 U882 ( .A1(n790), .A2(n789), .ZN(n794) );
  NAND2_X1 U883 ( .A1(G95), .A2(n895), .ZN(n792) );
  NAND2_X1 U884 ( .A1(G119), .A2(n888), .ZN(n791) );
  NAND2_X1 U885 ( .A1(n792), .A2(n791), .ZN(n793) );
  OR2_X1 U886 ( .A1(n794), .A2(n793), .ZN(n903) );
  NAND2_X1 U887 ( .A1(G1991), .A2(n903), .ZN(n795) );
  XNOR2_X1 U888 ( .A(n795), .B(KEYINPUT86), .ZN(n807) );
  NAND2_X1 U889 ( .A1(n888), .A2(G129), .ZN(n796) );
  XOR2_X1 U890 ( .A(KEYINPUT87), .B(n796), .Z(n798) );
  NAND2_X1 U891 ( .A1(n887), .A2(G117), .ZN(n797) );
  NAND2_X1 U892 ( .A1(n798), .A2(n797), .ZN(n799) );
  XNOR2_X1 U893 ( .A(KEYINPUT88), .B(n799), .ZN(n802) );
  NAND2_X1 U894 ( .A1(n895), .A2(G105), .ZN(n800) );
  XOR2_X1 U895 ( .A(KEYINPUT38), .B(n800), .Z(n801) );
  NOR2_X1 U896 ( .A1(n802), .A2(n801), .ZN(n804) );
  NAND2_X1 U897 ( .A1(n892), .A2(G141), .ZN(n803) );
  NAND2_X1 U898 ( .A1(n804), .A2(n803), .ZN(n805) );
  XOR2_X1 U899 ( .A(KEYINPUT89), .B(n805), .Z(n908) );
  NAND2_X1 U900 ( .A1(G1996), .A2(n908), .ZN(n806) );
  NAND2_X1 U901 ( .A1(n807), .A2(n806), .ZN(n1028) );
  NAND2_X1 U902 ( .A1(n808), .A2(n1028), .ZN(n809) );
  XNOR2_X1 U903 ( .A(n809), .B(KEYINPUT91), .ZN(n820) );
  NOR2_X1 U904 ( .A1(n810), .A2(n820), .ZN(n811) );
  XOR2_X1 U905 ( .A(KEYINPUT92), .B(n811), .Z(n812) );
  XNOR2_X1 U906 ( .A(G1986), .B(G290), .ZN(n960) );
  NOR2_X1 U907 ( .A1(G1996), .A2(n908), .ZN(n1021) );
  NOR2_X1 U908 ( .A1(G1991), .A2(n903), .ZN(n816) );
  XNOR2_X1 U909 ( .A(KEYINPUT106), .B(n816), .ZN(n1011) );
  NOR2_X1 U910 ( .A1(G1986), .A2(G290), .ZN(n817) );
  XOR2_X1 U911 ( .A(n817), .B(KEYINPUT105), .Z(n818) );
  NOR2_X1 U912 ( .A1(n1011), .A2(n818), .ZN(n819) );
  NOR2_X1 U913 ( .A1(n820), .A2(n819), .ZN(n821) );
  NOR2_X1 U914 ( .A1(n1021), .A2(n821), .ZN(n822) );
  XNOR2_X1 U915 ( .A(n822), .B(KEYINPUT39), .ZN(n824) );
  NAND2_X1 U916 ( .A1(n824), .A2(n823), .ZN(n826) );
  NAND2_X1 U917 ( .A1(n881), .A2(n825), .ZN(n1012) );
  NAND2_X1 U918 ( .A1(n826), .A2(n1012), .ZN(n828) );
  NAND2_X1 U919 ( .A1(n828), .A2(n827), .ZN(n829) );
  NAND2_X1 U920 ( .A1(n830), .A2(n829), .ZN(n831) );
  XNOR2_X1 U921 ( .A(n831), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U922 ( .A1(G2106), .A2(n832), .ZN(G217) );
  AND2_X1 U923 ( .A1(G15), .A2(G2), .ZN(n833) );
  NAND2_X1 U924 ( .A1(G661), .A2(n833), .ZN(G259) );
  NAND2_X1 U925 ( .A1(G3), .A2(G1), .ZN(n834) );
  NAND2_X1 U926 ( .A1(n835), .A2(n834), .ZN(G188) );
  INV_X1 U928 ( .A(G120), .ZN(G236) );
  INV_X1 U929 ( .A(G96), .ZN(G221) );
  INV_X1 U930 ( .A(G69), .ZN(G235) );
  NOR2_X1 U931 ( .A1(n837), .A2(n836), .ZN(G325) );
  INV_X1 U932 ( .A(G325), .ZN(G261) );
  INV_X1 U933 ( .A(n838), .ZN(G319) );
  XOR2_X1 U934 ( .A(G2100), .B(G2096), .Z(n840) );
  XNOR2_X1 U935 ( .A(KEYINPUT42), .B(G2678), .ZN(n839) );
  XNOR2_X1 U936 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U937 ( .A(KEYINPUT43), .B(G2072), .Z(n842) );
  XNOR2_X1 U938 ( .A(G2067), .B(G2090), .ZN(n841) );
  XNOR2_X1 U939 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U940 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U941 ( .A(G2078), .B(G2084), .ZN(n845) );
  XNOR2_X1 U942 ( .A(n846), .B(n845), .ZN(G227) );
  XNOR2_X1 U943 ( .A(G1961), .B(KEYINPUT108), .ZN(n856) );
  XOR2_X1 U944 ( .A(G1976), .B(G1971), .Z(n848) );
  XNOR2_X1 U945 ( .A(G1986), .B(G1956), .ZN(n847) );
  XNOR2_X1 U946 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U947 ( .A(G1981), .B(G1966), .Z(n850) );
  XNOR2_X1 U948 ( .A(G1996), .B(G1991), .ZN(n849) );
  XNOR2_X1 U949 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U950 ( .A(n852), .B(n851), .Z(n854) );
  XNOR2_X1 U951 ( .A(G2474), .B(KEYINPUT41), .ZN(n853) );
  XNOR2_X1 U952 ( .A(n854), .B(n853), .ZN(n855) );
  XNOR2_X1 U953 ( .A(n856), .B(n855), .ZN(G229) );
  XOR2_X1 U954 ( .A(n857), .B(G286), .Z(n860) );
  XNOR2_X1 U955 ( .A(n858), .B(G171), .ZN(n859) );
  XNOR2_X1 U956 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U957 ( .A(n963), .B(n861), .Z(n862) );
  NOR2_X1 U958 ( .A1(G37), .A2(n862), .ZN(G397) );
  NAND2_X1 U959 ( .A1(n888), .A2(G124), .ZN(n863) );
  XNOR2_X1 U960 ( .A(n863), .B(KEYINPUT44), .ZN(n865) );
  NAND2_X1 U961 ( .A1(G136), .A2(n892), .ZN(n864) );
  NAND2_X1 U962 ( .A1(n865), .A2(n864), .ZN(n866) );
  XNOR2_X1 U963 ( .A(n866), .B(KEYINPUT109), .ZN(n871) );
  NAND2_X1 U964 ( .A1(G100), .A2(n895), .ZN(n868) );
  NAND2_X1 U965 ( .A1(G112), .A2(n887), .ZN(n867) );
  NAND2_X1 U966 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U967 ( .A(KEYINPUT110), .B(n869), .Z(n870) );
  NAND2_X1 U968 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U969 ( .A(n872), .B(KEYINPUT111), .ZN(G162) );
  NAND2_X1 U970 ( .A1(G118), .A2(n887), .ZN(n874) );
  NAND2_X1 U971 ( .A1(G130), .A2(n888), .ZN(n873) );
  NAND2_X1 U972 ( .A1(n874), .A2(n873), .ZN(n880) );
  NAND2_X1 U973 ( .A1(G142), .A2(n892), .ZN(n876) );
  NAND2_X1 U974 ( .A1(G106), .A2(n895), .ZN(n875) );
  NAND2_X1 U975 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U976 ( .A(KEYINPUT45), .B(n877), .Z(n878) );
  XNOR2_X1 U977 ( .A(KEYINPUT112), .B(n878), .ZN(n879) );
  NOR2_X1 U978 ( .A1(n880), .A2(n879), .ZN(n882) );
  XNOR2_X1 U979 ( .A(n882), .B(n881), .ZN(n883) );
  XNOR2_X1 U980 ( .A(n883), .B(n1008), .ZN(n905) );
  XOR2_X1 U981 ( .A(KEYINPUT115), .B(KEYINPUT48), .Z(n885) );
  XNOR2_X1 U982 ( .A(KEYINPUT113), .B(KEYINPUT46), .ZN(n884) );
  XNOR2_X1 U983 ( .A(n885), .B(n884), .ZN(n886) );
  XOR2_X1 U984 ( .A(n886), .B(KEYINPUT117), .Z(n900) );
  NAND2_X1 U985 ( .A1(G115), .A2(n887), .ZN(n890) );
  NAND2_X1 U986 ( .A1(G127), .A2(n888), .ZN(n889) );
  NAND2_X1 U987 ( .A1(n890), .A2(n889), .ZN(n891) );
  XNOR2_X1 U988 ( .A(n891), .B(KEYINPUT47), .ZN(n894) );
  NAND2_X1 U989 ( .A1(G139), .A2(n892), .ZN(n893) );
  NAND2_X1 U990 ( .A1(n894), .A2(n893), .ZN(n898) );
  NAND2_X1 U991 ( .A1(n895), .A2(G103), .ZN(n896) );
  XOR2_X1 U992 ( .A(KEYINPUT114), .B(n896), .Z(n897) );
  NOR2_X1 U993 ( .A1(n898), .A2(n897), .ZN(n1016) );
  XNOR2_X1 U994 ( .A(n1016), .B(KEYINPUT116), .ZN(n899) );
  XNOR2_X1 U995 ( .A(n900), .B(n899), .ZN(n901) );
  XOR2_X1 U996 ( .A(G164), .B(n901), .Z(n902) );
  XNOR2_X1 U997 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U998 ( .A(n905), .B(n904), .Z(n907) );
  XNOR2_X1 U999 ( .A(G160), .B(G162), .ZN(n906) );
  XNOR2_X1 U1000 ( .A(n907), .B(n906), .ZN(n909) );
  XNOR2_X1 U1001 ( .A(n909), .B(n908), .ZN(n910) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n910), .ZN(n911) );
  XNOR2_X1 U1003 ( .A(KEYINPUT118), .B(n911), .ZN(G395) );
  XOR2_X1 U1004 ( .A(G2430), .B(G2451), .Z(n913) );
  XNOR2_X1 U1005 ( .A(G2446), .B(G2427), .ZN(n912) );
  XNOR2_X1 U1006 ( .A(n913), .B(n912), .ZN(n920) );
  XOR2_X1 U1007 ( .A(G2438), .B(KEYINPUT107), .Z(n915) );
  XNOR2_X1 U1008 ( .A(G2443), .B(G2454), .ZN(n914) );
  XNOR2_X1 U1009 ( .A(n915), .B(n914), .ZN(n916) );
  XOR2_X1 U1010 ( .A(n916), .B(G2435), .Z(n918) );
  XNOR2_X1 U1011 ( .A(G1341), .B(G1348), .ZN(n917) );
  XNOR2_X1 U1012 ( .A(n918), .B(n917), .ZN(n919) );
  XNOR2_X1 U1013 ( .A(n920), .B(n919), .ZN(n921) );
  NAND2_X1 U1014 ( .A1(n921), .A2(G14), .ZN(n927) );
  NAND2_X1 U1015 ( .A1(G319), .A2(n927), .ZN(n924) );
  NOR2_X1 U1016 ( .A1(G227), .A2(G229), .ZN(n922) );
  XNOR2_X1 U1017 ( .A(KEYINPUT49), .B(n922), .ZN(n923) );
  NOR2_X1 U1018 ( .A1(n924), .A2(n923), .ZN(n926) );
  NOR2_X1 U1019 ( .A1(G397), .A2(G395), .ZN(n925) );
  NAND2_X1 U1020 ( .A1(n926), .A2(n925), .ZN(G225) );
  INV_X1 U1021 ( .A(G225), .ZN(G308) );
  INV_X1 U1022 ( .A(G108), .ZN(G238) );
  INV_X1 U1023 ( .A(n927), .ZN(G401) );
  XOR2_X1 U1024 ( .A(G2067), .B(G26), .Z(n928) );
  NAND2_X1 U1025 ( .A1(n928), .A2(G28), .ZN(n937) );
  XNOR2_X1 U1026 ( .A(G1996), .B(G32), .ZN(n930) );
  XNOR2_X1 U1027 ( .A(G33), .B(G2072), .ZN(n929) );
  NOR2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(n935) );
  XNOR2_X1 U1029 ( .A(G1991), .B(G25), .ZN(n933) );
  XNOR2_X1 U1030 ( .A(G27), .B(n931), .ZN(n932) );
  NOR2_X1 U1031 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1032 ( .A1(n935), .A2(n934), .ZN(n936) );
  NOR2_X1 U1033 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1034 ( .A(n938), .B(KEYINPUT53), .ZN(n939) );
  XNOR2_X1 U1035 ( .A(n939), .B(KEYINPUT119), .ZN(n942) );
  XOR2_X1 U1036 ( .A(G2084), .B(KEYINPUT54), .Z(n940) );
  XNOR2_X1 U1037 ( .A(G34), .B(n940), .ZN(n941) );
  NAND2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n944) );
  XNOR2_X1 U1039 ( .A(G35), .B(G2090), .ZN(n943) );
  NOR2_X1 U1040 ( .A1(n944), .A2(n943), .ZN(n945) );
  XOR2_X1 U1041 ( .A(KEYINPUT55), .B(n945), .Z(n946) );
  NOR2_X1 U1042 ( .A1(G29), .A2(n946), .ZN(n1005) );
  XNOR2_X1 U1043 ( .A(G1966), .B(G168), .ZN(n948) );
  NAND2_X1 U1044 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1045 ( .A(KEYINPUT57), .B(n949), .ZN(n973) );
  INV_X1 U1046 ( .A(n950), .ZN(n951) );
  NAND2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n957) );
  XNOR2_X1 U1048 ( .A(G1956), .B(KEYINPUT121), .ZN(n953) );
  XNOR2_X1 U1049 ( .A(n953), .B(G299), .ZN(n955) );
  NAND2_X1 U1050 ( .A1(G1971), .A2(G303), .ZN(n954) );
  NAND2_X1 U1051 ( .A1(n955), .A2(n954), .ZN(n956) );
  NOR2_X1 U1052 ( .A1(n957), .A2(n956), .ZN(n962) );
  XNOR2_X1 U1053 ( .A(KEYINPUT122), .B(n958), .ZN(n959) );
  NOR2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1055 ( .A1(n962), .A2(n961), .ZN(n965) );
  XNOR2_X1 U1056 ( .A(G1341), .B(n963), .ZN(n964) );
  NOR2_X1 U1057 ( .A1(n965), .A2(n964), .ZN(n970) );
  XNOR2_X1 U1058 ( .A(n966), .B(G1348), .ZN(n968) );
  XNOR2_X1 U1059 ( .A(G301), .B(G1961), .ZN(n967) );
  NOR2_X1 U1060 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1061 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1062 ( .A(KEYINPUT123), .B(n971), .ZN(n972) );
  NAND2_X1 U1063 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1064 ( .A(n974), .B(KEYINPUT124), .ZN(n977) );
  XNOR2_X1 U1065 ( .A(G16), .B(KEYINPUT56), .ZN(n975) );
  XNOR2_X1 U1066 ( .A(n975), .B(KEYINPUT120), .ZN(n976) );
  NAND2_X1 U1067 ( .A1(n977), .A2(n976), .ZN(n1003) );
  XNOR2_X1 U1068 ( .A(G1986), .B(G24), .ZN(n979) );
  XNOR2_X1 U1069 ( .A(G1971), .B(G22), .ZN(n978) );
  NOR2_X1 U1070 ( .A1(n979), .A2(n978), .ZN(n981) );
  XOR2_X1 U1071 ( .A(G1976), .B(G23), .Z(n980) );
  NAND2_X1 U1072 ( .A1(n981), .A2(n980), .ZN(n983) );
  XOR2_X1 U1073 ( .A(KEYINPUT58), .B(KEYINPUT126), .Z(n982) );
  XNOR2_X1 U1074 ( .A(n983), .B(n982), .ZN(n987) );
  XNOR2_X1 U1075 ( .A(G1966), .B(G21), .ZN(n985) );
  XNOR2_X1 U1076 ( .A(G5), .B(G1961), .ZN(n984) );
  NOR2_X1 U1077 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1078 ( .A1(n987), .A2(n986), .ZN(n998) );
  XNOR2_X1 U1079 ( .A(G20), .B(n988), .ZN(n992) );
  XNOR2_X1 U1080 ( .A(G1341), .B(G19), .ZN(n990) );
  XNOR2_X1 U1081 ( .A(G1981), .B(G6), .ZN(n989) );
  NOR2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n995) );
  XOR2_X1 U1084 ( .A(KEYINPUT59), .B(G1348), .Z(n993) );
  XNOR2_X1 U1085 ( .A(G4), .B(n993), .ZN(n994) );
  NOR2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1087 ( .A(KEYINPUT60), .B(n996), .Z(n997) );
  NOR2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1089 ( .A(n999), .B(KEYINPUT61), .ZN(n1001) );
  XNOR2_X1 U1090 ( .A(G16), .B(KEYINPUT125), .ZN(n1000) );
  NAND2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NOR2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1094 ( .A1(G11), .A2(n1006), .ZN(n1007) );
  XNOR2_X1 U1095 ( .A(n1007), .B(KEYINPUT127), .ZN(n1034) );
  XNOR2_X1 U1096 ( .A(G160), .B(G2084), .ZN(n1009) );
  NAND2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NOR2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1013) );
  NAND2_X1 U1099 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1100 ( .A1(n1015), .A2(n1014), .ZN(n1026) );
  XOR2_X1 U1101 ( .A(G2072), .B(n1016), .Z(n1018) );
  XOR2_X1 U1102 ( .A(G164), .B(G2078), .Z(n1017) );
  NOR2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1104 ( .A(KEYINPUT50), .B(n1019), .Z(n1024) );
  XOR2_X1 U1105 ( .A(G2090), .B(G162), .Z(n1020) );
  NOR2_X1 U1106 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1107 ( .A(KEYINPUT51), .B(n1022), .ZN(n1023) );
  NOR2_X1 U1108 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1109 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1110 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1111 ( .A(KEYINPUT52), .B(n1029), .ZN(n1031) );
  INV_X1 U1112 ( .A(KEYINPUT55), .ZN(n1030) );
  NAND2_X1 U1113 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NAND2_X1 U1114 ( .A1(n1032), .A2(G29), .ZN(n1033) );
  NAND2_X1 U1115 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XOR2_X1 U1116 ( .A(KEYINPUT62), .B(n1035), .Z(G311) );
  INV_X1 U1117 ( .A(G311), .ZN(G150) );
endmodule

