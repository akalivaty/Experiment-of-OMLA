//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 1 0 1 1 0 1 1 1 0 1 0 1 0 1 0 0 0 1 1 1 1 0 0 1 1 1 1 1 1 0 0 1 0 0 0 1 1 0 1 1 0 1 0 0 1 1 0 0 1 0 0 1 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:01 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(G143), .ZN(new_n188));
  AND2_X1   g002(.A1(KEYINPUT65), .A2(G146), .ZN(new_n189));
  NOR2_X1   g003(.A1(KEYINPUT65), .A2(G146), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  AOI21_X1  g005(.A(new_n188), .B1(new_n191), .B2(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(KEYINPUT0), .A2(G128), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n195), .B1(new_n189), .B2(new_n190), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n187), .A2(G143), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n193), .A2(KEYINPUT64), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT64), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n200), .B1(KEYINPUT0), .B2(G128), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n199), .B1(new_n193), .B2(new_n201), .ZN(new_n202));
  AOI22_X1  g016(.A1(new_n192), .A2(new_n194), .B1(new_n198), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G137), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(KEYINPUT11), .A3(G134), .ZN(new_n205));
  INV_X1    g019(.A(G134), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G137), .ZN(new_n207));
  AND2_X1   g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G131), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT66), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n204), .A2(G134), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT11), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AOI211_X1 g027(.A(KEYINPUT66), .B(KEYINPUT11), .C1(new_n204), .C2(G134), .ZN(new_n214));
  OAI211_X1 g028(.A(new_n208), .B(new_n209), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n212), .B1(new_n206), .B2(G137), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(KEYINPUT66), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n211), .A2(new_n210), .A3(new_n212), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n209), .B1(new_n220), .B2(new_n208), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n203), .B1(new_n216), .B2(new_n221), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n209), .B1(new_n211), .B2(new_n207), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n205), .A2(new_n207), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n224), .B1(new_n218), .B2(new_n219), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n223), .B1(new_n225), .B2(new_n209), .ZN(new_n226));
  OR2_X1    g040(.A1(KEYINPUT65), .A2(G146), .ZN(new_n227));
  NAND2_X1  g041(.A1(KEYINPUT65), .A2(G146), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n227), .A2(G143), .A3(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n188), .ZN(new_n230));
  INV_X1    g044(.A(G128), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n231), .A2(KEYINPUT1), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n229), .A2(new_n230), .A3(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n231), .B1(new_n229), .B2(KEYINPUT1), .ZN(new_n234));
  INV_X1    g048(.A(new_n197), .ZN(new_n235));
  XNOR2_X1  g049(.A(KEYINPUT65), .B(G146), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n235), .B1(new_n236), .B2(new_n195), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n233), .B1(new_n234), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n226), .A2(new_n238), .ZN(new_n239));
  XOR2_X1   g053(.A(KEYINPUT2), .B(G113), .Z(new_n240));
  XNOR2_X1  g054(.A(G116), .B(G119), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g056(.A(KEYINPUT2), .B(G113), .ZN(new_n243));
  INV_X1    g057(.A(G116), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n244), .A2(G119), .ZN(new_n245));
  INV_X1    g059(.A(G119), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n246), .A2(G116), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n243), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT67), .ZN(new_n249));
  AND3_X1   g063(.A1(new_n242), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n249), .B1(new_n242), .B2(new_n248), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  AND3_X1   g066(.A1(new_n222), .A2(new_n239), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n242), .A2(new_n248), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n255), .B1(new_n222), .B2(new_n239), .ZN(new_n256));
  OAI21_X1  g070(.A(KEYINPUT28), .B1(new_n253), .B2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n222), .A2(new_n252), .A3(new_n239), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT28), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NOR2_X1   g074(.A1(G237), .A2(G953), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G210), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n262), .B(KEYINPUT27), .ZN(new_n263));
  XNOR2_X1  g077(.A(KEYINPUT26), .B(G101), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n263), .B(new_n264), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n257), .A2(KEYINPUT69), .A3(new_n260), .A4(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n265), .ZN(new_n267));
  NOR3_X1   g081(.A1(new_n189), .A2(new_n190), .A3(new_n195), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT1), .ZN(new_n269));
  OAI21_X1  g083(.A(G128), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  AOI22_X1  g084(.A1(new_n270), .A2(new_n198), .B1(new_n192), .B2(new_n232), .ZN(new_n271));
  INV_X1    g085(.A(new_n223), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n215), .A2(new_n272), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n229), .A2(new_n230), .A3(new_n194), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n200), .A2(KEYINPUT0), .A3(G128), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT0), .ZN(new_n277));
  AOI21_X1  g091(.A(KEYINPUT64), .B1(new_n277), .B2(new_n231), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n276), .B1(new_n278), .B2(new_n194), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n275), .B1(new_n237), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n208), .B1(new_n213), .B2(new_n214), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G131), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n280), .B1(new_n282), .B2(new_n215), .ZN(new_n283));
  OAI21_X1  g097(.A(KEYINPUT30), .B1(new_n274), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT30), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n222), .A2(new_n285), .A3(new_n239), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n255), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n267), .B1(new_n287), .B2(new_n253), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT29), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n266), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n282), .A2(new_n215), .ZN(new_n291));
  AOI22_X1  g105(.A1(new_n291), .A2(new_n203), .B1(new_n238), .B2(new_n226), .ZN(new_n292));
  AOI21_X1  g106(.A(KEYINPUT28), .B1(new_n292), .B2(new_n252), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n258), .B1(new_n292), .B2(new_n255), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n293), .B1(new_n294), .B2(KEYINPUT28), .ZN(new_n295));
  AOI21_X1  g109(.A(KEYINPUT69), .B1(new_n295), .B2(new_n265), .ZN(new_n296));
  OAI21_X1  g110(.A(KEYINPUT70), .B1(new_n290), .B2(new_n296), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n222), .A2(new_n285), .A3(new_n239), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n285), .B1(new_n222), .B2(new_n239), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n254), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(new_n258), .ZN(new_n301));
  AOI21_X1  g115(.A(KEYINPUT29), .B1(new_n301), .B2(new_n267), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n257), .A2(new_n260), .A3(new_n265), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT69), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT70), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n302), .A2(new_n305), .A3(new_n306), .A4(new_n266), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT71), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n258), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n292), .A2(KEYINPUT71), .A3(new_n252), .ZN(new_n310));
  OAI22_X1  g124(.A1(new_n274), .A2(new_n283), .B1(new_n251), .B2(new_n250), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT72), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n293), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n260), .A2(KEYINPUT72), .ZN(new_n315));
  AOI22_X1  g129(.A1(KEYINPUT28), .A2(new_n312), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n267), .A2(new_n289), .ZN(new_n317));
  AOI21_X1  g131(.A(G902), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n297), .A2(new_n307), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G472), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n284), .A2(new_n286), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n253), .B1(new_n321), .B2(new_n254), .ZN(new_n322));
  AOI21_X1  g136(.A(KEYINPUT31), .B1(new_n322), .B2(new_n265), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT31), .ZN(new_n324));
  NOR4_X1   g138(.A1(new_n287), .A2(new_n324), .A3(new_n253), .A4(new_n267), .ZN(new_n325));
  OAI22_X1  g139(.A1(new_n323), .A2(new_n325), .B1(new_n295), .B2(new_n265), .ZN(new_n326));
  INV_X1    g140(.A(G472), .ZN(new_n327));
  INV_X1    g141(.A(G902), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n326), .A2(KEYINPUT32), .A3(new_n327), .A4(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n330));
  XNOR2_X1  g144(.A(KEYINPUT68), .B(KEYINPUT32), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n320), .A2(new_n329), .A3(new_n332), .ZN(new_n333));
  XOR2_X1   g147(.A(KEYINPUT22), .B(G137), .Z(new_n334));
  XNOR2_X1  g148(.A(new_n334), .B(KEYINPUT76), .ZN(new_n335));
  INV_X1    g149(.A(G953), .ZN(new_n336));
  AND3_X1   g150(.A1(new_n336), .A2(G221), .A3(G234), .ZN(new_n337));
  XOR2_X1   g151(.A(new_n335), .B(new_n337), .Z(new_n338));
  NAND2_X1  g152(.A1(new_n231), .A2(G119), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT23), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n246), .A2(G128), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n231), .A2(KEYINPUT23), .A3(G119), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(G110), .ZN(new_n345));
  XNOR2_X1  g159(.A(KEYINPUT24), .B(G110), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT73), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n346), .B(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n339), .A2(new_n342), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n345), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(G125), .ZN(new_n351));
  NOR3_X1   g165(.A1(new_n351), .A2(KEYINPUT16), .A3(G140), .ZN(new_n352));
  XNOR2_X1  g166(.A(G125), .B(G140), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n352), .B1(new_n353), .B2(KEYINPUT16), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n354), .B(new_n187), .ZN(new_n355));
  OAI21_X1  g169(.A(KEYINPUT74), .B1(new_n350), .B2(new_n355), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n354), .B(G146), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT74), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n346), .B(KEYINPUT73), .ZN(new_n359));
  INV_X1    g173(.A(new_n349), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n357), .A2(new_n358), .A3(new_n361), .A4(new_n345), .ZN(new_n362));
  AND2_X1   g176(.A1(new_n356), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT75), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n344), .A2(G110), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n365), .B1(new_n348), .B2(new_n349), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n354), .A2(G146), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n191), .A2(new_n353), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n364), .B1(new_n366), .B2(new_n369), .ZN(new_n370));
  OAI22_X1  g184(.A1(new_n359), .A2(new_n360), .B1(G110), .B2(new_n344), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n371), .A2(KEYINPUT75), .A3(new_n367), .A4(new_n368), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n338), .B1(new_n363), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT25), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n370), .A2(new_n372), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n356), .A2(new_n362), .ZN(new_n377));
  INV_X1    g191(.A(new_n338), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n374), .A2(new_n375), .A3(new_n379), .A4(new_n328), .ZN(new_n380));
  INV_X1    g194(.A(G217), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n381), .B1(G234), .B2(new_n328), .ZN(new_n382));
  AND2_X1   g196(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n374), .A2(new_n328), .A3(new_n379), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT25), .ZN(new_n385));
  AND2_X1   g199(.A1(new_n374), .A2(new_n379), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n382), .A2(G902), .ZN(new_n387));
  AOI22_X1  g201(.A1(new_n383), .A2(new_n385), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT3), .ZN(new_n389));
  INV_X1    g203(.A(G107), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n389), .B1(new_n390), .B2(G104), .ZN(new_n391));
  INV_X1    g205(.A(G104), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n391), .B1(new_n392), .B2(G107), .ZN(new_n393));
  OR2_X1    g207(.A1(KEYINPUT78), .A2(G107), .ZN(new_n394));
  NAND2_X1  g208(.A1(KEYINPUT78), .A2(G107), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n394), .A2(new_n389), .A3(G104), .A4(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(G101), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n393), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(G104), .B1(new_n394), .B2(new_n395), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n392), .A2(G107), .ZN(new_n400));
  OAI21_X1  g214(.A(G101), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n231), .B1(new_n197), .B2(KEYINPUT1), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n402), .B1(new_n229), .B2(new_n230), .ZN(new_n403));
  AND3_X1   g217(.A1(new_n229), .A2(new_n230), .A3(new_n232), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n398), .B(new_n401), .C1(new_n403), .C2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT10), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AND2_X1   g221(.A1(new_n401), .A2(new_n398), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n408), .A2(KEYINPUT10), .A3(new_n238), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n389), .A2(G104), .ZN(new_n410));
  AND2_X1   g224(.A1(KEYINPUT78), .A2(G107), .ZN(new_n411));
  NOR2_X1   g225(.A1(KEYINPUT78), .A2(G107), .ZN(new_n412));
  NOR3_X1   g226(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(KEYINPUT3), .B1(new_n392), .B2(G107), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n414), .A2(new_n400), .ZN(new_n415));
  OAI21_X1  g229(.A(G101), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n416), .A2(KEYINPUT4), .A3(new_n398), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT4), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n418), .B(G101), .C1(new_n413), .C2(new_n415), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n417), .A2(new_n203), .A3(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n291), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n407), .A2(new_n409), .A3(new_n420), .A4(new_n421), .ZN(new_n422));
  XOR2_X1   g236(.A(G110), .B(G140), .Z(new_n423));
  XNOR2_X1  g237(.A(new_n423), .B(KEYINPUT77), .ZN(new_n424));
  INV_X1    g238(.A(G227), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n425), .A2(G953), .ZN(new_n426));
  XOR2_X1   g240(.A(new_n424), .B(new_n426), .Z(new_n427));
  NAND2_X1  g241(.A1(new_n422), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n407), .A2(new_n409), .A3(new_n420), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n291), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n422), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n401), .A2(new_n398), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n270), .A2(new_n198), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT79), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n434), .A2(new_n435), .A3(new_n436), .A4(new_n233), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n405), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n436), .B1(new_n271), .B2(new_n434), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n291), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT12), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  OAI211_X1 g256(.A(KEYINPUT12), .B(new_n291), .C1(new_n438), .C2(new_n439), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n433), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n432), .B(G469), .C1(new_n444), .C2(new_n427), .ZN(new_n445));
  INV_X1    g259(.A(G469), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n428), .B1(new_n442), .B2(new_n443), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n427), .B1(new_n431), .B2(new_n422), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n446), .B(new_n328), .C1(new_n447), .C2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(G469), .A2(G902), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n445), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n261), .A2(G143), .A3(G214), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(G143), .B1(new_n261), .B2(G214), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(KEYINPUT18), .A2(G131), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n351), .A2(G140), .ZN(new_n457));
  INV_X1    g271(.A(G140), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n458), .A2(G125), .ZN(new_n459));
  OAI21_X1  g273(.A(G146), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  AOI22_X1  g274(.A1(new_n455), .A2(new_n456), .B1(new_n368), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT87), .ZN(new_n462));
  OAI211_X1 g276(.A(KEYINPUT18), .B(G131), .C1(new_n453), .C2(new_n454), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n454), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n465), .A2(new_n452), .A3(new_n456), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n368), .A2(new_n460), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n463), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(KEYINPUT87), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n464), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n465), .A2(new_n452), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n471), .A2(KEYINPUT17), .A3(G131), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n455), .A2(new_n209), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n471), .A2(G131), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n355), .B(new_n472), .C1(new_n475), .C2(KEYINPUT17), .ZN(new_n476));
  XNOR2_X1  g290(.A(G113), .B(G122), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n477), .B(KEYINPUT89), .ZN(new_n478));
  XOR2_X1   g292(.A(KEYINPUT88), .B(G104), .Z(new_n479));
  XNOR2_X1  g293(.A(new_n478), .B(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n470), .A2(new_n476), .A3(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n480), .B1(new_n470), .B2(new_n476), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n328), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n484), .A2(G475), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n353), .B(KEYINPUT19), .ZN(new_n486));
  AOI22_X1  g300(.A1(new_n486), .A2(new_n191), .B1(G146), .B2(new_n354), .ZN(new_n487));
  AOI22_X1  g301(.A1(new_n464), .A2(new_n469), .B1(new_n487), .B2(new_n475), .ZN(new_n488));
  OAI21_X1  g302(.A(KEYINPUT90), .B1(new_n488), .B2(new_n480), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n487), .A2(new_n475), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n462), .B1(new_n461), .B2(new_n463), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n468), .A2(KEYINPUT87), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT90), .ZN(new_n494));
  INV_X1    g308(.A(new_n480), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n489), .A2(new_n496), .A3(new_n481), .ZN(new_n497));
  NOR2_X1   g311(.A1(G475), .A2(G902), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  XOR2_X1   g313(.A(KEYINPUT86), .B(KEYINPUT20), .Z(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT20), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n497), .A2(new_n503), .A3(new_n498), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n485), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n244), .A2(G122), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n244), .A2(G122), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n394), .A2(new_n395), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n231), .A2(G143), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n195), .A2(G128), .ZN(new_n513));
  OR3_X1    g327(.A1(new_n512), .A2(new_n513), .A3(G134), .ZN(new_n514));
  OAI21_X1  g328(.A(G134), .B1(new_n512), .B2(new_n513), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n511), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n508), .B1(new_n506), .B2(KEYINPUT14), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(KEYINPUT91), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT91), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n519), .B(new_n508), .C1(new_n506), .C2(KEYINPUT14), .ZN(new_n520));
  OR2_X1    g334(.A1(new_n508), .A2(KEYINPUT14), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n518), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT92), .ZN(new_n523));
  AND3_X1   g337(.A1(new_n522), .A2(new_n523), .A3(G107), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n523), .B1(new_n522), .B2(G107), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n516), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(KEYINPUT13), .B1(new_n195), .B2(G128), .ZN(new_n527));
  MUX2_X1   g341(.A(new_n527), .B(KEYINPUT13), .S(new_n512), .Z(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(G134), .ZN(new_n529));
  AND2_X1   g343(.A1(new_n509), .A2(new_n510), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n529), .B(new_n514), .C1(new_n530), .C2(new_n511), .ZN(new_n531));
  XNOR2_X1  g345(.A(KEYINPUT9), .B(G234), .ZN(new_n532));
  NOR3_X1   g346(.A1(new_n532), .A2(new_n381), .A3(G953), .ZN(new_n533));
  AND3_X1   g347(.A1(new_n526), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n533), .B1(new_n526), .B2(new_n531), .ZN(new_n535));
  OAI211_X1 g349(.A(KEYINPUT93), .B(new_n328), .C1(new_n534), .C2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(G478), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n537), .A2(KEYINPUT15), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n526), .A2(new_n531), .ZN(new_n540));
  INV_X1    g354(.A(new_n533), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n526), .A2(new_n531), .A3(new_n533), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n538), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n544), .A2(KEYINPUT93), .A3(new_n328), .A4(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(G234), .A2(G237), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n547), .A2(G952), .A3(new_n336), .ZN(new_n548));
  XNOR2_X1  g362(.A(KEYINPUT21), .B(G898), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n547), .A2(G902), .A3(G953), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n548), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AND3_X1   g366(.A1(new_n539), .A2(new_n546), .A3(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(G221), .B1(new_n532), .B2(G902), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n451), .A2(new_n505), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(G214), .B1(G237), .B2(G902), .ZN(new_n556));
  AOI21_X1  g370(.A(G125), .B1(new_n435), .B2(new_n233), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n275), .B(G125), .C1(new_n237), .C2(new_n279), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(KEYINPUT84), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n336), .A2(G224), .ZN(new_n561));
  XOR2_X1   g375(.A(new_n561), .B(KEYINPUT83), .Z(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n238), .A2(new_n351), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT84), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n564), .A2(new_n565), .A3(new_n558), .ZN(new_n566));
  AND3_X1   g380(.A1(new_n560), .A2(new_n563), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n563), .B1(new_n560), .B2(new_n566), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n417), .A2(new_n254), .A3(new_n419), .ZN(new_n570));
  INV_X1    g384(.A(G113), .ZN(new_n571));
  XOR2_X1   g385(.A(KEYINPUT80), .B(KEYINPUT5), .Z(new_n572));
  AOI21_X1  g386(.A(new_n571), .B1(new_n572), .B2(new_n245), .ZN(new_n573));
  XNOR2_X1  g387(.A(KEYINPUT80), .B(KEYINPUT5), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n241), .A2(new_n574), .ZN(new_n575));
  AOI22_X1  g389(.A1(new_n573), .A2(new_n575), .B1(new_n241), .B2(new_n240), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n408), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n570), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(G110), .B(G122), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  XOR2_X1   g394(.A(KEYINPUT82), .B(KEYINPUT6), .Z(new_n581));
  NAND3_X1  g395(.A1(new_n578), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n578), .A2(new_n580), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n570), .A2(new_n577), .A3(new_n579), .ZN(new_n584));
  AND4_X1   g398(.A1(KEYINPUT81), .A2(new_n583), .A3(KEYINPUT6), .A4(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT6), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n586), .B1(new_n578), .B2(new_n580), .ZN(new_n587));
  AOI21_X1  g401(.A(KEYINPUT81), .B1(new_n587), .B2(new_n584), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n569), .B(new_n582), .C1(new_n585), .C2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n584), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n562), .A2(KEYINPUT7), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n591), .B1(new_n557), .B2(new_n559), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n564), .A2(KEYINPUT7), .A3(new_n562), .A4(new_n558), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n241), .A2(KEYINPUT5), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n573), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n242), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n408), .ZN(new_n597));
  XOR2_X1   g411(.A(new_n579), .B(KEYINPUT8), .Z(new_n598));
  AOI21_X1  g412(.A(new_n598), .B1(new_n576), .B2(new_n434), .ZN(new_n599));
  AOI22_X1  g413(.A1(new_n592), .A2(new_n593), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n590), .B1(new_n600), .B2(KEYINPUT85), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n592), .A2(new_n593), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n599), .A2(new_n597), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT85), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(G902), .B1(new_n601), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(G210), .B1(G237), .B2(G902), .ZN(new_n608));
  AND3_X1   g422(.A1(new_n589), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n608), .B1(new_n589), .B2(new_n607), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n556), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n555), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n333), .A2(new_n388), .A3(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(G101), .ZN(G3));
  OAI211_X1 g428(.A(new_n556), .B(new_n552), .C1(new_n609), .C2(new_n610), .ZN(new_n615));
  INV_X1    g429(.A(new_n485), .ZN(new_n616));
  INV_X1    g430(.A(new_n504), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n500), .B1(new_n497), .B2(new_n498), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  AOI211_X1 g433(.A(G478), .B(G902), .C1(new_n542), .C2(new_n543), .ZN(new_n620));
  OAI21_X1  g434(.A(KEYINPUT33), .B1(new_n533), .B2(KEYINPUT94), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n621), .B1(new_n534), .B2(new_n535), .ZN(new_n622));
  INV_X1    g436(.A(new_n621), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n542), .A2(new_n543), .A3(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n622), .A2(new_n624), .A3(new_n328), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n620), .B1(new_n625), .B2(G478), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n619), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n615), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n451), .A2(new_n554), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n295), .A2(new_n265), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n300), .A2(new_n258), .A3(new_n265), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(new_n324), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n322), .A2(KEYINPUT31), .A3(new_n265), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n631), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g449(.A(G472), .B1(new_n635), .B2(G902), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n388), .A2(new_n636), .A3(new_n330), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n628), .A2(new_n630), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT34), .B(G104), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G6));
  INV_X1    g454(.A(new_n556), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n589), .A2(new_n607), .ZN(new_n642));
  INV_X1    g456(.A(new_n608), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n589), .A2(new_n607), .A3(new_n608), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n641), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n485), .B1(new_n546), .B2(new_n539), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n497), .A2(new_n498), .A3(new_n500), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n502), .A2(new_n648), .ZN(new_n649));
  AND2_X1   g463(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n646), .A2(new_n650), .A3(new_n552), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n636), .A2(new_n330), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n386), .A2(new_n387), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n384), .A2(KEYINPUT25), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n380), .A2(new_n382), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NOR3_X1   g471(.A1(new_n653), .A2(new_n657), .A3(new_n629), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n652), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT35), .B(G107), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G9));
  NAND2_X1  g475(.A1(new_n376), .A2(new_n377), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n338), .A2(KEYINPUT36), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n387), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n665), .B1(new_n655), .B2(new_n656), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n653), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n612), .ZN(new_n669));
  XNOR2_X1  g483(.A(KEYINPUT37), .B(G110), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(KEYINPUT95), .ZN(new_n671));
  XOR2_X1   g485(.A(new_n671), .B(KEYINPUT96), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n669), .B(new_n672), .ZN(G12));
  OR2_X1    g487(.A1(new_n551), .A2(G900), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n548), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n647), .A2(new_n649), .A3(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n676), .A2(new_n629), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n333), .A2(new_n646), .A3(new_n666), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G128), .ZN(G30));
  NAND2_X1  g493(.A1(new_n644), .A2(new_n645), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT98), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n644), .A2(KEYINPUT98), .A3(new_n645), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g498(.A(KEYINPUT97), .B(KEYINPUT38), .Z(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n675), .B(KEYINPUT39), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n630), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(KEYINPUT40), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT40), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n630), .A2(new_n690), .A3(new_n687), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n312), .A2(new_n267), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n632), .A2(new_n692), .A3(G472), .ZN(new_n693));
  NAND2_X1  g507(.A1(G472), .A2(G902), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT99), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n696), .A2(new_n332), .A3(new_n329), .ZN(new_n697));
  AND2_X1   g511(.A1(new_n539), .A2(new_n546), .ZN(new_n698));
  NOR4_X1   g512(.A1(new_n666), .A2(new_n505), .A3(new_n698), .A4(new_n641), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n689), .A2(new_n691), .A3(new_n697), .A4(new_n699), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n686), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(new_n195), .ZN(G45));
  NAND3_X1  g516(.A1(new_n619), .A2(new_n626), .A3(new_n675), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n703), .A2(new_n629), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n333), .A2(new_n646), .A3(new_n666), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G146), .ZN(G48));
  OAI21_X1  g520(.A(new_n328), .B1(new_n447), .B2(new_n448), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(G469), .ZN(new_n708));
  AND3_X1   g522(.A1(new_n708), .A2(new_n554), .A3(new_n449), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n333), .A2(new_n628), .A3(new_n388), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(KEYINPUT41), .B(G113), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G15));
  AND2_X1   g526(.A1(new_n333), .A2(new_n388), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT100), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n713), .A2(new_n714), .A3(new_n652), .A4(new_n709), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n333), .A2(new_n388), .A3(new_n709), .ZN(new_n716));
  OAI21_X1  g530(.A(KEYINPUT100), .B1(new_n716), .B2(new_n651), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G116), .ZN(G18));
  NAND3_X1  g533(.A1(new_n708), .A2(new_n554), .A3(new_n449), .ZN(new_n720));
  OAI21_X1  g534(.A(KEYINPUT101), .B1(new_n611), .B2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT101), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n646), .A2(new_n722), .A3(new_n709), .ZN(new_n723));
  AND2_X1   g537(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n505), .A2(new_n553), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n333), .A2(new_n725), .A3(new_n666), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(KEYINPUT102), .B(G119), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(G21));
  AOI21_X1  g543(.A(new_n327), .B1(new_n326), .B2(new_n328), .ZN(new_n730));
  NOR2_X1   g544(.A1(G472), .A2(G902), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n312), .A2(KEYINPUT28), .ZN(new_n733));
  AND2_X1   g547(.A1(new_n314), .A2(new_n315), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n267), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n633), .A2(new_n634), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n732), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n730), .A2(new_n657), .A3(new_n737), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n505), .A2(new_n698), .ZN(new_n739));
  INV_X1    g553(.A(new_n552), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n720), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n738), .A2(new_n646), .A3(new_n739), .A4(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G122), .ZN(G24));
  NAND2_X1  g557(.A1(new_n721), .A2(new_n723), .ZN(new_n744));
  INV_X1    g558(.A(new_n737), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n745), .A2(new_n636), .A3(new_n666), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n746), .A2(new_n703), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G125), .ZN(G27));
  NAND4_X1  g563(.A1(new_n644), .A2(new_n556), .A3(new_n645), .A4(new_n554), .ZN(new_n750));
  XOR2_X1   g564(.A(new_n450), .B(KEYINPUT103), .Z(new_n751));
  AND3_X1   g565(.A1(new_n445), .A2(new_n449), .A3(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(new_n703), .ZN(new_n754));
  AND3_X1   g568(.A1(new_n753), .A2(KEYINPUT42), .A3(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n330), .B(KEYINPUT32), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n657), .B1(new_n756), .B2(new_n320), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n333), .A2(new_n388), .A3(new_n753), .A4(new_n754), .ZN(new_n759));
  XOR2_X1   g573(.A(KEYINPUT104), .B(KEYINPUT42), .Z(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n758), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G131), .ZN(G33));
  INV_X1    g577(.A(new_n676), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n333), .A2(new_n764), .A3(new_n753), .A4(new_n388), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G134), .ZN(G36));
  NAND3_X1  g580(.A1(new_n644), .A2(new_n556), .A3(new_n645), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n505), .A2(new_n626), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT43), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(new_n653), .A3(new_n666), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT44), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n768), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(KEYINPUT107), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT107), .ZN(new_n776));
  OAI211_X1 g590(.A(new_n776), .B(new_n768), .C1(new_n772), .C2(new_n773), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n772), .A2(new_n773), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n775), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n432), .B1(new_n444), .B2(new_n427), .ZN(new_n781));
  OR2_X1    g595(.A1(new_n781), .A2(KEYINPUT45), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(KEYINPUT45), .ZN(new_n783));
  AOI211_X1 g597(.A(KEYINPUT105), .B(new_n446), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT105), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n781), .B(KEYINPUT45), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n785), .B1(new_n786), .B2(G469), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n751), .B1(new_n784), .B2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT46), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n449), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n786), .A2(G469), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(KEYINPUT105), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n786), .A2(new_n785), .A3(G469), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g608(.A(KEYINPUT46), .B1(new_n794), .B2(new_n751), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n554), .B(new_n687), .C1(new_n790), .C2(new_n795), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n796), .A2(KEYINPUT106), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n796), .A2(KEYINPUT106), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n780), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G137), .ZN(G39));
  NOR4_X1   g614(.A1(new_n333), .A2(new_n388), .A3(new_n703), .A4(new_n767), .ZN(new_n801));
  OAI211_X1 g615(.A(KEYINPUT47), .B(new_n554), .C1(new_n790), .C2(new_n795), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n794), .A2(KEYINPUT46), .A3(new_n751), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n788), .A2(new_n789), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n804), .A2(new_n805), .A3(new_n449), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT47), .B1(new_n806), .B2(new_n554), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n801), .B1(new_n803), .B2(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(KEYINPUT108), .B(G140), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n808), .B(new_n809), .ZN(G42));
  INV_X1    g624(.A(new_n697), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n708), .A2(new_n449), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n813), .A2(new_n750), .ZN(new_n814));
  INV_X1    g628(.A(new_n548), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n811), .A2(new_n388), .A3(new_n814), .A4(new_n815), .ZN(new_n816));
  XOR2_X1   g630(.A(new_n816), .B(KEYINPUT114), .Z(new_n817));
  INV_X1    g631(.A(new_n627), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n771), .A2(new_n815), .A3(new_n814), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(new_n757), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(KEYINPUT48), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n336), .A2(G952), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n771), .A2(new_n815), .A3(new_n738), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n823), .B1(new_n824), .B2(new_n744), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n819), .A2(new_n822), .A3(new_n825), .ZN(new_n826));
  XOR2_X1   g640(.A(new_n826), .B(KEYINPUT115), .Z(new_n827));
  NAND3_X1  g641(.A1(new_n824), .A2(new_n641), .A3(new_n709), .ZN(new_n828));
  INV_X1    g642(.A(new_n685), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n684), .B(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT50), .ZN(new_n831));
  OAI22_X1  g645(.A1(new_n828), .A2(new_n830), .B1(KEYINPUT113), .B2(new_n831), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n831), .A2(KEYINPUT113), .ZN(new_n833));
  OR2_X1    g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n619), .A2(new_n626), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n817), .A2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n746), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n820), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n832), .A2(new_n833), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n834), .A2(new_n836), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n554), .B1(new_n790), .B2(new_n795), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT47), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n843), .B(new_n802), .C1(new_n554), .C2(new_n813), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n824), .A2(new_n768), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n840), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n827), .B1(new_n846), .B2(KEYINPUT51), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n847), .B1(KEYINPUT51), .B2(new_n846), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n710), .B1(new_n724), .B2(new_n726), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n613), .A2(new_n638), .A3(new_n669), .A4(new_n742), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT109), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n502), .A2(new_n504), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n647), .A2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n851), .B1(new_n854), .B2(new_n615), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n646), .A2(new_n853), .A3(KEYINPUT109), .A4(new_n552), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n855), .A2(new_n658), .A3(new_n856), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n849), .A2(new_n850), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n747), .A2(new_n753), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n765), .A2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT110), .ZN(new_n861));
  INV_X1    g675(.A(new_n649), .ZN(new_n862));
  INV_X1    g676(.A(new_n675), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n863), .B1(new_n484), .B2(G475), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n864), .A2(new_n539), .A3(new_n546), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n861), .B1(new_n862), .B2(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n698), .A2(new_n649), .A3(KEYINPUT110), .A4(new_n864), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n767), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n667), .A2(new_n629), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n868), .A2(new_n333), .A3(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT111), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n868), .A2(new_n333), .A3(KEYINPUT111), .A4(new_n869), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n860), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n858), .A2(new_n718), .A3(new_n762), .A4(new_n874), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n611), .A2(new_n505), .A3(new_n698), .ZN(new_n876));
  INV_X1    g690(.A(new_n554), .ZN(new_n877));
  NOR4_X1   g691(.A1(new_n752), .A2(new_n666), .A3(new_n877), .A4(new_n863), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n876), .A2(new_n878), .A3(new_n697), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n748), .A2(new_n678), .A3(new_n879), .A4(new_n705), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(KEYINPUT52), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n875), .A2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT53), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g698(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n884), .B1(new_n882), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(KEYINPUT54), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n885), .B1(new_n875), .B2(new_n881), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n849), .A2(new_n850), .ZN(new_n889));
  INV_X1    g703(.A(new_n857), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n889), .A2(new_n718), .A3(new_n890), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n678), .A2(new_n705), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n892), .A2(KEYINPUT52), .A3(new_n748), .A4(new_n879), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT52), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n880), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n872), .A2(new_n873), .ZN(new_n897));
  AND4_X1   g711(.A1(new_n762), .A2(new_n897), .A3(new_n765), .A4(new_n859), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n891), .A2(KEYINPUT53), .A3(new_n896), .A4(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n888), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n887), .B1(KEYINPUT54), .B2(new_n900), .ZN(new_n901));
  OAI22_X1  g715(.A1(new_n848), .A2(new_n901), .B1(G952), .B2(G953), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n812), .B(KEYINPUT49), .ZN(new_n903));
  NOR4_X1   g717(.A1(new_n769), .A2(new_n657), .A3(new_n641), .A4(new_n877), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n686), .A2(new_n811), .A3(new_n903), .A4(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n902), .A2(new_n905), .ZN(G75));
  NAND3_X1  g720(.A1(new_n900), .A2(G210), .A3(G902), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(KEYINPUT117), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT117), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n582), .B1(new_n585), .B2(new_n588), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(new_n569), .Z(new_n913));
  XNOR2_X1  g727(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n913), .B(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n916), .A2(KEYINPUT56), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n909), .A2(new_n911), .A3(new_n917), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n916), .B1(new_n908), .B2(KEYINPUT56), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n336), .A2(G952), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n918), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(KEYINPUT118), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT118), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n918), .A2(new_n924), .A3(new_n919), .A4(new_n921), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n923), .A2(new_n925), .ZN(G51));
  XOR2_X1   g740(.A(new_n900), .B(KEYINPUT54), .Z(new_n927));
  XNOR2_X1  g741(.A(new_n751), .B(KEYINPUT119), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT57), .Z(new_n929));
  OAI22_X1  g743(.A1(new_n927), .A2(new_n929), .B1(new_n448), .B2(new_n447), .ZN(new_n930));
  INV_X1    g744(.A(new_n900), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n931), .A2(new_n328), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n932), .A2(new_n793), .A3(new_n792), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n920), .B1(new_n930), .B2(new_n933), .ZN(G54));
  NAND4_X1  g748(.A1(new_n932), .A2(KEYINPUT58), .A3(G475), .A4(new_n497), .ZN(new_n935));
  INV_X1    g749(.A(new_n497), .ZN(new_n936));
  INV_X1    g750(.A(new_n932), .ZN(new_n937));
  NAND2_X1  g751(.A1(KEYINPUT58), .A2(G475), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n935), .A2(new_n921), .A3(new_n939), .ZN(G60));
  AND2_X1   g754(.A1(new_n622), .A2(new_n624), .ZN(new_n941));
  NAND2_X1  g755(.A1(G478), .A2(G902), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT59), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n941), .B1(new_n901), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n941), .A2(new_n943), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n921), .B1(new_n927), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n944), .A2(new_n946), .ZN(G63));
  NAND2_X1  g761(.A1(G217), .A2(G902), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(KEYINPUT60), .Z(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n950), .B1(new_n888), .B2(new_n899), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n921), .B1(new_n951), .B2(new_n386), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n951), .A2(new_n664), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n953), .A2(KEYINPUT61), .A3(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT121), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n952), .A2(new_n956), .ZN(new_n957));
  OAI211_X1 g771(.A(KEYINPUT121), .B(new_n921), .C1(new_n951), .C2(new_n386), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT120), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n954), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n951), .A2(KEYINPUT120), .A3(new_n664), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n957), .A2(new_n958), .A3(new_n960), .A4(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT61), .ZN(new_n963));
  AND3_X1   g777(.A1(new_n962), .A2(KEYINPUT122), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(KEYINPUT122), .B1(new_n962), .B2(new_n963), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n955), .B1(new_n964), .B2(new_n965), .ZN(G66));
  NAND2_X1  g780(.A1(new_n891), .A2(new_n336), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n550), .A2(G224), .A3(G953), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n912), .B1(G898), .B2(new_n336), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n969), .B(new_n970), .Z(G69));
  INV_X1    g785(.A(KEYINPUT62), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n892), .A2(new_n748), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n972), .B1(new_n973), .B2(new_n701), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n689), .A2(new_n697), .A3(new_n699), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n975), .A2(new_n830), .A3(new_n691), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n976), .A2(KEYINPUT62), .A3(new_n748), .A4(new_n892), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  AOI211_X1 g792(.A(new_n767), .B(new_n688), .C1(new_n627), .C2(new_n854), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n979), .A2(new_n713), .ZN(new_n980));
  INV_X1    g794(.A(new_n980), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n808), .A2(new_n978), .A3(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(new_n798), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n796), .A2(KEYINPUT106), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n779), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n336), .B1(new_n982), .B2(new_n985), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n321), .B(new_n486), .Z(new_n987));
  XOR2_X1   g801(.A(new_n987), .B(KEYINPUT123), .Z(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n986), .A2(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT124), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n986), .A2(KEYINPUT124), .A3(new_n989), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n762), .A2(new_n748), .A3(new_n765), .A4(new_n892), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n843), .A2(new_n802), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n994), .B1(new_n995), .B2(new_n801), .ZN(new_n996));
  AND2_X1   g810(.A1(new_n757), .A2(new_n876), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n997), .B1(new_n797), .B2(new_n798), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n996), .A2(new_n799), .A3(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT125), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n996), .A2(new_n799), .A3(new_n998), .A4(KEYINPUT125), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n1001), .A2(new_n336), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n987), .B1(G900), .B2(G953), .ZN(new_n1004));
  AOI22_X1  g818(.A1(new_n992), .A2(new_n993), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(G900), .ZN(new_n1006));
  OAI21_X1  g820(.A(G953), .B1(new_n425), .B2(new_n1006), .ZN(new_n1007));
  OR2_X1    g821(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n992), .A2(new_n993), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1010));
  AND4_X1   g824(.A1(KEYINPUT126), .A2(new_n1009), .A3(new_n1007), .A4(new_n1010), .ZN(new_n1011));
  AOI21_X1  g825(.A(KEYINPUT126), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1008), .B1(new_n1011), .B2(new_n1012), .ZN(G72));
  NAND3_X1  g827(.A1(new_n1001), .A2(new_n891), .A3(new_n1002), .ZN(new_n1014));
  XOR2_X1   g828(.A(new_n694), .B(KEYINPUT63), .Z(new_n1015));
  AOI211_X1 g829(.A(new_n265), .B(new_n301), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g830(.A1(new_n982), .A2(new_n985), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1017), .A2(new_n891), .ZN(new_n1018));
  AOI211_X1 g832(.A(new_n267), .B(new_n322), .C1(new_n1018), .C2(new_n1015), .ZN(new_n1019));
  AOI21_X1  g833(.A(KEYINPUT127), .B1(new_n322), .B2(new_n265), .ZN(new_n1020));
  XOR2_X1   g834(.A(new_n1020), .B(new_n288), .Z(new_n1021));
  AND3_X1   g835(.A1(new_n886), .A2(new_n1015), .A3(new_n1021), .ZN(new_n1022));
  NOR4_X1   g836(.A1(new_n1016), .A2(new_n920), .A3(new_n1019), .A4(new_n1022), .ZN(G57));
endmodule


