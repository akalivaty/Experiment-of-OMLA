//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 0 1 1 1 0 1 0 0 0 1 1 1 1 1 0 1 0 1 1 1 1 0 0 1 0 1 0 1 1 1 1 1 0 1 1 0 1 0 1 0 0 0 0 1 0 1 0 1 1 1 0 1 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:55 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1274, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1342, new_n1343, new_n1344;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  XNOR2_X1  g0001(.A(new_n201), .B(KEYINPUT64), .ZN(new_n202));
  NOR2_X1   g0002(.A1(new_n202), .A2(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  XNOR2_X1  g0011(.A(KEYINPUT65), .B(G244), .ZN(new_n212));
  INV_X1    g0012(.A(G77), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G107), .B2(G264), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G68), .A2(G238), .B1(G97), .B2(G257), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G116), .A2(G270), .ZN(new_n218));
  NAND4_X1  g0018(.A1(new_n215), .A2(new_n216), .A3(new_n217), .A4(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n208), .B1(new_n214), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n221));
  OR2_X1    g0021(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n222));
  NOR2_X1   g0022(.A1(G58), .A2(G68), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(G50), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  AND2_X1   g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  NAND3_X1  g0027(.A1(new_n226), .A2(G20), .A3(new_n227), .ZN(new_n228));
  NAND4_X1  g0028(.A1(new_n211), .A2(new_n221), .A3(new_n222), .A4(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(KEYINPUT66), .Z(G361));
  XOR2_X1   g0030(.A(G238), .B(G244), .Z(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G226), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n235), .B(new_n238), .Z(G358));
  XOR2_X1   g0039(.A(G68), .B(G77), .Z(new_n240));
  XOR2_X1   g0040(.A(G50), .B(G58), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G351));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(G1), .A2(G13), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  OAI21_X1  g0049(.A(KEYINPUT23), .B1(new_n206), .B2(G107), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT23), .ZN(new_n251));
  INV_X1    g0051(.A(G107), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n251), .A2(new_n252), .A3(G20), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n206), .A2(G33), .A3(G116), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n250), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT87), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n255), .B(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT3), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n262), .A2(new_n206), .A3(G87), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(KEYINPUT22), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT22), .ZN(new_n265));
  NAND4_X1  g0065(.A1(new_n262), .A2(new_n265), .A3(new_n206), .A4(G87), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT24), .ZN(new_n268));
  AND3_X1   g0068(.A1(new_n257), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n268), .B1(new_n257), .B2(new_n267), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n249), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  AOI211_X1 g0073(.A(new_n249), .B(new_n273), .C1(new_n205), .C2(G33), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT25), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n275), .B1(new_n272), .B2(G107), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n273), .A2(KEYINPUT25), .A3(new_n252), .ZN(new_n277));
  AOI22_X1  g0077(.A1(new_n274), .A2(G107), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n271), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT88), .ZN(new_n280));
  AND2_X1   g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  NOR2_X1   g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  OAI211_X1 g0082(.A(G257), .B(G1698), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G1698), .ZN(new_n284));
  OAI211_X1 g0084(.A(G250), .B(new_n284), .C1(new_n281), .C2(new_n282), .ZN(new_n285));
  INV_X1    g0085(.A(G294), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n283), .B(new_n285), .C1(new_n259), .C2(new_n286), .ZN(new_n287));
  AND2_X1   g0087(.A1(G33), .A2(G41), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n288), .A2(new_n248), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT5), .B(G41), .ZN(new_n290));
  INV_X1    g0090(.A(G45), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n291), .A2(G1), .ZN(new_n292));
  NAND2_X1  g0092(.A1(G33), .A2(G41), .ZN(new_n293));
  AOI22_X1  g0093(.A1(new_n290), .A2(new_n292), .B1(new_n227), .B2(new_n293), .ZN(new_n294));
  AOI22_X1  g0094(.A1(new_n287), .A2(new_n289), .B1(G264), .B2(new_n294), .ZN(new_n295));
  AND2_X1   g0095(.A1(KEYINPUT5), .A2(G41), .ZN(new_n296));
  NOR2_X1   g0096(.A1(KEYINPUT5), .A2(G41), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n292), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  OAI21_X1  g0098(.A(G274), .B1(new_n288), .B2(new_n248), .ZN(new_n299));
  OAI21_X1  g0099(.A(KEYINPUT81), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G274), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n301), .B1(new_n227), .B2(new_n293), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT81), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n302), .A2(new_n303), .A3(new_n290), .A4(new_n292), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n300), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n295), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G179), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n280), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n295), .A2(KEYINPUT88), .A3(G179), .A4(new_n305), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n306), .A2(G169), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n279), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n306), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(G190), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n306), .A2(G200), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n271), .A2(new_n314), .A3(new_n278), .A4(new_n315), .ZN(new_n316));
  AND2_X1   g0116(.A1(new_n312), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT68), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n319));
  NOR3_X1   g0119(.A1(new_n299), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n319), .ZN(new_n321));
  AOI21_X1  g0121(.A(KEYINPUT68), .B1(new_n302), .B2(new_n321), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n227), .A2(new_n293), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n319), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n323), .B1(G226), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n262), .A2(new_n284), .ZN(new_n328));
  INV_X1    g0128(.A(G222), .ZN(new_n329));
  OAI22_X1  g0129(.A1(new_n328), .A2(new_n329), .B1(new_n213), .B2(new_n262), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n284), .B1(new_n260), .B2(new_n261), .ZN(new_n331));
  XOR2_X1   g0131(.A(new_n331), .B(KEYINPUT69), .Z(new_n332));
  AOI21_X1  g0132(.A(new_n330), .B1(new_n332), .B2(G223), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n327), .B1(new_n333), .B2(new_n324), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n273), .A2(new_n249), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n205), .A2(G20), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n335), .A2(G50), .A3(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G50), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n273), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  XNOR2_X1  g0140(.A(KEYINPUT8), .B(G58), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n206), .A2(G33), .ZN(new_n342));
  INV_X1    g0142(.A(G150), .ZN(new_n343));
  NOR2_X1   g0143(.A1(G20), .A2(G33), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  OAI22_X1  g0145(.A1(new_n341), .A2(new_n342), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n202), .A2(G20), .B1(new_n346), .B2(KEYINPUT70), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n347), .B1(KEYINPUT70), .B2(new_n346), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n340), .B1(new_n348), .B2(new_n249), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n334), .A2(G200), .B1(new_n349), .B2(KEYINPUT9), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(G190), .ZN(new_n352));
  OAI22_X1  g0152(.A1(new_n334), .A2(new_n352), .B1(new_n349), .B2(KEYINPUT9), .ZN(new_n353));
  OAI21_X1  g0153(.A(KEYINPUT10), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n353), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT10), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n355), .A2(new_n356), .A3(new_n350), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(G169), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n349), .B1(new_n334), .B2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT71), .ZN(new_n361));
  OR2_X1    g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT72), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n363), .B1(new_n334), .B2(G179), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n360), .A2(new_n361), .ZN(new_n365));
  OR3_X1    g0165(.A1(new_n334), .A2(new_n363), .A3(G179), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n362), .A2(new_n364), .A3(new_n365), .A4(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n318), .B1(new_n299), .B2(new_n319), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n302), .A2(KEYINPUT68), .A3(new_n321), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n370), .B1(new_n212), .B2(new_n325), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(G232), .ZN(new_n373));
  OAI22_X1  g0173(.A1(new_n328), .A2(new_n373), .B1(new_n252), .B2(new_n262), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n374), .B1(new_n332), .B2(G238), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n372), .B1(new_n375), .B2(new_n324), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G200), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(G87), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(KEYINPUT15), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT15), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(G87), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  OAI22_X1  g0185(.A1(new_n385), .A2(new_n342), .B1(new_n206), .B2(new_n213), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n341), .A2(new_n345), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n249), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n249), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n389), .A2(KEYINPUT73), .A3(new_n272), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT73), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(new_n273), .B2(new_n249), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n390), .A2(new_n392), .A3(G77), .A4(new_n336), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n388), .B(new_n393), .C1(G77), .C2(new_n272), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(new_n376), .B2(new_n352), .ZN(new_n396));
  OR2_X1    g0196(.A1(new_n379), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n377), .A2(new_n307), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n395), .B1(new_n376), .B2(new_n359), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n358), .A2(new_n367), .A3(new_n397), .A4(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT13), .ZN(new_n402));
  OAI211_X1 g0202(.A(G226), .B(new_n284), .C1(new_n281), .C2(new_n282), .ZN(new_n403));
  NAND2_X1  g0203(.A1(G33), .A2(G97), .ZN(new_n404));
  AND2_X1   g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT74), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n406), .B1(new_n331), .B2(G232), .ZN(new_n407));
  OAI211_X1 g0207(.A(G232), .B(G1698), .C1(new_n281), .C2(new_n282), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n408), .A2(KEYINPUT74), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n405), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n289), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n368), .A2(new_n369), .B1(new_n326), .B2(G238), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n402), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n408), .A2(KEYINPUT74), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n262), .A2(new_n406), .A3(G232), .A4(G1698), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n324), .B1(new_n416), .B2(new_n405), .ZN(new_n417));
  INV_X1    g0217(.A(G238), .ZN(new_n418));
  OAI22_X1  g0218(.A1(new_n320), .A2(new_n322), .B1(new_n418), .B2(new_n325), .ZN(new_n419));
  NOR3_X1   g0219(.A1(new_n417), .A2(KEYINPUT13), .A3(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(G169), .B1(new_n413), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT14), .ZN(new_n422));
  OAI21_X1  g0222(.A(KEYINPUT13), .B1(new_n417), .B2(new_n419), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n403), .A2(new_n404), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n424), .B1(new_n415), .B2(new_n414), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n412), .B(new_n402), .C1(new_n425), .C2(new_n324), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n423), .A2(new_n426), .A3(G179), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n423), .A2(new_n426), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT14), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n428), .A2(new_n429), .A3(G169), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n422), .A2(new_n427), .A3(new_n430), .ZN(new_n431));
  OAI22_X1  g0231(.A1(new_n342), .A2(new_n213), .B1(new_n206), .B2(G68), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT75), .ZN(new_n433));
  AOI22_X1  g0233(.A1(new_n432), .A2(new_n433), .B1(G50), .B2(new_n344), .ZN(new_n434));
  OAI221_X1 g0234(.A(KEYINPUT75), .B1(new_n206), .B2(G68), .C1(new_n342), .C2(new_n213), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n436), .A2(KEYINPUT11), .A3(new_n249), .ZN(new_n437));
  INV_X1    g0237(.A(G68), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n273), .A2(new_n438), .ZN(new_n439));
  XNOR2_X1  g0239(.A(new_n439), .B(KEYINPUT12), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n390), .A2(new_n392), .A3(G68), .A4(new_n336), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n389), .B1(new_n434), .B2(new_n435), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n442), .B1(new_n443), .B2(KEYINPUT11), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT76), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n423), .A2(new_n426), .A3(G190), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(new_n445), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n378), .B1(new_n423), .B2(new_n426), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n447), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n428), .A2(G200), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n452), .A2(KEYINPUT76), .A3(new_n448), .A4(new_n445), .ZN(new_n453));
  AOI22_X1  g0253(.A1(new_n431), .A2(new_n446), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  XNOR2_X1  g0255(.A(G58), .B(G68), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n456), .A2(G20), .B1(G159), .B2(new_n344), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n260), .A2(new_n206), .A3(new_n261), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT7), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(KEYINPUT77), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT77), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(KEYINPUT7), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(G68), .B1(new_n458), .B2(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n281), .A2(new_n282), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n459), .B1(new_n465), .B2(new_n206), .ZN(new_n466));
  OAI211_X1 g0266(.A(KEYINPUT16), .B(new_n457), .C1(new_n464), .C2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(G58), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n468), .A2(new_n438), .ZN(new_n469));
  OAI21_X1  g0269(.A(G20), .B1(new_n469), .B2(new_n223), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n344), .A2(G159), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n260), .A2(KEYINPUT7), .A3(new_n206), .A4(new_n261), .ZN(new_n473));
  NOR3_X1   g0273(.A1(new_n281), .A2(new_n282), .A3(G20), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n473), .B1(new_n474), .B2(new_n463), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n472), .B1(new_n475), .B2(G68), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n249), .B(new_n467), .C1(new_n476), .C2(KEYINPUT16), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n341), .B1(new_n205), .B2(G20), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n478), .A2(new_n335), .B1(new_n273), .B2(new_n341), .ZN(new_n479));
  INV_X1    g0279(.A(G226), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(G1698), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n481), .B1(G223), .B2(G1698), .ZN(new_n482));
  OAI22_X1  g0282(.A1(new_n482), .A2(new_n465), .B1(new_n259), .B2(new_n380), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n483), .A2(new_n289), .B1(new_n326), .B2(G232), .ZN(new_n484));
  XNOR2_X1  g0284(.A(KEYINPUT78), .B(G190), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n484), .A2(new_n485), .A3(new_n370), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n324), .A2(G232), .A3(new_n319), .ZN(new_n487));
  NOR2_X1   g0287(.A1(G223), .A2(G1698), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n488), .B1(new_n480), .B2(G1698), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n489), .A2(new_n262), .B1(G33), .B2(G87), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n487), .B1(new_n490), .B2(new_n324), .ZN(new_n491));
  OAI21_X1  g0291(.A(G200), .B1(new_n491), .B2(new_n323), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n477), .A2(new_n479), .A3(new_n486), .A4(new_n492), .ZN(new_n493));
  XNOR2_X1  g0293(.A(new_n493), .B(KEYINPUT17), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n477), .A2(new_n479), .ZN(new_n495));
  OAI21_X1  g0295(.A(G169), .B1(new_n491), .B2(new_n323), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n484), .A2(G179), .A3(new_n370), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT18), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n477), .A2(new_n479), .B1(new_n496), .B2(new_n497), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(KEYINPUT18), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  AND2_X1   g0304(.A1(new_n494), .A2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  NOR3_X1   g0306(.A1(new_n401), .A2(new_n455), .A3(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(G97), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n508), .A2(new_n252), .A3(KEYINPUT6), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n509), .B1(KEYINPUT6), .B2(new_n508), .ZN(new_n510));
  XOR2_X1   g0310(.A(KEYINPUT79), .B(G107), .Z(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g0312(.A(KEYINPUT79), .B(G107), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n513), .B(new_n509), .C1(KEYINPUT6), .C2(new_n508), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n512), .A2(new_n514), .A3(G20), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n344), .A2(G77), .ZN(new_n516));
  XNOR2_X1  g0316(.A(KEYINPUT77), .B(KEYINPUT7), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n458), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n252), .B1(new_n518), .B2(new_n473), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n515), .B(new_n516), .C1(new_n519), .C2(KEYINPUT80), .ZN(new_n520));
  AND2_X1   g0320(.A1(new_n519), .A2(KEYINPUT80), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n249), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n272), .A2(G97), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n523), .B1(new_n274), .B2(G97), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  AND2_X1   g0325(.A1(KEYINPUT4), .A2(G244), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n284), .B(new_n526), .C1(new_n281), .C2(new_n282), .ZN(new_n527));
  NAND2_X1  g0327(.A1(G33), .A2(G283), .ZN(new_n528));
  INV_X1    g0328(.A(G244), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n529), .B1(new_n260), .B2(new_n261), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n527), .B(new_n528), .C1(new_n530), .C2(KEYINPUT4), .ZN(new_n531));
  OAI21_X1  g0331(.A(G250), .B1(new_n281), .B2(new_n282), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n284), .B1(new_n532), .B2(KEYINPUT4), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n289), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n300), .A2(new_n304), .B1(new_n294), .B2(G257), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT82), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n294), .A2(G257), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n305), .A2(new_n536), .A3(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n352), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n378), .B1(new_n537), .B2(new_n539), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n525), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n206), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n380), .A2(new_n508), .A3(new_n252), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n206), .B(G68), .C1(new_n281), .C2(new_n282), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT19), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n549), .B1(new_n342), .B2(new_n508), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n547), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n249), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n384), .A2(new_n272), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(KEYINPUT85), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT85), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n552), .A2(new_n557), .A3(new_n554), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n418), .A2(new_n284), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n529), .A2(G1698), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n560), .B(new_n561), .C1(new_n281), .C2(new_n282), .ZN(new_n562));
  NAND2_X1  g0362(.A1(G33), .A2(G116), .ZN(new_n563));
  AND3_X1   g0363(.A1(new_n562), .A2(KEYINPUT84), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(KEYINPUT84), .B1(new_n562), .B2(new_n563), .ZN(new_n565));
  NOR3_X1   g0365(.A1(new_n564), .A2(new_n565), .A3(new_n324), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT83), .ZN(new_n567));
  INV_X1    g0367(.A(new_n292), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n567), .B1(new_n299), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n302), .A2(KEYINPUT83), .A3(new_n292), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n568), .A2(new_n324), .A3(G250), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OAI21_X1  g0373(.A(G200), .B1(new_n566), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n274), .A2(G87), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n562), .A2(new_n563), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT84), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n562), .A2(KEYINPUT84), .A3(new_n563), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n578), .A2(new_n289), .A3(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n572), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n581), .B1(new_n569), .B2(new_n570), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n580), .A2(G190), .A3(new_n582), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n559), .A2(new_n574), .A3(new_n575), .A4(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n274), .A2(new_n384), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n557), .B1(new_n552), .B2(new_n554), .ZN(new_n586));
  AOI211_X1 g0386(.A(KEYINPUT85), .B(new_n553), .C1(new_n551), .C2(new_n249), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n359), .B1(new_n566), .B2(new_n573), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n580), .A2(new_n307), .A3(new_n582), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n584), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(G169), .B1(new_n537), .B2(new_n539), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n305), .A2(new_n538), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(KEYINPUT82), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n535), .A2(new_n536), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n595), .A2(G179), .A3(new_n596), .A4(new_n534), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n593), .A2(new_n597), .B1(new_n522), .B2(new_n524), .ZN(new_n598));
  NOR3_X1   g0398(.A1(new_n543), .A2(new_n592), .A3(new_n598), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n300), .A2(new_n304), .B1(new_n294), .B2(G270), .ZN(new_n600));
  OAI211_X1 g0400(.A(G264), .B(G1698), .C1(new_n281), .C2(new_n282), .ZN(new_n601));
  OAI211_X1 g0401(.A(G257), .B(new_n284), .C1(new_n281), .C2(new_n282), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n260), .A2(G303), .A3(new_n261), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n289), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n600), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n606), .A2(new_n307), .ZN(new_n607));
  INV_X1    g0407(.A(G116), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n608), .B1(new_n205), .B2(G33), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n390), .A2(new_n392), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n273), .A2(new_n608), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n247), .A2(new_n248), .B1(G20), .B2(new_n608), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n528), .B(new_n206), .C1(G33), .C2(new_n508), .ZN(new_n613));
  AOI21_X1  g0413(.A(KEYINPUT20), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n612), .A2(KEYINPUT20), .A3(new_n613), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n610), .B(new_n611), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n607), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n359), .B1(new_n600), .B2(new_n605), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT21), .ZN(new_n619));
  AND3_X1   g0419(.A1(new_n618), .A2(new_n619), .A3(new_n616), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n619), .B1(new_n618), .B2(new_n616), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n617), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n616), .B1(G200), .B2(new_n606), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n294), .A2(G270), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n305), .A2(new_n605), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n485), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT86), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n623), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n623), .A2(new_n626), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(KEYINPUT86), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n622), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  AND4_X1   g0431(.A1(new_n317), .A2(new_n507), .A3(new_n599), .A4(new_n631), .ZN(G372));
  INV_X1    g0432(.A(new_n367), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n400), .B1(new_n451), .B2(new_n453), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n430), .A2(new_n427), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n429), .B1(new_n428), .B2(G169), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n446), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n494), .B1(new_n634), .B2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT92), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n495), .A2(KEYINPUT18), .A3(new_n498), .ZN(new_n641));
  AOI21_X1  g0441(.A(KEYINPUT18), .B1(new_n495), .B2(new_n498), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n501), .A2(KEYINPUT92), .A3(new_n503), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n639), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n633), .B1(new_n645), .B2(new_n358), .ZN(new_n646));
  INV_X1    g0446(.A(new_n507), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n593), .A2(new_n597), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n648), .A2(new_n584), .A3(new_n591), .A4(new_n525), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT26), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n598), .A2(KEYINPUT26), .A3(new_n591), .A4(new_n584), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n591), .A2(KEYINPUT90), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT90), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n588), .A2(new_n589), .A3(new_n655), .A4(new_n590), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n653), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(KEYINPUT91), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n657), .B1(new_n651), .B2(new_n652), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT91), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n622), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n312), .A2(KEYINPUT89), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT89), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n666), .B1(new_n279), .B2(new_n311), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n664), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n599), .A2(new_n316), .ZN(new_n669));
  AOI22_X1  g0469(.A1(new_n660), .A2(new_n663), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n646), .B1(new_n647), .B2(new_n670), .ZN(G369));
  NAND3_X1  g0471(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(G213), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(G343), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n616), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n678), .B(KEYINPUT93), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n630), .A2(new_n628), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n664), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n679), .B1(new_n681), .B2(KEYINPUT94), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n682), .B1(KEYINPUT94), .B2(new_n681), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n622), .A2(new_n679), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(G330), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n279), .A2(new_n677), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n317), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n279), .A2(new_n311), .A3(new_n677), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g0491(.A(new_n677), .B(KEYINPUT95), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  OR3_X1    g0493(.A1(new_n665), .A2(new_n667), .A3(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n664), .A2(new_n677), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n317), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  OR2_X1    g0497(.A1(new_n691), .A2(new_n697), .ZN(G399));
  INV_X1    g0498(.A(new_n209), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(G41), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n546), .A2(G116), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n701), .A2(G1), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n703), .B1(new_n225), .B2(new_n701), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT28), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n306), .B1(new_n537), .B2(new_n539), .ZN(new_n706));
  AOI21_X1  g0506(.A(G179), .B1(new_n600), .B2(new_n605), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT96), .ZN(new_n708));
  AND3_X1   g0508(.A1(new_n580), .A2(new_n708), .A3(new_n582), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n708), .B1(new_n580), .B2(new_n582), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n707), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT97), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI211_X1 g0513(.A(new_n707), .B(KEYINPUT97), .C1(new_n709), .C2(new_n710), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n706), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT30), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n625), .A2(new_n295), .A3(new_n580), .A4(new_n582), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n716), .B1(new_n597), .B2(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n580), .A2(new_n295), .A3(new_n582), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(new_n606), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n720), .A2(new_n540), .A3(KEYINPUT30), .A4(G179), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n677), .B1(new_n715), .B2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT31), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n599), .A2(new_n317), .A3(new_n631), .A4(new_n692), .ZN(new_n726));
  INV_X1    g0526(.A(new_n706), .ZN(new_n727));
  INV_X1    g0527(.A(new_n714), .ZN(new_n728));
  OAI21_X1  g0528(.A(KEYINPUT96), .B1(new_n566), .B2(new_n573), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n580), .A2(new_n708), .A3(new_n582), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(KEYINPUT97), .B1(new_n731), .B2(new_n707), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n727), .B1(new_n728), .B2(new_n732), .ZN(new_n733));
  AND2_X1   g0533(.A1(new_n718), .A2(new_n721), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n692), .A2(new_n724), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n725), .A2(new_n726), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G330), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT98), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n738), .A2(KEYINPUT98), .A3(G330), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT99), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n744), .B1(new_n670), .B2(new_n693), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT29), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n668), .A2(new_n316), .A3(new_n599), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n662), .B1(new_n653), .B2(new_n658), .ZN(new_n748));
  AOI211_X1 g0548(.A(KEYINPUT91), .B(new_n657), .C1(new_n651), .C2(new_n652), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n750), .A2(KEYINPUT99), .A3(new_n692), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n745), .A2(new_n746), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n664), .A2(new_n312), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n669), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n677), .B1(new_n754), .B2(new_n661), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(KEYINPUT29), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n743), .B1(new_n752), .B2(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n705), .B1(new_n757), .B2(G1), .ZN(G364));
  AOI21_X1  g0558(.A(new_n248), .B1(G20), .B2(new_n359), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n206), .A2(G179), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n760), .A2(G190), .A3(G200), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G87), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(new_n262), .ZN(new_n764));
  OR2_X1    g0564(.A1(new_n764), .A2(KEYINPUT102), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(KEYINPUT102), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n760), .A2(new_n352), .A3(G200), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(new_n252), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n352), .A2(G179), .A3(G200), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n206), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G97), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n765), .A2(new_n766), .A3(new_n769), .A4(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(G20), .A2(G179), .ZN(new_n775));
  XOR2_X1   g0575(.A(new_n775), .B(KEYINPUT100), .Z(new_n776));
  NAND3_X1  g0576(.A1(new_n776), .A2(new_n352), .A3(G200), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n776), .A2(new_n352), .A3(new_n378), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI22_X1  g0580(.A1(G68), .A2(new_n778), .B1(new_n780), .B2(G77), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n760), .A2(new_n352), .A3(new_n378), .ZN(new_n782));
  INV_X1    g0582(.A(G159), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT32), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n776), .A2(G200), .A3(new_n485), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n781), .B(new_n785), .C1(new_n338), .C2(new_n786), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n776), .A2(new_n378), .A3(new_n485), .ZN(new_n788));
  AND2_X1   g0588(.A1(new_n788), .A2(KEYINPUT101), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n788), .A2(KEYINPUT101), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  AOI211_X1 g0592(.A(new_n774), .B(new_n787), .C1(G58), .C2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(G303), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n465), .B1(new_n761), .B2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n767), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n795), .B1(G283), .B2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n782), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n772), .A2(G294), .B1(new_n798), .B2(G329), .ZN(new_n799));
  INV_X1    g0599(.A(G326), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n797), .B(new_n799), .C1(new_n800), .C2(new_n786), .ZN(new_n801));
  INV_X1    g0601(.A(G311), .ZN(new_n802));
  XOR2_X1   g0602(.A(KEYINPUT33), .B(G317), .Z(new_n803));
  OAI22_X1  g0603(.A1(new_n802), .A2(new_n779), .B1(new_n777), .B2(new_n803), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n801), .B(new_n804), .C1(new_n792), .C2(G322), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n759), .B1(new_n793), .B2(new_n805), .ZN(new_n806));
  AND2_X1   g0606(.A1(new_n206), .A2(G13), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n205), .B1(new_n807), .B2(G45), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n700), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n209), .A2(G116), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n699), .A2(new_n262), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(G45), .B2(new_n225), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(G45), .B2(new_n242), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n699), .A2(new_n465), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n812), .B(new_n815), .C1(G355), .C2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(G13), .A2(G33), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n820), .A2(G20), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(new_n759), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n811), .B1(new_n818), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n821), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n806), .B(new_n823), .C1(new_n685), .C2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n810), .B1(new_n685), .B2(G330), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n685), .A2(G330), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n825), .B1(new_n827), .B2(new_n828), .ZN(G396));
  INV_X1    g0629(.A(new_n677), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n379), .A2(new_n396), .B1(new_n395), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(new_n400), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n398), .A2(new_n399), .A3(new_n830), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n745), .A2(new_n751), .A3(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n834), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n750), .A2(new_n692), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n743), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n840), .B(KEYINPUT106), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n810), .B1(new_n838), .B2(new_n839), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n465), .B1(new_n761), .B2(new_n252), .ZN(new_n844));
  XOR2_X1   g0644(.A(new_n844), .B(KEYINPUT104), .Z(new_n845));
  NOR2_X1   g0645(.A1(new_n767), .A2(new_n380), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n773), .B1(new_n802), .B2(new_n782), .ZN(new_n847));
  NOR3_X1   g0647(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n608), .A2(new_n779), .B1(new_n786), .B2(new_n794), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(G283), .B2(new_n778), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n848), .B(new_n850), .C1(new_n286), .C2(new_n791), .ZN(new_n851));
  INV_X1    g0651(.A(new_n786), .ZN(new_n852));
  AOI22_X1  g0652(.A1(G137), .A2(new_n852), .B1(new_n778), .B2(G150), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n783), .B2(new_n779), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n854), .B1(G143), .B2(new_n792), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(KEYINPUT34), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n767), .A2(new_n438), .ZN(new_n857));
  INV_X1    g0657(.A(G132), .ZN(new_n858));
  OAI221_X1 g0658(.A(new_n262), .B1(new_n761), .B2(new_n338), .C1(new_n858), .C2(new_n782), .ZN(new_n859));
  AOI211_X1 g0659(.A(new_n857), .B(new_n859), .C1(G58), .C2(new_n772), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n856), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n855), .A2(KEYINPUT34), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n851), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT105), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n863), .A2(new_n864), .ZN(new_n867));
  INV_X1    g0667(.A(new_n759), .ZN(new_n868));
  NOR3_X1   g0668(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n759), .A2(new_n819), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n810), .B1(G77), .B2(new_n871), .ZN(new_n872));
  XOR2_X1   g0672(.A(new_n872), .B(KEYINPUT103), .Z(new_n873));
  OAI21_X1  g0673(.A(new_n873), .B1(new_n836), .B2(new_n820), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n843), .B1(new_n869), .B2(new_n874), .ZN(G384));
  NOR3_X1   g0675(.A1(new_n248), .A2(new_n206), .A3(new_n608), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n512), .A2(new_n514), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT35), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n876), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n880), .B1(new_n879), .B2(new_n878), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n881), .B(KEYINPUT36), .ZN(new_n882));
  OR3_X1    g0682(.A1(new_n225), .A2(new_n213), .A3(new_n469), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n338), .A2(G68), .ZN(new_n884));
  AOI211_X1 g0684(.A(new_n205), .B(G13), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n438), .B1(new_n474), .B2(new_n517), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n458), .A2(KEYINPUT7), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n472), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n889), .A2(KEYINPUT16), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n467), .A2(new_n249), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n479), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n675), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n894), .B1(new_n494), .B2(new_n504), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n495), .A2(new_n893), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n499), .A2(new_n896), .A3(new_n493), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT37), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n892), .B1(new_n498), .B2(new_n893), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n900), .A2(KEYINPUT37), .A3(new_n493), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT38), .ZN(new_n903));
  OR3_X1    g0703(.A1(new_n895), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n479), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n389), .B1(new_n889), .B2(KEYINPUT16), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT16), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n438), .B1(new_n518), .B2(new_n473), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n907), .B1(new_n908), .B2(new_n472), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n905), .B1(new_n906), .B2(new_n909), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n493), .B(new_n640), .C1(new_n910), .C2(new_n675), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(KEYINPUT37), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n897), .ZN(new_n913));
  INV_X1    g0713(.A(new_n493), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n675), .B1(new_n477), .B2(new_n479), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n916), .A2(KEYINPUT92), .A3(KEYINPUT37), .A4(new_n499), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n913), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n643), .A2(new_n644), .A3(new_n494), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n918), .B1(new_n915), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n904), .B1(new_n920), .B2(KEYINPUT38), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n446), .A2(new_n677), .ZN(new_n922));
  INV_X1    g0722(.A(new_n431), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n451), .A2(new_n453), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT108), .B1(new_n454), .B2(new_n922), .ZN(new_n927));
  AND4_X1   g0727(.A1(KEYINPUT108), .A2(new_n924), .A3(new_n637), .A4(new_n922), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  OAI211_X1 g0729(.A(KEYINPUT31), .B(new_n677), .C1(new_n715), .C2(new_n722), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n725), .A2(new_n726), .A3(new_n930), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n921), .A2(new_n836), .A3(new_n929), .A4(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(KEYINPUT40), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n931), .A2(new_n836), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n924), .A2(new_n637), .A3(new_n922), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT108), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n454), .A2(KEYINPUT108), .A3(new_n922), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n925), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n934), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n903), .B1(new_n895), .B2(new_n902), .ZN(new_n941));
  AOI21_X1  g0741(.A(KEYINPUT40), .B1(new_n904), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n933), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT109), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n507), .A2(new_n931), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n945), .A2(new_n946), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n947), .A2(G330), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n638), .A2(new_n830), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n904), .A2(KEYINPUT39), .A3(new_n941), .ZN(new_n952));
  NOR3_X1   g0752(.A1(new_n895), .A2(new_n902), .A3(new_n903), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n919), .A2(new_n915), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n916), .A2(new_n499), .B1(new_n911), .B2(KEYINPUT37), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n896), .A2(new_n493), .ZN(new_n956));
  NOR4_X1   g0756(.A1(new_n956), .A2(new_n640), .A3(new_n898), .A4(new_n502), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n953), .B1(new_n959), .B2(new_n903), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n951), .B(new_n952), .C1(new_n960), .C2(KEYINPUT39), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n643), .A2(new_n644), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n675), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n904), .A2(new_n941), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n833), .B(KEYINPUT107), .Z(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n939), .B1(new_n837), .B2(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n964), .B1(new_n965), .B2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n752), .A2(new_n507), .A3(new_n756), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n646), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n970), .B(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n949), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(new_n205), .B2(new_n807), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n949), .A2(new_n973), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n886), .B1(new_n975), .B2(new_n976), .ZN(G367));
  OAI21_X1  g0777(.A(new_n822), .B1(new_n209), .B2(new_n385), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n978), .B1(new_n813), .B2(new_n238), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT111), .Z(new_n980));
  AOI22_X1  g0780(.A1(G283), .A2(new_n780), .B1(new_n852), .B2(G311), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n286), .B2(new_n777), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n761), .A2(new_n608), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT46), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n262), .B1(new_n798), .B2(G317), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n985), .B1(new_n508), .B2(new_n767), .C1(new_n252), .C2(new_n771), .ZN(new_n986));
  NOR3_X1   g0786(.A1(new_n982), .A2(new_n984), .A3(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n794), .B2(new_n791), .ZN(new_n988));
  INV_X1    g0788(.A(G137), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n262), .B1(new_n761), .B2(new_n468), .C1(new_n989), .C2(new_n782), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n772), .A2(G68), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n213), .B2(new_n767), .ZN(new_n992));
  AOI211_X1 g0792(.A(new_n990), .B(new_n992), .C1(G159), .C2(new_n778), .ZN(new_n993));
  AOI22_X1  g0793(.A1(G50), .A2(new_n780), .B1(new_n852), .B2(G143), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n993), .B(new_n994), .C1(new_n343), .C2(new_n791), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n988), .A2(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT47), .ZN(new_n997));
  AOI211_X1 g0797(.A(new_n811), .B(new_n980), .C1(new_n997), .C2(new_n759), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n559), .A2(new_n575), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(new_n677), .ZN(new_n1000));
  MUX2_X1   g0800(.A(new_n658), .B(new_n592), .S(new_n1000), .Z(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n998), .B1(new_n824), .B2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1003), .B(KEYINPUT112), .Z(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n541), .A2(new_n542), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n525), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n598), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n1008), .B(new_n1009), .C1(new_n1007), .C2(new_n692), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n598), .A2(new_n693), .ZN(new_n1011));
  AND2_X1   g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1012), .A2(new_n696), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT110), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1009), .B1(new_n1010), .B2(new_n312), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n1014), .A2(KEYINPUT42), .B1(new_n692), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(KEYINPUT42), .B2(new_n1014), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1002), .A2(KEYINPUT43), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1002), .A2(KEYINPUT43), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1017), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1019), .B1(new_n1017), .B2(new_n1020), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n691), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n1022), .A2(new_n1023), .B1(new_n1024), .B2(new_n1012), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1023), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1024), .A2(new_n1012), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1026), .A2(new_n1027), .A3(new_n1021), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1025), .A2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n697), .A2(new_n1012), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT45), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n697), .A2(new_n1012), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT44), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1032), .B(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1031), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(new_n691), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1024), .A2(new_n1031), .A3(new_n1034), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n690), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n696), .B1(new_n1039), .B2(new_n695), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(new_n686), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n757), .B1(new_n1038), .B2(new_n1041), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n700), .B(KEYINPUT41), .Z(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n809), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1005), .B1(new_n1029), .B2(new_n1045), .ZN(G387));
  INV_X1    g0846(.A(new_n1041), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n701), .B1(new_n757), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT114), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1050), .B(new_n1051), .C1(new_n757), .C2(new_n1047), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n771), .A2(new_n385), .B1(new_n782), .B2(new_n343), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n762), .A2(G77), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1054), .B(new_n262), .C1(new_n508), .C2(new_n767), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n341), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n1053), .B(new_n1055), .C1(new_n1056), .C2(new_n778), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(G68), .A2(new_n780), .B1(new_n852), .B2(G159), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1057), .B(new_n1058), .C1(new_n338), .C2(new_n791), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n262), .B1(new_n798), .B2(G326), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(G303), .A2(new_n780), .B1(new_n852), .B2(G322), .ZN(new_n1061));
  INV_X1    g0861(.A(G317), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1061), .B1(new_n802), .B2(new_n777), .C1(new_n791), .C2(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT48), .ZN(new_n1064));
  OR2_X1    g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n772), .A2(G283), .B1(new_n762), .B2(G294), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT49), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n1060), .B1(new_n608), .B2(new_n767), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1070));
  AND2_X1   g0870(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1059), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n759), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n816), .B1(G116), .B2(new_n546), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n235), .A2(new_n291), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1056), .A2(new_n338), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT50), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n702), .B(new_n291), .C1(new_n438), .C2(new_n213), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n813), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n1074), .B1(G107), .B2(new_n209), .C1(new_n1075), .C2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n811), .B1(new_n1080), .B2(new_n822), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1073), .B(new_n1081), .C1(new_n1039), .C2(new_n824), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT113), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(new_n809), .B2(new_n1047), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1052), .A2(new_n1084), .ZN(G393));
  NAND2_X1  g0885(.A1(new_n1012), .A2(new_n821), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n791), .A2(new_n802), .B1(new_n1062), .B2(new_n786), .ZN(new_n1087));
  XOR2_X1   g0887(.A(new_n1087), .B(KEYINPUT52), .Z(new_n1088));
  AOI211_X1 g0888(.A(new_n262), .B(new_n768), .C1(G283), .C2(new_n762), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n772), .A2(G116), .B1(new_n798), .B2(G322), .ZN(new_n1090));
  AND2_X1   g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n1091), .B1(new_n286), .B2(new_n779), .C1(new_n794), .C2(new_n777), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n791), .A2(new_n783), .B1(new_n343), .B2(new_n786), .ZN(new_n1093));
  XOR2_X1   g0893(.A(new_n1093), .B(KEYINPUT51), .Z(new_n1094));
  AOI211_X1 g0894(.A(new_n465), .B(new_n846), .C1(G68), .C2(new_n762), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n772), .A2(G77), .B1(new_n798), .B2(G143), .ZN(new_n1096));
  AND2_X1   g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n1097), .B1(new_n338), .B2(new_n777), .C1(new_n341), .C2(new_n779), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n1088), .A2(new_n1092), .B1(new_n1094), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n759), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n813), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n822), .B1(new_n508), .B2(new_n209), .C1(new_n1101), .C2(new_n245), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1086), .A2(new_n1100), .A3(new_n810), .A4(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n1038), .B2(new_n808), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(KEYINPUT115), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT115), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1106), .B(new_n1103), .C1(new_n1038), .C2(new_n808), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n757), .A2(new_n1047), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n700), .B1(new_n1109), .B2(new_n1038), .ZN(new_n1110));
  AND2_X1   g0910(.A1(new_n1038), .A2(new_n1109), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1108), .B1(new_n1110), .B2(new_n1111), .ZN(G390));
  AOI22_X1  g0912(.A1(G97), .A2(new_n780), .B1(new_n778), .B2(G107), .ZN(new_n1113));
  INV_X1    g0913(.A(G283), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1113), .B1(new_n1114), .B2(new_n786), .ZN(new_n1115));
  XOR2_X1   g0915(.A(new_n1115), .B(KEYINPUT117), .Z(new_n1116));
  AOI22_X1  g0916(.A1(new_n772), .A2(G77), .B1(new_n798), .B2(G294), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n857), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1117), .A2(new_n465), .A3(new_n763), .A4(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(new_n792), .B2(G116), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n465), .B1(new_n798), .B2(G125), .ZN(new_n1121));
  OAI221_X1 g0921(.A(new_n1121), .B1(new_n338), .B2(new_n767), .C1(new_n783), .C2(new_n771), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(KEYINPUT54), .B(G143), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(G128), .A2(new_n852), .B1(new_n780), .B2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(new_n989), .B2(new_n777), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT53), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1127), .B1(new_n761), .B2(new_n343), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n762), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n1122), .B(new_n1126), .C1(new_n1128), .C2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n792), .A2(G132), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n1116), .A2(new_n1120), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n810), .B1(new_n1056), .B2(new_n871), .C1(new_n1132), .C2(new_n868), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n952), .B1(new_n960), .B2(KEYINPUT39), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1133), .B1(new_n1134), .B2(new_n819), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT118), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1134), .B1(new_n968), .B2(new_n951), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n834), .B1(new_n741), .B2(new_n742), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(new_n929), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n966), .B1(new_n755), .B2(new_n836), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n950), .B(new_n921), .C1(new_n1141), .C2(new_n939), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1138), .A2(new_n1140), .A3(new_n1142), .ZN(new_n1143));
  AND2_X1   g0943(.A1(new_n1138), .A2(new_n1142), .ZN(new_n1144));
  INV_X1    g0944(.A(G330), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n934), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n929), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1143), .B1(new_n1144), .B2(new_n1147), .ZN(new_n1148));
  OAI211_X1 g0948(.A(KEYINPUT119), .B(new_n1137), .C1(new_n1148), .C2(new_n808), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT119), .ZN(new_n1150));
  AND3_X1   g0950(.A1(new_n1138), .A2(new_n1140), .A3(new_n1142), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1147), .B1(new_n1138), .B2(new_n1142), .ZN(new_n1152));
  NOR3_X1   g0952(.A1(new_n1151), .A2(new_n1152), .A3(new_n808), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1150), .B1(new_n1153), .B2(new_n1136), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n507), .A2(G330), .A3(new_n931), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n971), .A2(new_n646), .A3(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n837), .A2(new_n967), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n723), .A2(new_n724), .B1(new_n735), .B2(new_n736), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n740), .B(new_n1145), .C1(new_n1158), .C2(new_n726), .ZN(new_n1159));
  AOI21_X1  g0959(.A(KEYINPUT98), .B1(new_n738), .B2(G330), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n836), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1161), .A2(KEYINPUT116), .A3(new_n939), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n1147), .ZN(new_n1163));
  AOI21_X1  g0963(.A(KEYINPUT116), .B1(new_n1161), .B2(new_n939), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1157), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1141), .B1(new_n929), .B2(new_n1146), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(new_n929), .B2(new_n1139), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1156), .B1(new_n1165), .B2(new_n1168), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n700), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT116), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1172), .B1(new_n1139), .B2(new_n929), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1173), .A2(new_n1162), .A3(new_n1147), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1167), .B1(new_n1174), .B2(new_n1157), .ZN(new_n1175));
  NOR3_X1   g0975(.A1(new_n1148), .A2(new_n1175), .A3(new_n1156), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1149), .B(new_n1154), .C1(new_n1171), .C2(new_n1176), .ZN(G378));
  INV_X1    g0977(.A(KEYINPUT57), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1165), .A2(new_n1168), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1156), .B1(new_n1179), .B2(new_n1170), .ZN(new_n1180));
  OR2_X1    g0980(.A1(new_n349), .A2(new_n675), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1181), .B(KEYINPUT55), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(new_n358), .B2(new_n367), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  XOR2_X1   g0984(.A(KEYINPUT120), .B(KEYINPUT56), .Z(new_n1185));
  NAND3_X1  g0985(.A1(new_n358), .A2(new_n367), .A3(new_n1182), .ZN(new_n1186));
  AND3_X1   g0986(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1185), .B1(new_n1184), .B2(new_n1186), .ZN(new_n1188));
  OR2_X1    g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(new_n944), .B2(G330), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n932), .A2(KEYINPUT40), .B1(new_n940), .B2(new_n942), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1192));
  NOR3_X1   g0992(.A1(new_n1191), .A2(new_n1145), .A3(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n970), .B1(new_n1190), .B2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1192), .B1(new_n1191), .B2(new_n1145), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT40), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(new_n940), .B2(new_n921), .ZN(new_n1197));
  AND4_X1   g0997(.A1(new_n836), .A2(new_n942), .A3(new_n929), .A4(new_n931), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1189), .B(G330), .C1(new_n1197), .C2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1195), .A2(new_n1199), .A3(new_n969), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1194), .A2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1178), .B1(new_n1180), .B2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1156), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n1148), .B2(new_n1175), .ZN(new_n1204));
  AND3_X1   g1004(.A1(new_n1195), .A2(new_n969), .A3(new_n1199), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n969), .B1(new_n1195), .B2(new_n1199), .ZN(new_n1206));
  NOR3_X1   g1006(.A1(new_n1205), .A2(new_n1206), .A3(new_n1178), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n701), .B1(new_n1204), .B2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1202), .A2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1194), .A2(new_n809), .A3(new_n1200), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n468), .A2(new_n767), .B1(new_n782), .B2(new_n1114), .ZN(new_n1211));
  INV_X1    g1011(.A(G41), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n991), .A2(new_n1212), .A3(new_n465), .A4(new_n1054), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n1211), .B(new_n1213), .C1(new_n384), .C2(new_n780), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(G97), .A2(new_n778), .B1(new_n852), .B2(G116), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1214), .B(new_n1215), .C1(new_n252), .C2(new_n791), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT58), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n465), .A2(new_n1212), .ZN(new_n1218));
  AOI21_X1  g1018(.A(G50), .B1(new_n259), .B2(new_n1212), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n1216), .A2(new_n1217), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(G132), .A2(new_n778), .B1(new_n780), .B2(G137), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n852), .A2(G125), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n772), .A2(G150), .B1(new_n762), .B2(new_n1124), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1221), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(G128), .B2(new_n792), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(KEYINPUT59), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n796), .A2(G159), .ZN(new_n1228));
  AOI211_X1 g1028(.A(G33), .B(G41), .C1(new_n798), .C2(G124), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1227), .A2(new_n1228), .A3(new_n1229), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1226), .A2(KEYINPUT59), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1220), .B1(new_n1217), .B2(new_n1216), .C1(new_n1230), .C2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(new_n759), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n811), .B1(new_n338), .B2(new_n870), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1233), .B(new_n1234), .C1(new_n1192), .C2(new_n820), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1210), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1209), .A2(new_n1237), .ZN(G375));
  AOI21_X1  g1038(.A(new_n811), .B1(new_n438), .B2(new_n870), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n262), .B1(new_n761), .B2(new_n783), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(G58), .B2(new_n796), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n772), .A2(G50), .B1(new_n798), .B2(G128), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1241), .B(new_n1242), .C1(new_n343), .C2(new_n779), .ZN(new_n1243));
  XOR2_X1   g1043(.A(new_n1243), .B(KEYINPUT121), .Z(new_n1244));
  OAI22_X1  g1044(.A1(new_n858), .A2(new_n786), .B1(new_n777), .B2(new_n1123), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(new_n792), .B2(G137), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n792), .A2(G283), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n608), .A2(new_n777), .B1(new_n786), .B2(new_n286), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n779), .A2(new_n252), .ZN(new_n1249));
  OAI221_X1 g1049(.A(new_n465), .B1(new_n761), .B2(new_n508), .C1(new_n213), .C2(new_n767), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n771), .A2(new_n385), .B1(new_n782), .B2(new_n794), .ZN(new_n1251));
  NOR4_X1   g1051(.A1(new_n1248), .A2(new_n1249), .A3(new_n1250), .A4(new_n1251), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n1244), .A2(new_n1246), .B1(new_n1247), .B2(new_n1252), .ZN(new_n1253));
  OAI221_X1 g1053(.A(new_n1239), .B1(new_n868), .B2(new_n1253), .C1(new_n929), .C2(new_n820), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1255), .B1(new_n1179), .B2(new_n809), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1179), .A2(new_n1203), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1044), .B1(new_n1175), .B2(new_n1156), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1256), .B1(new_n1257), .B2(new_n1258), .ZN(G381));
  INV_X1    g1059(.A(G396), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1052), .A2(new_n1260), .A3(new_n1084), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1261), .A2(G384), .ZN(new_n1262));
  XOR2_X1   g1062(.A(new_n1262), .B(KEYINPUT122), .Z(new_n1263));
  NOR2_X1   g1063(.A1(new_n1153), .A2(new_n1136), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1264), .B1(new_n1171), .B2(new_n1176), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NOR3_X1   g1066(.A1(G387), .A2(G390), .A3(G381), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1263), .A2(new_n1266), .A3(new_n1267), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1268), .A2(G375), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT123), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NOR3_X1   g1071(.A1(new_n1268), .A2(KEYINPUT123), .A3(G375), .ZN(new_n1272));
  OR2_X1    g1072(.A1(new_n1271), .A2(new_n1272), .ZN(G407));
  NAND4_X1  g1073(.A1(new_n1266), .A2(new_n1209), .A3(new_n676), .A4(new_n1237), .ZN(new_n1274));
  OAI211_X1 g1074(.A(G213), .B(new_n1274), .C1(new_n1271), .C2(new_n1272), .ZN(G409));
  INV_X1    g1075(.A(new_n1029), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1045), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1004), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  OAI21_X1  g1078(.A(G390), .B1(new_n1278), .B2(KEYINPUT126), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(G393), .A2(G396), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(new_n1261), .ZN(new_n1281));
  INV_X1    g1081(.A(G390), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT126), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1282), .A2(G387), .A3(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1279), .A2(new_n1281), .A3(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT125), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(G390), .A2(new_n1286), .ZN(new_n1287));
  OAI211_X1 g1087(.A(new_n1108), .B(KEYINPUT125), .C1(new_n1110), .C2(new_n1111), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1278), .A2(new_n1287), .A3(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(G387), .A2(G390), .A3(new_n1286), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1289), .A2(new_n1261), .A3(new_n1280), .A4(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1285), .A2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1209), .A2(G378), .A3(new_n1237), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT124), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1194), .A2(new_n1044), .A3(new_n1200), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1236), .B1(new_n1204), .B2(new_n1297), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1295), .B1(new_n1298), .B2(new_n1265), .ZN(new_n1299));
  OAI211_X1 g1099(.A(new_n1210), .B(new_n1235), .C1(new_n1180), .C2(new_n1296), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1148), .B1(new_n1175), .B2(new_n1156), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1301), .A2(new_n1302), .A3(new_n700), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1300), .A2(KEYINPUT124), .A3(new_n1303), .A4(new_n1264), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1294), .A2(new_n1299), .A3(new_n1304), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1169), .A2(new_n701), .ZN(new_n1306));
  NOR3_X1   g1106(.A1(new_n1179), .A2(KEYINPUT60), .A3(new_n1203), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT60), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1308), .B1(new_n1175), .B2(new_n1156), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1306), .B1(new_n1307), .B2(new_n1309), .ZN(new_n1310));
  AND3_X1   g1110(.A1(new_n1310), .A2(G384), .A3(new_n1256), .ZN(new_n1311));
  AOI21_X1  g1111(.A(G384), .B1(new_n1310), .B2(new_n1256), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n676), .A2(G213), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1305), .A2(new_n1313), .A3(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT62), .ZN(new_n1316));
  AND2_X1   g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT127), .ZN(new_n1318));
  AND3_X1   g1118(.A1(new_n1305), .A2(new_n1318), .A3(new_n1314), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1318), .B1(new_n1305), .B2(new_n1314), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1313), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1322), .A2(new_n1316), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1317), .B1(new_n1321), .B2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(G2897), .ZN(new_n1325));
  NOR2_X1   g1125(.A1(new_n1314), .A2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1313), .A2(new_n1326), .ZN(new_n1327));
  OAI22_X1  g1127(.A1(new_n1311), .A2(new_n1312), .B1(new_n1325), .B2(new_n1314), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1329), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT61), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1293), .B1(new_n1324), .B2(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1292), .A2(new_n1331), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1305), .A2(new_n1314), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1334), .B1(new_n1335), .B2(new_n1329), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1321), .A2(KEYINPUT63), .A3(new_n1313), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT63), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1315), .A2(new_n1338), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1336), .A2(new_n1337), .A3(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1333), .A2(new_n1340), .ZN(G405));
  NAND2_X1  g1141(.A1(G375), .A2(new_n1266), .ZN(new_n1342));
  AND2_X1   g1142(.A1(new_n1342), .A2(new_n1294), .ZN(new_n1343));
  XNOR2_X1  g1143(.A(new_n1343), .B(new_n1322), .ZN(new_n1344));
  XNOR2_X1  g1144(.A(new_n1344), .B(new_n1293), .ZN(G402));
endmodule


