//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 0 0 1 0 0 0 1 1 0 1 1 1 0 0 0 0 0 0 1 1 0 0 1 1 0 0 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0 0 0 0 1 0 1 1 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:43 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n444, new_n445, new_n446, new_n451, new_n453,
    new_n456, new_n457, new_n458, new_n459, new_n460, new_n461, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n492, new_n493,
    new_n494, new_n495, new_n496, new_n497, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n566, new_n568, new_n569, new_n570, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n628, new_n629, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n833, new_n834, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1136,
    new_n1137, new_n1138;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  XOR2_X1   g017(.A(KEYINPUT66), .B(G108), .Z(G238));
  INV_X1    g018(.A(G2072), .ZN(new_n444));
  INV_X1    g019(.A(G2078), .ZN(new_n445));
  NOR2_X1   g020(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g021(.A1(new_n446), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g022(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g023(.A(G452), .Z(G391));
  AND2_X1   g024(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g025(.A1(G7), .A2(G661), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g027(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT67), .ZN(G234));
  NAND3_X1  g029(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g030(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n456));
  XOR2_X1   g031(.A(KEYINPUT68), .B(KEYINPUT2), .Z(new_n457));
  XNOR2_X1  g032(.A(new_n456), .B(new_n457), .ZN(new_n458));
  NOR4_X1   g033(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT69), .Z(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n458), .A2(new_n461), .ZN(G325));
  INV_X1    g037(.A(G325), .ZN(G261));
  NAND2_X1  g038(.A1(new_n458), .A2(G2106), .ZN(new_n464));
  OR2_X1    g039(.A1(new_n464), .A2(KEYINPUT70), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(KEYINPUT70), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n461), .A2(G567), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  XNOR2_X1  g043(.A(new_n468), .B(KEYINPUT71), .ZN(G319));
  INV_X1    g044(.A(KEYINPUT73), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT72), .ZN(new_n471));
  INV_X1    g046(.A(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(KEYINPUT72), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G2105), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n470), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AND2_X1   g052(.A1(KEYINPUT72), .A2(G2104), .ZN(new_n478));
  NOR2_X1   g053(.A1(KEYINPUT72), .A2(G2104), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n470), .B(new_n476), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  OAI21_X1  g056(.A(G101), .B1(new_n477), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n473), .A2(KEYINPUT3), .A3(new_n474), .ZN(new_n483));
  OR2_X1    g058(.A1(new_n472), .A2(KEYINPUT3), .ZN(new_n484));
  NAND4_X1  g059(.A1(new_n483), .A2(G137), .A3(new_n476), .A4(new_n484), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n482), .A2(KEYINPUT74), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT74), .ZN(new_n487));
  INV_X1    g062(.A(G101), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n476), .B1(new_n478), .B2(new_n479), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(KEYINPUT73), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n488), .B1(new_n490), .B2(new_n480), .ZN(new_n491));
  INV_X1    g066(.A(new_n485), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n487), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  XNOR2_X1  g068(.A(KEYINPUT3), .B(G2104), .ZN(new_n494));
  AOI22_X1  g069(.A1(new_n494), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n495));
  OR2_X1    g070(.A1(new_n495), .A2(new_n476), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n486), .A2(new_n493), .A3(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G160));
  NAND3_X1  g073(.A1(new_n483), .A2(new_n476), .A3(new_n484), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G136), .ZN(new_n501));
  AND3_X1   g076(.A1(new_n483), .A2(G2105), .A3(new_n484), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G124), .ZN(new_n503));
  MUX2_X1   g078(.A(G100), .B(G112), .S(G2105), .Z(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G2104), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n501), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G162));
  MUX2_X1   g082(.A(G102), .B(G114), .S(G2105), .Z(new_n508));
  AOI22_X1  g083(.A1(new_n502), .A2(G126), .B1(G2104), .B2(new_n508), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n483), .A2(G138), .A3(new_n476), .A4(new_n484), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT75), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n510), .A2(new_n511), .A3(KEYINPUT4), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT4), .ZN(new_n513));
  NAND4_X1  g088(.A1(new_n494), .A2(new_n513), .A3(G138), .A4(new_n476), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n511), .B1(new_n510), .B2(KEYINPUT4), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n509), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(G164));
  AND2_X1   g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G543), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G50), .ZN(new_n524));
  OR2_X1    g099(.A1(new_n519), .A2(new_n520), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT5), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(new_n522), .ZN(new_n527));
  NAND2_X1  g102(.A1(KEYINPUT5), .A2(G543), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n525), .A2(new_n529), .ZN(new_n530));
  XOR2_X1   g105(.A(KEYINPUT76), .B(G88), .Z(new_n531));
  INV_X1    g106(.A(G651), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n529), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n533));
  OAI221_X1 g108(.A(new_n524), .B1(new_n530), .B2(new_n531), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT77), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n534), .A2(new_n535), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(G166));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT7), .ZN(new_n540));
  INV_X1    g115(.A(new_n523), .ZN(new_n541));
  INV_X1    g116(.A(G51), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AND2_X1   g118(.A1(new_n527), .A2(new_n528), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n525), .A2(G89), .ZN(new_n545));
  NAND2_X1  g120(.A1(G63), .A2(G651), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n543), .A2(new_n547), .ZN(G168));
  NAND2_X1  g123(.A1(G77), .A2(G543), .ZN(new_n549));
  INV_X1    g124(.A(G64), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n549), .B1(new_n544), .B2(new_n550), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n532), .B1(new_n551), .B2(KEYINPUT78), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n552), .B1(KEYINPUT78), .B2(new_n551), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n544), .A2(new_n521), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n554), .A2(G90), .B1(G52), .B2(new_n523), .ZN(new_n555));
  AND2_X1   g130(.A1(new_n553), .A2(new_n555), .ZN(G171));
  AOI22_X1  g131(.A1(new_n529), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n557));
  OR2_X1    g132(.A1(new_n557), .A2(KEYINPUT79), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(KEYINPUT79), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n558), .A2(G651), .A3(new_n559), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n554), .A2(G81), .B1(G43), .B2(new_n523), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT80), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(G153));
  AND3_X1   g140(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G36), .ZN(G176));
  XNOR2_X1  g142(.A(KEYINPUT81), .B(KEYINPUT8), .ZN(new_n568));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n568), .B(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n566), .A2(new_n570), .ZN(G188));
  NAND2_X1  g146(.A1(G78), .A2(G543), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n529), .B(KEYINPUT83), .ZN(new_n573));
  INV_X1    g148(.A(G65), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G651), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT82), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n523), .A2(new_n577), .A3(KEYINPUT9), .A4(G53), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT9), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n577), .A2(G53), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n541), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n554), .A2(G91), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n576), .A2(new_n578), .A3(new_n581), .A4(new_n582), .ZN(G299));
  XNOR2_X1  g158(.A(G171), .B(KEYINPUT84), .ZN(G301));
  INV_X1    g159(.A(G168), .ZN(G286));
  INV_X1    g160(.A(G166), .ZN(G303));
  OAI211_X1 g161(.A(G49), .B(G543), .C1(new_n519), .C2(new_n520), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n587), .B(KEYINPUT85), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(new_n589));
  OAI21_X1  g164(.A(G651), .B1(new_n529), .B2(G74), .ZN(new_n590));
  INV_X1    g165(.A(G87), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n530), .B2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n589), .A2(new_n593), .ZN(G288));
  NAND3_X1  g169(.A1(new_n525), .A2(G48), .A3(G543), .ZN(new_n595));
  INV_X1    g170(.A(G86), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n530), .B2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(G61), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n598), .B1(new_n527), .B2(new_n528), .ZN(new_n599));
  AND2_X1   g174(.A1(G73), .A2(G543), .ZN(new_n600));
  OAI21_X1  g175(.A(G651), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n597), .A2(new_n602), .ZN(new_n603));
  XOR2_X1   g178(.A(new_n603), .B(KEYINPUT86), .Z(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(G305));
  NAND2_X1  g180(.A1(new_n523), .A2(G47), .ZN(new_n606));
  INV_X1    g181(.A(G85), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(new_n530), .ZN(new_n608));
  AND2_X1   g183(.A1(new_n608), .A2(KEYINPUT87), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n608), .A2(KEYINPUT87), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n529), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n611));
  OAI22_X1  g186(.A1(new_n609), .A2(new_n610), .B1(new_n532), .B2(new_n611), .ZN(G290));
  NAND2_X1  g187(.A1(new_n554), .A2(G92), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT10), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n614), .B1(G54), .B2(new_n523), .ZN(new_n615));
  INV_X1    g190(.A(G66), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n573), .A2(new_n616), .ZN(new_n617));
  AND2_X1   g192(.A1(G79), .A2(G543), .ZN(new_n618));
  OAI21_X1  g193(.A(G651), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(G868), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(G301), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(new_n621), .ZN(G284));
  OAI21_X1  g199(.A(new_n622), .B1(new_n623), .B2(new_n621), .ZN(G321));
  MUX2_X1   g200(.A(G286), .B(G299), .S(new_n621), .Z(G297));
  MUX2_X1   g201(.A(G286), .B(G299), .S(new_n621), .Z(G280));
  INV_X1    g202(.A(new_n620), .ZN(new_n628));
  INV_X1    g203(.A(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(new_n629), .B2(G860), .ZN(G148));
  NAND2_X1  g205(.A1(new_n628), .A2(new_n629), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT88), .ZN(new_n632));
  MUX2_X1   g207(.A(new_n563), .B(new_n632), .S(G868), .Z(G323));
  XNOR2_X1  g208(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g209(.A1(new_n490), .A2(new_n480), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(new_n494), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(KEYINPUT12), .Z(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(KEYINPUT13), .Z(new_n638));
  INV_X1    g213(.A(G2100), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  MUX2_X1   g216(.A(G99), .B(G111), .S(G2105), .Z(new_n642));
  AOI22_X1  g217(.A1(new_n502), .A2(G123), .B1(G2104), .B2(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(G135), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n643), .B1(new_n644), .B2(new_n499), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(G2096), .Z(new_n646));
  NAND3_X1  g221(.A1(new_n640), .A2(new_n641), .A3(new_n646), .ZN(G156));
  INV_X1    g222(.A(KEYINPUT14), .ZN(new_n648));
  XOR2_X1   g223(.A(KEYINPUT15), .B(G2435), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2438), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2427), .ZN(new_n651));
  INV_X1    g226(.A(G2430), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n648), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n653), .B1(new_n652), .B2(new_n651), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2451), .B(G2454), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(KEYINPUT89), .B(KEYINPUT16), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G1341), .B(G1348), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n654), .A2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(G14), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n663), .B1(new_n654), .B2(new_n661), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT90), .ZN(G401));
  XOR2_X1   g241(.A(G2072), .B(G2078), .Z(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT17), .Z(new_n668));
  XNOR2_X1  g243(.A(G2067), .B(G2678), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT91), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n670), .A2(new_n667), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2084), .B(G2090), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT92), .ZN(new_n676));
  OR3_X1    g251(.A1(new_n668), .A2(new_n671), .A3(new_n674), .ZN(new_n677));
  NOR3_X1   g252(.A1(new_n670), .A2(new_n667), .A3(new_n674), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT18), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n676), .A2(new_n677), .A3(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(KEYINPUT93), .Z(new_n681));
  XOR2_X1   g256(.A(G2096), .B(G2100), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(G227));
  XNOR2_X1  g259(.A(G1956), .B(G2474), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT94), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1961), .B(G1966), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1971), .B(G1976), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT19), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT20), .Z(new_n693));
  NOR2_X1   g268(.A1(new_n686), .A2(new_n688), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n695), .A2(new_n691), .A3(new_n689), .ZN(new_n696));
  OAI211_X1 g271(.A(new_n693), .B(new_n696), .C1(new_n691), .C2(new_n695), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT95), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1991), .B(G1996), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1981), .B(G1986), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n700), .B(new_n703), .ZN(G229));
  NAND2_X1  g279(.A1(new_n628), .A2(G16), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G4), .B2(G16), .ZN(new_n706));
  INV_X1    g281(.A(G1348), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(G29), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G26), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT28), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n500), .A2(G140), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n502), .A2(G128), .ZN(new_n713));
  MUX2_X1   g288(.A(G104), .B(G116), .S(G2105), .Z(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G2104), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n712), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n711), .B1(new_n717), .B2(new_n709), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT100), .B(G2067), .Z(new_n719));
  AOI21_X1  g294(.A(new_n708), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(G16), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G19), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(new_n564), .B2(new_n721), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(G1341), .Z(new_n724));
  NOR2_X1   g299(.A1(new_n718), .A2(new_n719), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(new_n706), .B2(new_n707), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n720), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT101), .Z(new_n728));
  NOR2_X1   g303(.A1(G27), .A2(G29), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G164), .B2(G29), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(new_n445), .ZN(new_n731));
  AOI22_X1  g306(.A1(new_n494), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n732), .A2(new_n476), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n476), .A2(G103), .A3(G2104), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT102), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT25), .Z(new_n736));
  AOI211_X1 g311(.A(new_n733), .B(new_n736), .C1(G139), .C2(new_n500), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(G29), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G29), .B2(G33), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n739), .A2(new_n444), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT103), .Z(new_n741));
  NOR2_X1   g316(.A1(G29), .A2(G35), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(G162), .B2(G29), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT29), .Z(new_n744));
  INV_X1    g319(.A(G2090), .ZN(new_n745));
  INV_X1    g320(.A(G2084), .ZN(new_n746));
  AND2_X1   g321(.A1(KEYINPUT24), .A2(G34), .ZN(new_n747));
  NOR2_X1   g322(.A1(KEYINPUT24), .A2(G34), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n709), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(new_n497), .B2(new_n709), .ZN(new_n750));
  AOI22_X1  g325(.A1(new_n744), .A2(new_n745), .B1(new_n746), .B2(new_n750), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n741), .B(new_n751), .C1(new_n745), .C2(new_n744), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n721), .A2(G5), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G171), .B2(new_n721), .ZN(new_n754));
  AOI22_X1  g329(.A1(new_n739), .A2(new_n444), .B1(new_n754), .B2(G1961), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n721), .A2(G20), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT23), .Z(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G299), .B2(G16), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G1956), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT104), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT31), .B(G11), .ZN(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT30), .B(G28), .ZN(new_n762));
  AOI22_X1  g337(.A1(new_n760), .A2(new_n761), .B1(new_n762), .B2(new_n709), .ZN(new_n763));
  OAI221_X1 g338(.A(new_n763), .B1(new_n760), .B2(new_n761), .C1(new_n645), .C2(new_n709), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n721), .A2(G21), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G168), .B2(new_n721), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n764), .B1(new_n766), .B2(G1966), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n766), .A2(G1966), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT105), .ZN(new_n769));
  NAND4_X1  g344(.A1(new_n755), .A2(new_n759), .A3(new_n767), .A4(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n754), .A2(G1961), .ZN(new_n771));
  AOI22_X1  g346(.A1(G141), .A2(new_n500), .B1(new_n502), .B2(G129), .ZN(new_n772));
  NAND3_X1  g347(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT26), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n635), .B2(G105), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n777), .A2(new_n709), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n709), .B2(G32), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT27), .B(G1996), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n771), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OAI221_X1 g356(.A(new_n781), .B1(new_n746), .B2(new_n750), .C1(new_n779), .C2(new_n780), .ZN(new_n782));
  NOR3_X1   g357(.A1(new_n752), .A2(new_n770), .A3(new_n782), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n728), .A2(new_n731), .A3(new_n783), .ZN(new_n784));
  MUX2_X1   g359(.A(G24), .B(G290), .S(G16), .Z(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G1986), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n500), .A2(G131), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n502), .A2(G119), .ZN(new_n788));
  AND2_X1   g363(.A1(G107), .A2(G2105), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G95), .B2(new_n476), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n787), .B(new_n788), .C1(new_n472), .C2(new_n790), .ZN(new_n791));
  MUX2_X1   g366(.A(G25), .B(new_n791), .S(G29), .Z(new_n792));
  XOR2_X1   g367(.A(KEYINPUT35), .B(G1991), .Z(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n792), .B(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n786), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(G6), .A2(G16), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(new_n604), .B2(G16), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT32), .B(G1981), .Z(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n721), .A2(G22), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G166), .B2(new_n721), .ZN(new_n802));
  INV_X1    g377(.A(G1971), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n800), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(G16), .A2(G23), .ZN(new_n806));
  OR3_X1    g381(.A1(new_n588), .A2(new_n592), .A3(KEYINPUT96), .ZN(new_n807));
  OAI21_X1  g382(.A(KEYINPUT96), .B1(new_n588), .B2(new_n592), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n806), .B1(new_n809), .B2(G16), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT33), .B(G1976), .Z(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n805), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n796), .B1(new_n813), .B2(KEYINPUT34), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n805), .A2(new_n812), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT34), .ZN(new_n816));
  OAI21_X1  g391(.A(KEYINPUT97), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT97), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n813), .A2(new_n818), .A3(KEYINPUT34), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n814), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT99), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT98), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n823), .A2(KEYINPUT36), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n821), .A2(new_n822), .A3(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(KEYINPUT99), .B1(new_n820), .B2(new_n824), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT36), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n828), .B1(KEYINPUT98), .B2(new_n829), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n826), .A2(new_n823), .A3(KEYINPUT36), .A4(new_n827), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n784), .B1(new_n830), .B2(new_n831), .ZN(G311));
  NAND2_X1  g407(.A1(new_n830), .A2(new_n831), .ZN(new_n833));
  INV_X1    g408(.A(new_n784), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(G150));
  NAND2_X1  g410(.A1(new_n628), .A2(G559), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT38), .ZN(new_n837));
  XOR2_X1   g412(.A(KEYINPUT106), .B(G55), .Z(new_n838));
  INV_X1    g413(.A(G93), .ZN(new_n839));
  OAI22_X1  g414(.A1(new_n541), .A2(new_n838), .B1(new_n530), .B2(new_n839), .ZN(new_n840));
  AOI22_X1  g415(.A1(new_n529), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n841), .A2(new_n532), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n564), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n562), .A2(new_n843), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n837), .B(new_n847), .ZN(new_n848));
  OR2_X1    g423(.A1(new_n848), .A2(KEYINPUT39), .ZN(new_n849));
  INV_X1    g424(.A(G860), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n848), .A2(KEYINPUT39), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n843), .A2(new_n850), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT37), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n852), .A2(new_n854), .ZN(G145));
  XNOR2_X1  g430(.A(KEYINPUT109), .B(G37), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n637), .B(new_n791), .ZN(new_n858));
  MUX2_X1   g433(.A(G106), .B(G118), .S(G2105), .Z(new_n859));
  AOI22_X1  g434(.A1(new_n502), .A2(G130), .B1(G2104), .B2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(G142), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n860), .B1(new_n861), .B2(new_n499), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n858), .B(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n517), .B(new_n716), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n863), .B(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT108), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n737), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n776), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n865), .B(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n497), .B(KEYINPUT107), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n645), .B(new_n506), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n870), .B(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n857), .B1(new_n869), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n873), .B1(new_n872), .B2(new_n869), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g450(.A1(new_n844), .A2(G868), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n632), .B(new_n847), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n620), .B(G299), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT41), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n880), .B1(new_n878), .B2(new_n877), .ZN(new_n881));
  XOR2_X1   g456(.A(new_n809), .B(G290), .Z(new_n882));
  XNOR2_X1  g457(.A(new_n604), .B(G166), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n882), .B(new_n883), .Z(new_n884));
  XOR2_X1   g459(.A(new_n884), .B(KEYINPUT42), .Z(new_n885));
  XNOR2_X1  g460(.A(new_n881), .B(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n876), .B1(new_n886), .B2(G868), .ZN(G295));
  AOI21_X1  g462(.A(new_n876), .B1(new_n886), .B2(G868), .ZN(G331));
  NAND2_X1  g463(.A1(G301), .A2(G168), .ZN(new_n889));
  NAND2_X1  g464(.A1(G171), .A2(G286), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(new_n847), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n889), .A2(new_n845), .A3(new_n846), .A4(new_n890), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n894), .A2(new_n878), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT111), .ZN(new_n896));
  OR2_X1    g471(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n893), .A2(new_n896), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n897), .A2(new_n898), .A3(new_n892), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n895), .B1(new_n899), .B2(new_n879), .ZN(new_n900));
  INV_X1    g475(.A(new_n884), .ZN(new_n901));
  OR2_X1    g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(G37), .B1(new_n900), .B2(new_n901), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(KEYINPUT114), .B1(new_n904), .B2(KEYINPUT43), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n879), .A2(new_n894), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(KEYINPUT112), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT112), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n879), .A2(new_n894), .A3(new_n908), .ZN(new_n909));
  OAI211_X1 g484(.A(new_n907), .B(new_n909), .C1(new_n878), .C2(new_n899), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(new_n884), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n857), .B1(new_n900), .B2(new_n901), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(KEYINPUT43), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT114), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT43), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n902), .A2(new_n903), .A3(new_n915), .A4(new_n916), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n905), .A2(new_n914), .A3(KEYINPUT44), .A4(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT113), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n919), .B1(new_n913), .B2(KEYINPUT43), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n911), .A2(KEYINPUT113), .A3(new_n912), .A4(new_n916), .ZN(new_n921));
  AOI22_X1  g496(.A1(new_n920), .A2(new_n921), .B1(KEYINPUT43), .B2(new_n904), .ZN(new_n922));
  XOR2_X1   g497(.A(KEYINPUT110), .B(KEYINPUT44), .Z(new_n923));
  OAI21_X1  g498(.A(new_n918), .B1(new_n922), .B2(new_n923), .ZN(G397));
  AND4_X1   g499(.A1(G40), .A2(new_n486), .A3(new_n493), .A4(new_n496), .ZN(new_n925));
  INV_X1    g500(.A(G1384), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n517), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT45), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n925), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n929), .A2(G1996), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(new_n777), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n931), .B(KEYINPUT115), .ZN(new_n932));
  INV_X1    g507(.A(new_n929), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n716), .B(G2067), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n934), .B(KEYINPUT116), .ZN(new_n935));
  INV_X1    g510(.A(G1996), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n777), .A2(new_n936), .ZN(new_n937));
  OR2_X1    g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n932), .B1(new_n933), .B2(new_n938), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n791), .A2(new_n794), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n791), .A2(new_n794), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n933), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n939), .A2(new_n942), .ZN(new_n943));
  XNOR2_X1  g518(.A(G290), .B(G1986), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(new_n933), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT122), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n510), .A2(KEYINPUT4), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(KEYINPUT75), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n949), .A2(new_n512), .A3(new_n514), .ZN(new_n950));
  AOI21_X1  g525(.A(G1384), .B1(new_n950), .B2(new_n509), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n925), .B1(new_n951), .B2(KEYINPUT45), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n927), .A2(new_n928), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n803), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT117), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n486), .A2(new_n493), .A3(G40), .A4(new_n496), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n956), .B1(new_n927), .B2(new_n928), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n951), .A2(KEYINPUT45), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT117), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n959), .A2(new_n960), .A3(new_n803), .ZN(new_n961));
  XOR2_X1   g536(.A(KEYINPUT118), .B(KEYINPUT50), .Z(new_n962));
  AOI21_X1  g537(.A(new_n956), .B1(new_n951), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT119), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n964), .B1(new_n927), .B2(KEYINPUT50), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT50), .ZN(new_n966));
  AOI211_X1 g541(.A(KEYINPUT119), .B(new_n966), .C1(new_n517), .C2(new_n926), .ZN(new_n967));
  OAI211_X1 g542(.A(new_n745), .B(new_n963), .C1(new_n965), .C2(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n955), .A2(new_n961), .A3(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(G8), .ZN(new_n970));
  NOR2_X1   g545(.A1(G166), .A2(new_n970), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n971), .B(KEYINPUT55), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n807), .A2(G1976), .A3(new_n808), .ZN(new_n973));
  OAI211_X1 g548(.A(new_n973), .B(G8), .C1(new_n927), .C2(new_n956), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(KEYINPUT52), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n925), .A2(new_n951), .ZN(new_n976));
  INV_X1    g551(.A(G1976), .ZN(new_n977));
  AOI21_X1  g552(.A(KEYINPUT52), .B1(G288), .B2(new_n977), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n976), .A2(G8), .A3(new_n973), .A4(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(G1981), .B1(new_n597), .B2(new_n602), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n554), .A2(G86), .ZN(new_n981));
  INV_X1    g556(.A(G1981), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n981), .A2(new_n982), .A3(new_n601), .A4(new_n595), .ZN(new_n983));
  AND3_X1   g558(.A1(new_n980), .A2(KEYINPUT49), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(KEYINPUT49), .B1(new_n980), .B2(new_n983), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n986), .A2(new_n976), .A3(G8), .ZN(new_n987));
  AND3_X1   g562(.A1(new_n975), .A2(new_n979), .A3(new_n987), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n969), .A2(G8), .A3(new_n972), .A4(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n976), .A2(G8), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n987), .ZN(new_n992));
  NOR3_X1   g567(.A1(new_n992), .A2(G1976), .A3(G288), .ZN(new_n993));
  INV_X1    g568(.A(new_n983), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n991), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n989), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(KEYINPUT120), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT120), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n989), .A2(new_n998), .A3(new_n995), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT121), .ZN(new_n1000));
  INV_X1    g575(.A(new_n962), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n925), .B1(new_n927), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g577(.A(KEYINPUT119), .B1(new_n951), .B2(new_n966), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n927), .A2(new_n964), .A3(KEYINPUT50), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1002), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  AOI22_X1  g580(.A1(new_n1005), .A2(new_n745), .B1(new_n954), .B2(KEYINPUT117), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n970), .B1(new_n1006), .B2(new_n961), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n1000), .B(new_n988), .C1(new_n1007), .C2(new_n972), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n972), .B1(new_n969), .B2(G8), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n975), .A2(new_n979), .A3(new_n987), .ZN(new_n1010));
  OAI21_X1  g585(.A(KEYINPUT121), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(G1966), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n959), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n963), .B1(new_n965), .B2(new_n967), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1013), .B1(G2084), .B2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g590(.A1(G286), .A2(new_n970), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1015), .A2(KEYINPUT63), .A3(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1017), .B1(new_n1007), .B2(new_n972), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1008), .A2(new_n1011), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT63), .ZN(new_n1020));
  INV_X1    g595(.A(new_n972), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n925), .B1(new_n927), .B2(KEYINPUT50), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n951), .A2(new_n962), .ZN(new_n1023));
  NOR3_X1   g598(.A1(new_n1022), .A2(new_n1023), .A3(G2090), .ZN(new_n1024));
  AOI21_X1  g599(.A(G1971), .B1(new_n957), .B2(new_n958), .ZN(new_n1025));
  OAI21_X1  g600(.A(G8), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1010), .B1(new_n1021), .B2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n969), .A2(G8), .A3(new_n972), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1020), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  AOI221_X4 g606(.A(new_n947), .B1(new_n997), .B2(new_n999), .C1(new_n1019), .C2(new_n1031), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n957), .A2(KEYINPUT53), .A3(new_n445), .A4(new_n958), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1033), .B1(new_n1005), .B2(G1961), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT53), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1035), .B1(new_n959), .B2(G2078), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n623), .B1(new_n1034), .B2(new_n1037), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1029), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT51), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1040), .B1(new_n1015), .B2(G286), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1013), .B(G168), .C1(G2084), .C2(new_n1014), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(G8), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1040), .B1(new_n1042), .B2(G8), .ZN(new_n1045));
  OAI21_X1  g620(.A(KEYINPUT62), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1043), .A2(KEYINPUT51), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT62), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1047), .B(new_n1048), .C1(new_n1043), .C2(new_n1041), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1039), .A2(new_n1046), .A3(new_n1049), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n976), .A2(G2067), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1051), .B1(new_n1014), .B2(new_n707), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1052), .A2(new_n620), .ZN(new_n1053));
  AOI211_X1 g628(.A(new_n1051), .B(new_n628), .C1(new_n1014), .C2(new_n707), .ZN(new_n1054));
  OAI21_X1  g629(.A(KEYINPUT60), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(G1956), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1056), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1057));
  AND2_X1   g632(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1058));
  NOR2_X1   g633(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  XOR2_X1   g635(.A(KEYINPUT56), .B(G2072), .Z(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n957), .A2(new_n958), .A3(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1057), .A2(new_n1060), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT61), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1051), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n620), .A2(KEYINPUT60), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1066), .B(new_n1067), .C1(new_n1005), .C2(G1348), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT61), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1057), .A2(new_n1060), .A3(new_n1063), .A4(new_n1069), .ZN(new_n1070));
  AND3_X1   g645(.A1(new_n1065), .A2(new_n1068), .A3(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT124), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT59), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n957), .A2(new_n936), .A3(new_n958), .ZN(new_n1074));
  XOR2_X1   g649(.A(KEYINPUT58), .B(G1341), .Z(new_n1075));
  NAND2_X1  g650(.A1(new_n976), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(new_n564), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT125), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1072), .B(new_n1073), .C1(new_n1078), .C2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1077), .A2(KEYINPUT124), .A3(new_n564), .ZN(new_n1081));
  AOI211_X1 g656(.A(new_n1079), .B(new_n563), .C1(new_n1074), .C2(new_n1076), .ZN(new_n1082));
  OAI211_X1 g657(.A(KEYINPUT59), .B(new_n1081), .C1(new_n1082), .C2(KEYINPUT124), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1055), .A2(new_n1071), .A3(new_n1080), .A4(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1060), .B1(new_n1057), .B2(new_n1063), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT123), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1086), .B1(new_n1052), .B2(new_n620), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1066), .B1(new_n1005), .B2(G1348), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1088), .A2(KEYINPUT123), .A3(new_n628), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1085), .B1(new_n1090), .B2(new_n1064), .ZN(new_n1091));
  AND2_X1   g666(.A1(new_n1084), .A2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1047), .B1(new_n1043), .B2(new_n1041), .ZN(new_n1093));
  INV_X1    g668(.A(G1961), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1014), .A2(new_n1094), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1095), .A2(new_n1036), .A3(G301), .A4(new_n1033), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1038), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1029), .ZN(new_n1100));
  OAI21_X1  g675(.A(G171), .B1(new_n1034), .B2(new_n1037), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1101), .A2(KEYINPUT54), .A3(new_n1096), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1093), .A2(new_n1099), .A3(new_n1100), .A4(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1050), .B1(new_n1092), .B2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1032), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1019), .A2(new_n1031), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n997), .A2(new_n999), .ZN(new_n1107));
  AOI21_X1  g682(.A(KEYINPUT122), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n946), .B1(new_n1105), .B2(new_n1109), .ZN(new_n1110));
  NOR3_X1   g685(.A1(new_n929), .A2(G1986), .A3(G290), .ZN(new_n1111));
  XOR2_X1   g686(.A(new_n1111), .B(KEYINPUT48), .Z(new_n1112));
  NAND2_X1  g687(.A1(new_n943), .A2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n933), .B1(new_n935), .B2(new_n776), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n930), .A2(KEYINPUT46), .ZN(new_n1115));
  OR2_X1    g690(.A1(new_n930), .A2(KEYINPUT46), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1114), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g692(.A(new_n1117), .B(KEYINPUT47), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1113), .A2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n716), .A2(G2067), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1120), .B1(new_n939), .B2(new_n941), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1121), .A2(new_n929), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1119), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(KEYINPUT126), .B1(new_n1110), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT126), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1106), .A2(KEYINPUT122), .A3(new_n1107), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1084), .A2(new_n1091), .ZN(new_n1128));
  AND2_X1   g703(.A1(new_n1099), .A2(new_n1102), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1128), .A2(new_n1129), .A3(new_n1100), .A4(new_n1093), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1127), .A2(new_n1130), .A3(new_n1050), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1131), .A2(new_n1108), .ZN(new_n1132));
  OAI211_X1 g707(.A(new_n1126), .B(new_n1123), .C1(new_n1132), .C2(new_n946), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1125), .A2(new_n1133), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g709(.A(new_n665), .ZN(new_n1136));
  NOR4_X1   g710(.A1(G229), .A2(G227), .A3(new_n468), .A4(new_n1136), .ZN(new_n1137));
  NAND2_X1  g711(.A1(new_n874), .A2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g712(.A1(new_n922), .A2(new_n1138), .ZN(G308));
  OR2_X1    g713(.A1(new_n922), .A2(new_n1138), .ZN(G225));
endmodule


