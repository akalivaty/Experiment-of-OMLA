//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 1 1 0 0 0 1 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 1 0 1 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n808, new_n809, new_n810, new_n811, new_n813, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n903, new_n904, new_n905, new_n906,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n953, new_n954, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1008, new_n1009, new_n1010, new_n1011, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027;
  INV_X1    g000(.A(G227gat), .ZN(new_n202));
  INV_X1    g001(.A(G233gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NOR2_X1   g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT65), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT26), .ZN(new_n208));
  NAND2_X1  g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT26), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n205), .A2(new_n206), .A3(new_n210), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n208), .A2(new_n209), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213));
  INV_X1    g012(.A(G190gat), .ZN(new_n214));
  AND2_X1   g013(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT28), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT28), .ZN(new_n219));
  OAI211_X1 g018(.A(new_n219), .B(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n212), .A2(new_n213), .A3(new_n218), .A4(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT23), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI211_X1 g023(.A(KEYINPUT64), .B(KEYINPUT23), .C1(G169gat), .C2(G176gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n209), .B1(new_n213), .B2(KEYINPUT24), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  NOR2_X1   g027(.A1(G183gat), .A2(G190gat), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n230), .A2(KEYINPUT24), .A3(new_n213), .ZN(new_n231));
  AND4_X1   g030(.A1(KEYINPUT25), .A2(new_n226), .A3(new_n228), .A4(new_n231), .ZN(new_n232));
  AND2_X1   g031(.A1(G183gat), .A2(G190gat), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n233), .A2(new_n229), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n227), .B1(new_n234), .B2(KEYINPUT24), .ZN(new_n235));
  AOI21_X1  g034(.A(KEYINPUT25), .B1(new_n235), .B2(new_n226), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n221), .B1(new_n232), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT1), .ZN(new_n239));
  AND2_X1   g038(.A1(G127gat), .A2(G134gat), .ZN(new_n240));
  NOR2_X1   g039(.A1(G127gat), .A2(G134gat), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n239), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(G113gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(G120gat), .ZN(new_n244));
  AND2_X1   g043(.A1(KEYINPUT66), .A2(G120gat), .ZN(new_n245));
  NOR2_X1   g044(.A1(KEYINPUT66), .A2(G120gat), .ZN(new_n246));
  OAI21_X1  g045(.A(G113gat), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n242), .B1(new_n244), .B2(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(G127gat), .B(G134gat), .ZN(new_n249));
  INV_X1    g048(.A(G120gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(G113gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n244), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n249), .B1(new_n239), .B2(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n238), .B1(new_n248), .B2(new_n253), .ZN(new_n254));
  OR2_X1    g053(.A1(G127gat), .A2(G134gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(G127gat), .A2(G134gat), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT1), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT66), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(new_n250), .ZN(new_n259));
  NAND2_X1  g058(.A1(KEYINPUT66), .A2(G120gat), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n243), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n244), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n257), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G113gat), .B(G120gat), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n255), .B(new_n256), .C1(new_n264), .C2(KEYINPUT1), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n263), .A2(KEYINPUT67), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n254), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n237), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n226), .A2(new_n228), .A3(new_n231), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT25), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n235), .A2(KEYINPUT25), .A3(new_n226), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n273), .A2(new_n254), .A3(new_n266), .A4(new_n221), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n204), .B1(new_n268), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n268), .A2(new_n274), .A3(new_n204), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT34), .ZN(new_n277));
  AND3_X1   g076(.A1(new_n276), .A2(KEYINPUT32), .A3(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n277), .B1(new_n276), .B2(KEYINPUT32), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n275), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n276), .A2(KEYINPUT32), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT34), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n276), .A2(KEYINPUT32), .A3(new_n277), .ZN(new_n283));
  INV_X1    g082(.A(new_n275), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G15gat), .B(G43gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n286), .B(KEYINPUT68), .ZN(new_n287));
  XNOR2_X1  g086(.A(G71gat), .B(G99gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n287), .B(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT33), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n289), .B1(new_n276), .B2(new_n290), .ZN(new_n291));
  AND3_X1   g090(.A1(new_n280), .A2(new_n285), .A3(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n291), .B1(new_n280), .B2(new_n285), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT36), .ZN(new_n294));
  NOR3_X1   g093(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n291), .ZN(new_n296));
  NOR3_X1   g095(.A1(new_n278), .A2(new_n279), .A3(new_n275), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n284), .B1(new_n282), .B2(new_n283), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n296), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n280), .A2(new_n285), .A3(new_n291), .ZN(new_n300));
  AOI21_X1  g099(.A(KEYINPUT36), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n295), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(G78gat), .B(G106gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n303), .B(G50gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(KEYINPUT77), .B(KEYINPUT31), .ZN(new_n305));
  INV_X1    g104(.A(G22gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n305), .B(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n304), .B(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT78), .ZN(new_n310));
  XNOR2_X1  g109(.A(G141gat), .B(G148gat), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT2), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n312), .B1(G155gat), .B2(G162gat), .ZN(new_n313));
  OAI21_X1  g112(.A(KEYINPUT73), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G155gat), .B(G162gat), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(G155gat), .A2(G162gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(KEYINPUT2), .ZN(new_n319));
  INV_X1    g118(.A(G141gat), .ZN(new_n320));
  INV_X1    g119(.A(G148gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(G141gat), .A2(G148gat), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n319), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n324), .A2(KEYINPUT73), .A3(new_n315), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n317), .A2(KEYINPUT3), .A3(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT69), .ZN(new_n327));
  AND2_X1   g126(.A1(G197gat), .A2(G204gat), .ZN(new_n328));
  NOR2_X1   g127(.A1(G197gat), .A2(G204gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n327), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n331), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n333), .B(KEYINPUT69), .C1(new_n329), .C2(new_n328), .ZN(new_n334));
  XOR2_X1   g133(.A(G211gat), .B(G218gat), .Z(new_n335));
  NAND3_X1  g134(.A1(new_n332), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(G211gat), .B(G218gat), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n337), .B(new_n333), .C1(new_n329), .C2(new_n328), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(KEYINPUT70), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  NAND4_X1  g139(.A1(new_n332), .A2(new_n334), .A3(KEYINPUT70), .A4(new_n335), .ZN(new_n341));
  AND2_X1   g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT29), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n317), .A2(new_n343), .A3(new_n325), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n310), .B(new_n326), .C1(new_n342), .C2(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n344), .B1(new_n340), .B2(new_n341), .ZN(new_n346));
  INV_X1    g145(.A(new_n326), .ZN(new_n347));
  OAI21_X1  g146(.A(KEYINPUT78), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(KEYINPUT75), .B(KEYINPUT3), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  AND3_X1   g149(.A1(new_n324), .A2(KEYINPUT73), .A3(new_n315), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n315), .B1(new_n324), .B2(KEYINPUT73), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n350), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(new_n343), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n342), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n345), .A2(new_n348), .A3(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(G228gat), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n357), .A2(new_n203), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n335), .B1(new_n331), .B2(new_n330), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(new_n338), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n349), .B1(new_n361), .B2(new_n343), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n317), .A2(new_n325), .ZN(new_n363));
  OAI22_X1  g162(.A1(new_n362), .A2(new_n363), .B1(new_n357), .B2(new_n203), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n364), .B1(new_n354), .B2(new_n342), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n309), .B1(new_n359), .B2(new_n366), .ZN(new_n367));
  AOI211_X1 g166(.A(new_n365), .B(new_n308), .C1(new_n356), .C2(new_n358), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(G8gat), .B(G36gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(G64gat), .B(G92gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n370), .B(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n340), .A2(new_n341), .ZN(new_n373));
  NAND2_X1  g172(.A1(G226gat), .A2(G233gat), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n375), .B1(new_n237), .B2(new_n343), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n374), .B(KEYINPUT71), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n377), .B1(new_n273), .B2(new_n221), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n373), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT72), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n237), .A2(new_n375), .ZN(new_n381));
  AOI21_X1  g180(.A(KEYINPUT29), .B1(new_n273), .B2(new_n221), .ZN(new_n382));
  INV_X1    g181(.A(new_n377), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n381), .B(new_n342), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  AND3_X1   g183(.A1(new_n379), .A2(new_n380), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n380), .B1(new_n379), .B2(new_n384), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n372), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n379), .A2(new_n384), .ZN(new_n388));
  INV_X1    g187(.A(new_n372), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n387), .A2(KEYINPUT30), .A3(new_n390), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n390), .A2(KEYINPUT30), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(G225gat), .A2(G233gat), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n248), .A2(new_n253), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n363), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT4), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n396), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n267), .A2(KEYINPUT4), .A3(new_n363), .ZN(new_n401));
  NOR3_X1   g200(.A1(new_n248), .A2(new_n253), .A3(KEYINPUT74), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT74), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n403), .B1(new_n263), .B2(new_n265), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n353), .B(new_n326), .C1(new_n402), .C2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n400), .A2(new_n401), .A3(new_n405), .ZN(new_n406));
  OAI21_X1  g205(.A(KEYINPUT74), .B1(new_n248), .B2(new_n253), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n263), .A2(new_n403), .A3(new_n265), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n363), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n398), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n396), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n406), .A2(KEYINPUT5), .A3(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n267), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n351), .A2(new_n352), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n399), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n396), .A2(KEYINPUT5), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n363), .A2(new_n397), .A3(KEYINPUT4), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n415), .A2(new_n405), .A3(new_n416), .A4(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n412), .A2(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(G1gat), .B(G29gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n420), .B(G85gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(KEYINPUT0), .B(G57gat), .ZN(new_n422));
  XOR2_X1   g221(.A(new_n421), .B(new_n422), .Z(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n419), .A2(new_n424), .ZN(new_n425));
  XOR2_X1   g224(.A(KEYINPUT76), .B(KEYINPUT6), .Z(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n412), .A2(new_n418), .A3(new_n423), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n425), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n423), .B1(new_n412), .B2(new_n418), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(new_n426), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n369), .B1(new_n394), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g232(.A(KEYINPUT79), .B1(new_n302), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n369), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT30), .ZN(new_n436));
  NOR4_X1   g235(.A1(KEYINPUT65), .A2(KEYINPUT26), .A3(G169gat), .A4(G176gat), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n210), .B1(new_n205), .B2(new_n206), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n233), .B1(new_n439), .B2(new_n209), .ZN(new_n440));
  AND2_X1   g239(.A1(new_n218), .A2(new_n220), .ZN(new_n441));
  AOI22_X1  g240(.A1(new_n271), .A2(new_n272), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n374), .B1(new_n442), .B2(KEYINPUT29), .ZN(new_n443));
  INV_X1    g242(.A(new_n378), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n342), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n383), .B1(new_n237), .B2(new_n343), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n374), .B1(new_n273), .B2(new_n221), .ZN(new_n447));
  NOR3_X1   g246(.A1(new_n446), .A2(new_n373), .A3(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(KEYINPUT72), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n379), .A2(new_n380), .A3(new_n384), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n436), .B1(new_n451), .B2(new_n372), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n392), .B1(new_n452), .B2(new_n390), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n414), .B1(new_n254), .B2(new_n266), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n405), .B(new_n417), .C1(new_n454), .C2(KEYINPUT4), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(new_n396), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n414), .B1(new_n402), .B2(new_n404), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT80), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n457), .A2(new_n458), .A3(new_n395), .A4(new_n398), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n457), .A2(new_n395), .A3(new_n398), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT80), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n456), .A2(KEYINPUT39), .A3(new_n459), .A4(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT39), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n455), .A2(new_n463), .A3(new_n396), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n462), .A2(new_n423), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(KEYINPUT40), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT40), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n462), .A2(new_n467), .A3(new_n423), .A4(new_n464), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT81), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n425), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n430), .A2(KEYINPUT81), .ZN(new_n471));
  AOI22_X1  g270(.A1(new_n466), .A2(new_n468), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n435), .B1(new_n453), .B2(new_n472), .ZN(new_n473));
  AND2_X1   g272(.A1(new_n428), .A2(new_n427), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n430), .A2(KEYINPUT81), .ZN(new_n475));
  AOI211_X1 g274(.A(new_n469), .B(new_n423), .C1(new_n412), .C2(new_n418), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT82), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT82), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n474), .B(new_n479), .C1(new_n475), .C2(new_n476), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n478), .A2(new_n431), .A3(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n342), .B1(new_n376), .B2(new_n378), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT83), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n381), .B(new_n373), .C1(new_n382), .C2(new_n383), .ZN(new_n485));
  OAI211_X1 g284(.A(KEYINPUT83), .B(new_n342), .C1(new_n376), .C2(new_n378), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT37), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT84), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT38), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT37), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n389), .B1(new_n388), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n487), .A2(KEYINPUT84), .A3(KEYINPUT37), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n490), .A2(new_n491), .A3(new_n493), .A4(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(KEYINPUT37), .B1(new_n385), .B2(new_n386), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(new_n493), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT38), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n495), .A2(new_n390), .A3(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n473), .B1(new_n481), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n294), .B1(new_n292), .B2(new_n293), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n299), .A2(KEYINPUT36), .A3(new_n300), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT79), .ZN(new_n504));
  AOI22_X1  g303(.A1(new_n391), .A2(new_n393), .B1(new_n429), .B2(new_n431), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n503), .B(new_n504), .C1(new_n369), .C2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n434), .A2(new_n500), .A3(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n299), .A2(new_n369), .A3(new_n300), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT85), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT85), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n299), .A2(new_n369), .A3(new_n510), .A4(new_n300), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n509), .A2(new_n511), .A3(new_n505), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(KEYINPUT35), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT35), .ZN(new_n514));
  INV_X1    g313(.A(new_n508), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n481), .A2(new_n514), .A3(new_n515), .A4(new_n394), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  AND3_X1   g316(.A1(new_n507), .A2(new_n517), .A3(KEYINPUT86), .ZN(new_n518));
  AOI21_X1  g317(.A(KEYINPUT86), .B1(new_n507), .B2(new_n517), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(G15gat), .B(G22gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(KEYINPUT92), .ZN(new_n522));
  INV_X1    g321(.A(G1gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n521), .A2(KEYINPUT92), .A3(G1gat), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT16), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n521), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n524), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(G8gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(G50gat), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n531), .A2(G43gat), .ZN(new_n532));
  INV_X1    g331(.A(G43gat), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n533), .A2(G50gat), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT15), .ZN(new_n535));
  NOR3_X1   g334(.A1(new_n532), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NOR2_X1   g335(.A1(G29gat), .A2(G36gat), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT14), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g338(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(G36gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(KEYINPUT88), .B(G29gat), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n536), .B1(new_n544), .B2(KEYINPUT89), .ZN(new_n545));
  XOR2_X1   g344(.A(KEYINPUT88), .B(G29gat), .Z(new_n546));
  AOI22_X1  g345(.A1(new_n546), .A2(G36gat), .B1(new_n540), .B2(new_n539), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT89), .ZN(new_n548));
  OR3_X1    g347(.A1(new_n532), .A2(new_n534), .A3(new_n535), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT90), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n551), .B1(new_n531), .B2(G43gat), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n533), .A2(KEYINPUT90), .A3(G50gat), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n552), .B(new_n553), .C1(new_n533), .C2(G50gat), .ZN(new_n554));
  AND2_X1   g353(.A1(new_n554), .A2(new_n535), .ZN(new_n555));
  AOI22_X1  g354(.A1(new_n545), .A2(new_n550), .B1(new_n547), .B2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT91), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n556), .A2(new_n557), .A3(KEYINPUT17), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(KEYINPUT17), .B1(new_n556), .B2(new_n557), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n530), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(G229gat), .A2(G233gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n528), .B(G8gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(new_n556), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n561), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT18), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n564), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT17), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n545), .A2(new_n550), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n547), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n569), .B1(new_n572), .B2(KEYINPUT91), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(new_n558), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n568), .B1(new_n574), .B2(new_n530), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n575), .A2(KEYINPUT18), .A3(new_n562), .ZN(new_n576));
  AOI21_X1  g375(.A(KEYINPUT93), .B1(new_n530), .B2(new_n572), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n577), .B1(new_n530), .B2(new_n572), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n562), .B(KEYINPUT13), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n563), .A2(KEYINPUT93), .A3(new_n556), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n578), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n567), .A2(new_n576), .A3(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(G113gat), .B(G141gat), .ZN(new_n584));
  INV_X1    g383(.A(G197gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(KEYINPUT11), .B(G169gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XOR2_X1   g387(.A(new_n588), .B(KEYINPUT87), .Z(new_n589));
  INV_X1    g388(.A(KEYINPUT12), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n583), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n567), .A2(new_n591), .A3(new_n576), .A4(new_n582), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT94), .ZN(new_n596));
  XOR2_X1   g395(.A(G57gat), .B(G64gat), .Z(new_n597));
  INV_X1    g396(.A(KEYINPUT9), .ZN(new_n598));
  INV_X1    g397(.A(G71gat), .ZN(new_n599));
  INV_X1    g398(.A(G78gat), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G71gat), .B(G78gat), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n597), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n602), .B1(new_n597), .B2(new_n601), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n596), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n597), .A2(new_n601), .ZN(new_n607));
  INV_X1    g406(.A(new_n602), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n609), .A2(KEYINPUT94), .A3(new_n603), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n563), .B1(new_n611), .B2(KEYINPUT21), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(KEYINPUT95), .ZN(new_n613));
  INV_X1    g412(.A(G127gat), .ZN(new_n614));
  INV_X1    g413(.A(new_n610), .ZN(new_n615));
  AOI21_X1  g414(.A(KEYINPUT94), .B1(new_n609), .B2(new_n603), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT21), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n530), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT95), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n613), .A2(new_n614), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n614), .B1(new_n613), .B2(new_n621), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n617), .A2(new_n618), .ZN(new_n625));
  XOR2_X1   g424(.A(G183gat), .B(G211gat), .Z(new_n626));
  OR2_X1    g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n625), .A2(new_n626), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(G231gat), .A2(G233gat), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n627), .A2(new_n628), .A3(G231gat), .A4(G233gat), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n624), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(G155gat), .ZN(new_n636));
  OAI211_X1 g435(.A(new_n631), .B(new_n632), .C1(new_n622), .C2(new_n623), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n634), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n636), .B1(new_n634), .B2(new_n637), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(G190gat), .B(G218gat), .ZN(new_n642));
  AOI21_X1  g441(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n642), .B(new_n643), .Z(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(G85gat), .A2(G92gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(KEYINPUT7), .ZN(new_n647));
  OR2_X1    g446(.A1(G85gat), .A2(G92gat), .ZN(new_n648));
  INV_X1    g447(.A(G99gat), .ZN(new_n649));
  INV_X1    g448(.A(G106gat), .ZN(new_n650));
  OAI21_X1  g449(.A(KEYINPUT8), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n647), .A2(new_n648), .A3(new_n651), .ZN(new_n652));
  XOR2_X1   g451(.A(G99gat), .B(G106gat), .Z(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n653), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n655), .A2(new_n648), .A3(new_n647), .A4(new_n651), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n574), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n556), .A2(new_n656), .A3(new_n654), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g460(.A(G134gat), .B(G162gat), .Z(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT96), .ZN(new_n663));
  AND2_X1   g462(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n661), .A2(new_n663), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n645), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n661), .A2(new_n663), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n661), .A2(new_n663), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n667), .A2(new_n644), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n520), .A2(new_n595), .A3(new_n641), .A4(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT98), .ZN(new_n672));
  XNOR2_X1  g471(.A(KEYINPUT97), .B(KEYINPUT10), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n611), .A2(new_n657), .ZN(new_n674));
  OAI211_X1 g473(.A(new_n654), .B(new_n656), .C1(new_n605), .C2(new_n604), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n673), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n611), .A2(KEYINPUT10), .A3(new_n656), .A4(new_n654), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n672), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n673), .ZN(new_n680));
  AOI22_X1  g479(.A1(new_n606), .A2(new_n610), .B1(new_n656), .B2(new_n654), .ZN(new_n681));
  INV_X1    g480(.A(new_n675), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n680), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n683), .A2(KEYINPUT98), .A3(new_n677), .ZN(new_n684));
  NAND2_X1  g483(.A1(G230gat), .A2(G233gat), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n679), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(G120gat), .B(G148gat), .ZN(new_n687));
  XNOR2_X1  g486(.A(G176gat), .B(G204gat), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n685), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n674), .A2(new_n691), .A3(new_n675), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n686), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n685), .B1(new_n676), .B2(new_n678), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(new_n692), .ZN(new_n695));
  AOI21_X1  g494(.A(KEYINPUT99), .B1(new_n695), .B2(new_n689), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT99), .ZN(new_n697));
  AOI211_X1 g496(.A(new_n697), .B(new_n690), .C1(new_n694), .C2(new_n692), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n693), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n671), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n432), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(G1gat), .ZN(G1324gat));
  NOR3_X1   g502(.A1(new_n671), .A2(new_n699), .A3(new_n394), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n526), .A2(new_n529), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n526), .A2(new_n529), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n704), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT42), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n704), .A2(KEYINPUT42), .A3(new_n706), .A4(new_n707), .ZN(new_n711));
  OAI211_X1 g510(.A(new_n710), .B(new_n711), .C1(new_n529), .C2(new_n704), .ZN(G1325gat));
  NOR2_X1   g511(.A1(new_n292), .A2(new_n293), .ZN(new_n713));
  AOI21_X1  g512(.A(G15gat), .B1(new_n700), .B2(new_n713), .ZN(new_n714));
  AND2_X1   g513(.A1(new_n302), .A2(G15gat), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n714), .B1(new_n700), .B2(new_n715), .ZN(G1326gat));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n435), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(G22gat), .ZN(new_n718));
  XNOR2_X1  g517(.A(KEYINPUT100), .B(KEYINPUT43), .ZN(new_n719));
  NOR4_X1   g518(.A1(new_n671), .A2(G22gat), .A3(new_n699), .A4(new_n369), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n718), .A2(new_n719), .A3(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n719), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n306), .B1(new_n700), .B2(new_n435), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n723), .B1(new_n724), .B2(new_n720), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n722), .A2(new_n725), .ZN(G1327gat));
  NAND2_X1  g525(.A1(new_n507), .A2(new_n517), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT86), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n507), .A2(new_n517), .A3(KEYINPUT86), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n641), .A2(new_n699), .A3(new_n670), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n729), .A2(new_n730), .A3(new_n595), .A4(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n733), .A2(new_n701), .A3(new_n543), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT45), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT44), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n670), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n729), .A2(new_n730), .A3(new_n737), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n302), .A2(new_n433), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n500), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n517), .A2(new_n740), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n666), .A2(new_n669), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n736), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT101), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n745), .B1(new_n639), .B2(new_n640), .ZN(new_n746));
  INV_X1    g545(.A(new_n640), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n747), .A2(KEYINPUT101), .A3(new_n638), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n750), .A2(new_n699), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n738), .A2(new_n744), .A3(new_n595), .A4(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n546), .B1(new_n752), .B2(new_n432), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n735), .A2(new_n753), .ZN(G1328gat));
  INV_X1    g553(.A(KEYINPUT104), .ZN(new_n755));
  OAI21_X1  g554(.A(G36gat), .B1(new_n752), .B2(new_n394), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n394), .A2(G36gat), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n732), .A2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT46), .ZN(new_n760));
  AOI21_X1  g559(.A(KEYINPUT103), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT103), .ZN(new_n762));
  NOR4_X1   g561(.A1(new_n732), .A2(new_n762), .A3(KEYINPUT46), .A4(new_n758), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n756), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT102), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n520), .A2(new_n595), .A3(new_n731), .A4(new_n757), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n765), .B1(new_n766), .B2(KEYINPUT46), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n765), .B(KEYINPUT46), .C1(new_n732), .C2(new_n758), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n755), .B1(new_n764), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(KEYINPUT102), .B1(new_n759), .B2(new_n760), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n768), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n762), .B1(new_n766), .B2(KEYINPUT46), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n759), .A2(KEYINPUT103), .A3(new_n760), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n773), .A2(new_n776), .A3(KEYINPUT104), .A4(new_n756), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n771), .A2(new_n777), .ZN(G1329gat));
  OAI21_X1  g577(.A(G43gat), .B1(new_n752), .B2(new_n503), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT47), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(KEYINPUT105), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n733), .A2(new_n533), .A3(new_n713), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n779), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  OR2_X1    g582(.A1(new_n780), .A2(KEYINPUT105), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n783), .B(new_n784), .ZN(G1330gat));
  OAI21_X1  g584(.A(G50gat), .B1(new_n752), .B2(new_n369), .ZN(new_n786));
  AOI21_X1  g585(.A(KEYINPUT48), .B1(new_n786), .B2(KEYINPUT107), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n369), .A2(G50gat), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(KEYINPUT106), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n733), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n786), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n786), .B(new_n790), .C1(KEYINPUT107), .C2(KEYINPUT48), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(G1331gat));
  NAND3_X1  g593(.A1(new_n747), .A2(new_n670), .A3(new_n638), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n795), .A2(new_n595), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n699), .ZN(new_n797));
  XOR2_X1   g596(.A(new_n797), .B(KEYINPUT108), .Z(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n741), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(new_n701), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n801), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g601(.A1(new_n799), .A2(new_n394), .ZN(new_n803));
  NOR2_X1   g602(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n804));
  AND2_X1   g603(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n803), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n806), .B1(new_n803), .B2(new_n804), .ZN(G1333gat));
  NAND3_X1  g606(.A1(new_n800), .A2(new_n599), .A3(new_n713), .ZN(new_n808));
  OAI21_X1  g607(.A(G71gat), .B1(new_n799), .B2(new_n503), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT50), .ZN(new_n811));
  XNOR2_X1  g610(.A(new_n810), .B(new_n811), .ZN(G1334gat));
  NOR2_X1   g611(.A1(new_n799), .A2(new_n369), .ZN(new_n813));
  XNOR2_X1  g612(.A(new_n813), .B(new_n600), .ZN(G1335gat));
  NOR2_X1   g613(.A1(new_n641), .A2(new_n595), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n738), .A2(new_n744), .A3(new_n699), .A4(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(G85gat), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n816), .A2(new_n817), .A3(new_n432), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n741), .A2(new_n742), .A3(new_n815), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT51), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(KEYINPUT110), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT110), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n819), .A2(new_n823), .A3(new_n820), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n741), .A2(KEYINPUT51), .A3(new_n742), .A4(new_n815), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n826), .B(KEYINPUT109), .ZN(new_n827));
  OAI211_X1 g626(.A(new_n701), .B(new_n699), .C1(new_n825), .C2(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n818), .B1(new_n828), .B2(new_n817), .ZN(G1336gat));
  NOR2_X1   g628(.A1(new_n394), .A2(G92gat), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n699), .B(new_n830), .C1(new_n825), .C2(new_n827), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT52), .ZN(new_n832));
  OAI21_X1  g631(.A(G92gat), .B1(new_n816), .B2(new_n394), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n831), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n821), .A2(new_n826), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n835), .A2(new_n699), .A3(new_n830), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n834), .B1(new_n837), .B2(new_n832), .ZN(G1337gat));
  NOR3_X1   g637(.A1(new_n292), .A2(new_n293), .A3(G99gat), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n699), .B(new_n839), .C1(new_n825), .C2(new_n827), .ZN(new_n840));
  OAI21_X1  g639(.A(G99gat), .B1(new_n816), .B2(new_n503), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT111), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n840), .A2(KEYINPUT111), .A3(new_n841), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(G1338gat));
  NAND3_X1  g645(.A1(new_n699), .A2(new_n435), .A3(new_n650), .ZN(new_n847));
  XOR2_X1   g646(.A(new_n847), .B(KEYINPUT112), .Z(new_n848));
  OAI21_X1  g647(.A(new_n848), .B1(new_n825), .B2(new_n827), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT53), .ZN(new_n850));
  OAI21_X1  g649(.A(G106gat), .B1(new_n816), .B2(new_n369), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n835), .A2(new_n848), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n852), .B1(new_n854), .B2(new_n850), .ZN(G1339gat));
  INV_X1    g654(.A(new_n693), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT54), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n676), .A2(new_n678), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n857), .B1(new_n858), .B2(new_n691), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n686), .A2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(new_n694), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n690), .B1(new_n861), .B2(new_n857), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(KEYINPUT55), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT55), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n860), .A2(new_n862), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n856), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  AND3_X1   g666(.A1(new_n567), .A2(new_n582), .A3(new_n576), .ZN(new_n868));
  OAI21_X1  g667(.A(KEYINPUT113), .B1(new_n575), .B2(new_n562), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n561), .A2(new_n564), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT113), .ZN(new_n871));
  INV_X1    g670(.A(new_n562), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n578), .A2(new_n581), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(new_n579), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n869), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  AOI22_X1  g675(.A1(new_n868), .A2(new_n591), .B1(new_n876), .B2(new_n588), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n742), .A2(new_n867), .A3(new_n877), .ZN(new_n878));
  AOI22_X1  g677(.A1(new_n867), .A2(new_n595), .B1(new_n877), .B2(new_n699), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n878), .B1(new_n879), .B2(new_n742), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(new_n749), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n795), .A2(new_n699), .A3(new_n595), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n453), .A2(new_n432), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n884), .A2(new_n515), .A3(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(new_n595), .ZN(new_n887));
  OAI21_X1  g686(.A(G113gat), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n509), .A2(new_n511), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n884), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n885), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n595), .A2(new_n243), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n888), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n893), .B(KEYINPUT114), .ZN(G1340gat));
  INV_X1    g693(.A(new_n699), .ZN(new_n895));
  OAI21_X1  g694(.A(G120gat), .B1(new_n886), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n699), .B1(new_n246), .B2(new_n245), .ZN(new_n897));
  XOR2_X1   g696(.A(new_n897), .B(KEYINPUT115), .Z(new_n898));
  OAI21_X1  g697(.A(new_n896), .B1(new_n891), .B2(new_n898), .ZN(G1341gat));
  NOR3_X1   g698(.A1(new_n886), .A2(new_n614), .A3(new_n749), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n890), .A2(new_n641), .A3(new_n885), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n900), .B1(new_n901), .B2(new_n614), .ZN(G1342gat));
  NOR3_X1   g701(.A1(new_n891), .A2(G134gat), .A3(new_n670), .ZN(new_n903));
  XNOR2_X1  g702(.A(KEYINPUT116), .B(KEYINPUT56), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n903), .B(new_n904), .ZN(new_n905));
  OAI21_X1  g704(.A(G134gat), .B1(new_n886), .B2(new_n670), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(G1343gat));
  AND3_X1   g706(.A1(new_n742), .A2(new_n867), .A3(new_n877), .ZN(new_n908));
  AOI21_X1  g707(.A(KEYINPUT55), .B1(new_n863), .B2(KEYINPUT118), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT118), .ZN(new_n910));
  AOI211_X1 g709(.A(new_n910), .B(new_n865), .C1(new_n860), .C2(new_n862), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n595), .B(new_n693), .C1(new_n909), .C2(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT117), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n877), .A2(new_n913), .A3(new_n699), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n876), .A2(new_n588), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n915), .A2(new_n699), .A3(new_n594), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(KEYINPUT117), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n912), .A2(new_n914), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n908), .B1(new_n918), .B2(new_n670), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n883), .B1(new_n919), .B2(new_n641), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(new_n435), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(KEYINPUT57), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n882), .B1(new_n880), .B2(new_n749), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n923), .A2(KEYINPUT57), .A3(new_n369), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n885), .A2(new_n503), .ZN(new_n926));
  INV_X1    g725(.A(new_n926), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n922), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(G141gat), .B1(new_n928), .B2(new_n887), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n923), .A2(new_n369), .A3(new_n926), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n930), .A2(new_n320), .A3(new_n595), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(KEYINPUT58), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT58), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n929), .A2(new_n934), .A3(new_n931), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n933), .A2(new_n935), .ZN(G1344gat));
  NAND3_X1  g735(.A1(new_n930), .A2(new_n321), .A3(new_n699), .ZN(new_n937));
  XOR2_X1   g736(.A(new_n937), .B(KEYINPUT119), .Z(new_n938));
  INV_X1    g737(.A(new_n928), .ZN(new_n939));
  AOI211_X1 g738(.A(KEYINPUT59), .B(new_n321), .C1(new_n939), .C2(new_n699), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT59), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT57), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n920), .A2(new_n942), .A3(new_n435), .ZN(new_n943));
  OAI21_X1  g742(.A(KEYINPUT57), .B1(new_n923), .B2(new_n369), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n945), .A2(new_n895), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(new_n927), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n941), .B1(new_n947), .B2(G148gat), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n938), .B1(new_n940), .B2(new_n948), .ZN(G1345gat));
  AOI21_X1  g748(.A(G155gat), .B1(new_n930), .B2(new_n641), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n750), .A2(G155gat), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n950), .B1(new_n939), .B2(new_n951), .ZN(G1346gat));
  AOI21_X1  g751(.A(G162gat), .B1(new_n930), .B2(new_n742), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n742), .A2(G162gat), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n953), .B1(new_n939), .B2(new_n954), .ZN(G1347gat));
  NOR2_X1   g754(.A1(new_n701), .A2(new_n394), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n884), .A2(new_n515), .A3(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT122), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND4_X1  g758(.A1(new_n884), .A2(KEYINPUT122), .A3(new_n515), .A4(new_n956), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n959), .A2(new_n595), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(G169gat), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT123), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n961), .A2(KEYINPUT123), .A3(G169gat), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n884), .A2(new_n889), .A3(new_n956), .ZN(new_n966));
  OR2_X1    g765(.A1(new_n966), .A2(KEYINPUT120), .ZN(new_n967));
  INV_X1    g766(.A(G169gat), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n966), .A2(KEYINPUT120), .ZN(new_n969));
  NAND4_X1  g768(.A1(new_n967), .A2(new_n968), .A3(new_n595), .A4(new_n969), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT121), .ZN(new_n971));
  AND2_X1   g770(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n970), .A2(new_n971), .ZN(new_n973));
  OAI211_X1 g772(.A(new_n964), .B(new_n965), .C1(new_n972), .C2(new_n973), .ZN(G1348gat));
  AND2_X1   g773(.A1(new_n959), .A2(new_n960), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n975), .A2(G176gat), .A3(new_n699), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT124), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n967), .A2(new_n699), .A3(new_n969), .ZN(new_n979));
  INV_X1    g778(.A(G176gat), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND4_X1  g780(.A1(new_n975), .A2(KEYINPUT124), .A3(G176gat), .A4(new_n699), .ZN(new_n982));
  AND3_X1   g781(.A1(new_n978), .A2(new_n981), .A3(new_n982), .ZN(G1349gat));
  NAND3_X1  g782(.A1(new_n959), .A2(new_n750), .A3(new_n960), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n984), .A2(G183gat), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n641), .B1(new_n216), .B2(new_n215), .ZN(new_n986));
  OR2_X1    g785(.A1(new_n966), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  XNOR2_X1  g787(.A(new_n988), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g788(.A1(new_n959), .A2(new_n742), .A3(new_n960), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n990), .A2(G190gat), .ZN(new_n991));
  INV_X1    g790(.A(KEYINPUT61), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n990), .A2(KEYINPUT61), .A3(G190gat), .ZN(new_n994));
  NAND4_X1  g793(.A1(new_n967), .A2(new_n214), .A3(new_n742), .A4(new_n969), .ZN(new_n995));
  INV_X1    g794(.A(KEYINPUT125), .ZN(new_n996));
  AND2_X1   g795(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NOR2_X1   g796(.A1(new_n995), .A2(new_n996), .ZN(new_n998));
  OAI211_X1 g797(.A(new_n993), .B(new_n994), .C1(new_n997), .C2(new_n998), .ZN(G1351gat));
  NAND2_X1  g798(.A1(new_n956), .A2(new_n503), .ZN(new_n1000));
  NOR2_X1   g799(.A1(new_n945), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g800(.A(new_n585), .B1(new_n1001), .B2(new_n595), .ZN(new_n1002));
  NOR2_X1   g801(.A1(new_n923), .A2(new_n369), .ZN(new_n1003));
  INV_X1    g802(.A(new_n1000), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NOR3_X1   g804(.A1(new_n1005), .A2(G197gat), .A3(new_n887), .ZN(new_n1006));
  OR2_X1    g805(.A1(new_n1002), .A2(new_n1006), .ZN(G1352gat));
  NOR3_X1   g806(.A1(new_n1005), .A2(G204gat), .A3(new_n895), .ZN(new_n1008));
  XNOR2_X1  g807(.A(new_n1008), .B(KEYINPUT62), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n946), .A2(new_n1004), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n1010), .A2(G204gat), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n1009), .A2(new_n1011), .ZN(G1353gat));
  INV_X1    g811(.A(G211gat), .ZN(new_n1013));
  NAND4_X1  g812(.A1(new_n1003), .A2(new_n1013), .A3(new_n641), .A4(new_n1004), .ZN(new_n1014));
  NAND4_X1  g813(.A1(new_n943), .A2(new_n641), .A3(new_n944), .A4(new_n1004), .ZN(new_n1015));
  AND3_X1   g814(.A1(new_n1015), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1016));
  AOI21_X1  g815(.A(KEYINPUT63), .B1(new_n1015), .B2(G211gat), .ZN(new_n1017));
  OAI21_X1  g816(.A(new_n1014), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g817(.A(KEYINPUT126), .ZN(new_n1019));
  NAND2_X1  g818(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  OAI211_X1 g819(.A(KEYINPUT126), .B(new_n1014), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1021));
  NAND2_X1  g820(.A1(new_n1020), .A2(new_n1021), .ZN(G1354gat));
  INV_X1    g821(.A(G218gat), .ZN(new_n1023));
  OAI21_X1  g822(.A(new_n1023), .B1(new_n1005), .B2(new_n670), .ZN(new_n1024));
  NOR2_X1   g823(.A1(new_n1024), .A2(KEYINPUT127), .ZN(new_n1025));
  AND2_X1   g824(.A1(new_n1024), .A2(KEYINPUT127), .ZN(new_n1026));
  NOR2_X1   g825(.A1(new_n670), .A2(new_n1023), .ZN(new_n1027));
  AOI211_X1 g826(.A(new_n1025), .B(new_n1026), .C1(new_n1001), .C2(new_n1027), .ZN(G1355gat));
endmodule


