//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 0 0 1 1 0 1 0 0 1 1 0 1 0 1 0 0 1 1 0 0 0 0 1 0 1 0 0 1 0 0 1 1 1 0 1 0 1 1 0 0 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:13 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n553, new_n555, new_n556, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n626, new_n627, new_n630, new_n632, new_n633,
    new_n634, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1225, new_n1226,
    new_n1227;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT65), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT66), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n454), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI211_X1 g039(.A(G137), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  AOI21_X1  g043(.A(KEYINPUT68), .B1(new_n465), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n465), .A2(KEYINPUT68), .A3(new_n468), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n463), .A2(new_n464), .ZN(new_n472));
  INV_X1    g047(.A(G125), .ZN(new_n473));
  INV_X1    g048(.A(G113), .ZN(new_n474));
  OAI22_X1  g049(.A1(new_n472), .A2(new_n473), .B1(new_n474), .B2(new_n466), .ZN(new_n475));
  AOI22_X1  g050(.A1(new_n470), .A2(new_n471), .B1(G2105), .B2(new_n475), .ZN(new_n476));
  XOR2_X1   g051(.A(new_n476), .B(KEYINPUT69), .Z(G160));
  OR2_X1    g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT70), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(G112), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n485), .B1(new_n486), .B2(G2105), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n472), .A2(G2105), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n487), .B1(new_n488), .B2(G136), .ZN(new_n489));
  AND2_X1   g064(.A1(new_n484), .A2(new_n489), .ZN(G162));
  OAI211_X1 g065(.A(G126), .B(G2105), .C1(new_n463), .C2(new_n464), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n493), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n462), .A2(G138), .ZN(new_n496));
  OAI21_X1  g071(.A(KEYINPUT4), .B1(new_n472), .B2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  INV_X1    g073(.A(new_n496), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n480), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n495), .B1(new_n497), .B2(new_n500), .ZN(G164));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n506), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n507));
  OR2_X1    g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT71), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  OR2_X1    g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g092(.A(KEYINPUT71), .B1(new_n507), .B2(new_n511), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n514), .A2(new_n517), .A3(new_n518), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  NAND3_X1  g095(.A1(new_n508), .A2(KEYINPUT72), .A3(new_n509), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT72), .ZN(new_n522));
  AND2_X1   g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  NOR2_X1   g098(.A1(KEYINPUT6), .A2(G651), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n521), .A2(new_n525), .A3(G543), .ZN(new_n526));
  INV_X1    g101(.A(G51), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n506), .A2(G63), .A3(G651), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n510), .A2(new_n506), .ZN(new_n532));
  INV_X1    g107(.A(G89), .ZN(new_n533));
  OAI211_X1 g108(.A(new_n529), .B(new_n531), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n528), .A2(new_n534), .ZN(G168));
  AOI22_X1  g110(.A1(new_n506), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n536), .A2(new_n516), .ZN(new_n537));
  AND3_X1   g112(.A1(new_n521), .A2(new_n525), .A3(G543), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G52), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n508), .A2(new_n509), .B1(new_n504), .B2(new_n505), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G90), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n537), .A2(new_n539), .A3(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  NAND2_X1  g118(.A1(new_n540), .A2(G81), .ZN(new_n544));
  INV_X1    g119(.A(G56), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n545), .B1(new_n504), .B2(new_n505), .ZN(new_n546));
  AND2_X1   g121(.A1(G68), .A2(G543), .ZN(new_n547));
  OAI21_X1  g122(.A(G651), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(G43), .ZN(new_n549));
  OAI211_X1 g124(.A(new_n544), .B(new_n548), .C1(new_n526), .C2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT73), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  AOI21_X1  g132(.A(new_n503), .B1(new_n510), .B2(new_n522), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT9), .ZN(new_n559));
  NAND4_X1  g134(.A1(new_n558), .A2(new_n559), .A3(G53), .A4(new_n521), .ZN(new_n560));
  NAND4_X1  g135(.A1(new_n521), .A2(new_n525), .A3(G53), .A4(G543), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(KEYINPUT9), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(G65), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n564), .B1(new_n504), .B2(new_n505), .ZN(new_n565));
  AND2_X1   g140(.A1(G78), .A2(G543), .ZN(new_n566));
  OAI21_X1  g141(.A(G651), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT75), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OAI211_X1 g144(.A(KEYINPUT75), .B(G651), .C1(new_n565), .C2(new_n566), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT74), .ZN(new_n572));
  INV_X1    g147(.A(G91), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n532), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n540), .A2(KEYINPUT74), .A3(G91), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n563), .A2(new_n571), .A3(new_n576), .ZN(G299));
  INV_X1    g152(.A(G168), .ZN(G286));
  OAI21_X1  g153(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n579));
  OR2_X1    g154(.A1(new_n579), .A2(KEYINPUT76), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n538), .A2(G49), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n579), .A2(KEYINPUT76), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n540), .A2(G87), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n580), .A2(new_n581), .A3(new_n582), .A4(new_n583), .ZN(G288));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  INV_X1    g160(.A(new_n505), .ZN(new_n586));
  NOR2_X1   g161(.A1(KEYINPUT5), .A2(G543), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(G61), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n585), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(G651), .ZN(new_n591));
  NAND2_X1  g166(.A1(G48), .A2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G86), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n588), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(new_n510), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n591), .A2(new_n595), .ZN(G305));
  NAND2_X1  g171(.A1(new_n540), .A2(G85), .ZN(new_n597));
  INV_X1    g172(.A(G60), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n598), .B1(new_n504), .B2(new_n505), .ZN(new_n599));
  AND2_X1   g174(.A1(G72), .A2(G543), .ZN(new_n600));
  OAI21_X1  g175(.A(G651), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n597), .B1(new_n601), .B2(KEYINPUT77), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(G47), .A2(new_n538), .B1(new_n601), .B2(KEYINPUT77), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n603), .A2(KEYINPUT78), .A3(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(new_n606));
  AOI21_X1  g181(.A(KEYINPUT78), .B1(new_n603), .B2(new_n604), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(G290));
  NAND2_X1  g184(.A1(G301), .A2(G868), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT10), .ZN(new_n611));
  INV_X1    g186(.A(G92), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n532), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n540), .A2(KEYINPUT10), .A3(G92), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n613), .A2(new_n614), .B1(new_n538), .B2(G54), .ZN(new_n615));
  INV_X1    g190(.A(G66), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n616), .B1(new_n504), .B2(new_n505), .ZN(new_n617));
  AND2_X1   g192(.A1(G79), .A2(G543), .ZN(new_n618));
  OR3_X1    g193(.A1(new_n617), .A2(KEYINPUT79), .A3(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(KEYINPUT79), .B1(new_n617), .B2(new_n618), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n619), .A2(G651), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n615), .A2(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n610), .B1(new_n623), .B2(G868), .ZN(G284));
  OAI21_X1  g199(.A(new_n610), .B1(new_n623), .B2(G868), .ZN(G321));
  NAND2_X1  g200(.A1(G286), .A2(G868), .ZN(new_n626));
  INV_X1    g201(.A(G299), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(G868), .ZN(G297));
  OAI21_X1  g203(.A(new_n626), .B1(new_n627), .B2(G868), .ZN(G280));
  INV_X1    g204(.A(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n623), .B1(new_n630), .B2(G860), .ZN(G148));
  OAI21_X1  g206(.A(KEYINPUT80), .B1(new_n551), .B2(G868), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n623), .A2(new_n630), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(G868), .ZN(new_n634));
  MUX2_X1   g209(.A(KEYINPUT80), .B(new_n632), .S(new_n634), .Z(G323));
  XNOR2_X1  g210(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g211(.A1(new_n480), .A2(new_n467), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT12), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT13), .ZN(new_n639));
  INV_X1    g214(.A(G2100), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  AOI22_X1  g217(.A1(new_n482), .A2(G123), .B1(new_n488), .B2(G135), .ZN(new_n643));
  OAI21_X1  g218(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n644));
  INV_X1    g219(.A(KEYINPUT81), .ZN(new_n645));
  INV_X1    g220(.A(G111), .ZN(new_n646));
  AOI22_X1  g221(.A1(new_n644), .A2(new_n645), .B1(new_n646), .B2(G2105), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n647), .B1(new_n645), .B2(new_n644), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n643), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(G2096), .Z(new_n650));
  NAND3_X1  g225(.A1(new_n641), .A2(new_n642), .A3(new_n650), .ZN(G156));
  XNOR2_X1  g226(.A(KEYINPUT15), .B(G2435), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2438), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2427), .B(G2430), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n655), .A2(KEYINPUT14), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT82), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n657), .B1(new_n653), .B2(new_n654), .ZN(new_n658));
  XOR2_X1   g233(.A(G2443), .B(G2446), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2451), .B(G2454), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT16), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n660), .A2(new_n663), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1341), .B(G1348), .ZN(new_n667));
  OAI21_X1  g242(.A(KEYINPUT83), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(KEYINPUT83), .ZN(new_n669));
  INV_X1    g244(.A(new_n667), .ZN(new_n670));
  NAND4_X1  g245(.A1(new_n664), .A2(new_n665), .A3(new_n669), .A4(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(G14), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(new_n666), .B2(new_n667), .ZN(new_n674));
  AND2_X1   g249(.A1(new_n672), .A2(new_n674), .ZN(G401));
  XOR2_X1   g250(.A(G2084), .B(G2090), .Z(new_n676));
  XNOR2_X1  g251(.A(G2067), .B(G2678), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT84), .Z(new_n678));
  NOR2_X1   g253(.A1(G2072), .A2(G2078), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n442), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n676), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(KEYINPUT17), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n681), .B1(new_n678), .B2(new_n682), .ZN(new_n683));
  OAI211_X1 g258(.A(new_n676), .B(new_n677), .C1(new_n442), .C2(new_n679), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT18), .Z(new_n685));
  NAND3_X1  g260(.A1(new_n678), .A2(new_n682), .A3(new_n676), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n683), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(G2096), .B(G2100), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(G227));
  XNOR2_X1  g264(.A(G1981), .B(G1986), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(G1971), .B(G1976), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT19), .ZN(new_n693));
  XOR2_X1   g268(.A(G1956), .B(G2474), .Z(new_n694));
  XOR2_X1   g269(.A(G1961), .B(G1966), .Z(new_n695));
  NAND3_X1  g270(.A1(new_n694), .A2(new_n695), .A3(KEYINPUT85), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n694), .A2(new_n695), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT85), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n693), .A2(new_n696), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT20), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n694), .A2(new_n695), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n693), .A2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n702), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(new_n697), .ZN(new_n705));
  OAI211_X1 g280(.A(new_n701), .B(new_n703), .C1(new_n693), .C2(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(G1991), .B(G1996), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT86), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n708), .A2(new_n711), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n691), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n714), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n716), .A2(new_n712), .A3(new_n690), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n715), .A2(new_n717), .ZN(G229));
  INV_X1    g293(.A(G16), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G23), .ZN(new_n720));
  INV_X1    g295(.A(G288), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n720), .B1(new_n721), .B2(new_n719), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT33), .B(G1976), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n724), .A2(KEYINPUT91), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(KEYINPUT91), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n719), .A2(G22), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G166), .B2(new_n719), .ZN(new_n728));
  INV_X1    g303(.A(G1971), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n719), .A2(G6), .ZN(new_n731));
  INV_X1    g306(.A(G305), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n731), .B1(new_n732), .B2(new_n719), .ZN(new_n733));
  XOR2_X1   g308(.A(KEYINPUT32), .B(G1981), .Z(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT90), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n733), .B(new_n735), .ZN(new_n736));
  NAND4_X1  g311(.A1(new_n725), .A2(new_n726), .A3(new_n730), .A4(new_n736), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT89), .B(KEYINPUT34), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(G29), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(G25), .ZN(new_n741));
  OAI21_X1  g316(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n742));
  INV_X1    g317(.A(G107), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n742), .B1(new_n743), .B2(G2105), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT87), .ZN(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(G119), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n480), .A2(new_n462), .ZN(new_n748));
  INV_X1    g323(.A(G131), .ZN(new_n749));
  OAI22_X1  g324(.A1(new_n747), .A2(new_n481), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n746), .A2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n741), .B1(new_n752), .B2(new_n740), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT35), .B(G1991), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT88), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n753), .B(new_n755), .Z(new_n756));
  NAND2_X1  g331(.A1(new_n719), .A2(G24), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n608), .B2(new_n719), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n758), .A2(G1986), .ZN(new_n759));
  AND2_X1   g334(.A1(new_n758), .A2(G1986), .ZN(new_n760));
  NOR3_X1   g335(.A1(new_n756), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n737), .A2(new_n738), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n739), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(KEYINPUT92), .A2(KEYINPUT36), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  OR2_X1    g340(.A1(KEYINPUT92), .A2(KEYINPUT36), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n763), .A2(new_n764), .A3(new_n766), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT25), .Z(new_n769));
  INV_X1    g344(.A(G139), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n769), .B1(new_n770), .B2(new_n748), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT95), .ZN(new_n772));
  AOI22_X1  g347(.A1(new_n480), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n772), .B1(new_n462), .B2(new_n773), .ZN(new_n774));
  MUX2_X1   g349(.A(G33), .B(new_n774), .S(G29), .Z(new_n775));
  AND2_X1   g350(.A1(new_n775), .A2(G2072), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n775), .A2(G2072), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT31), .B(G11), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT98), .B(G28), .ZN(new_n779));
  INV_X1    g354(.A(KEYINPUT30), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n740), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT99), .ZN(new_n782));
  AND2_X1   g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n779), .A2(new_n780), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n781), .B2(new_n782), .ZN(new_n785));
  OAI221_X1 g360(.A(new_n778), .B1(new_n783), .B2(new_n785), .C1(new_n649), .C2(new_n740), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n740), .A2(G32), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n462), .A2(G105), .A3(G2104), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT96), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(G141), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n790), .B1(new_n791), .B2(new_n748), .ZN(new_n792));
  NAND3_X1  g367(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n793), .A2(KEYINPUT26), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n793), .A2(KEYINPUT26), .ZN(new_n795));
  INV_X1    g370(.A(G129), .ZN(new_n796));
  OAI211_X1 g371(.A(new_n794), .B(new_n795), .C1(new_n481), .C2(new_n796), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n792), .A2(new_n797), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n787), .B1(new_n798), .B2(new_n740), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  XNOR2_X1  g375(.A(KEYINPUT27), .B(G1996), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n786), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(new_n800), .B2(new_n801), .ZN(new_n803));
  NOR3_X1   g378(.A1(new_n776), .A2(new_n777), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n719), .A2(G5), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G171), .B2(new_n719), .ZN(new_n806));
  INV_X1    g381(.A(G1961), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(G29), .A2(G35), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G162), .B2(G29), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT29), .B(G2090), .Z(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n740), .A2(G26), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT94), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT28), .ZN(new_n815));
  OR2_X1    g390(.A1(G104), .A2(G2105), .ZN(new_n816));
  OAI211_X1 g391(.A(new_n816), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT93), .Z(new_n818));
  AOI22_X1  g393(.A1(new_n482), .A2(G128), .B1(new_n488), .B2(G140), .ZN(new_n819));
  AND2_X1   g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n815), .B1(new_n820), .B2(new_n740), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(G2067), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n740), .A2(G27), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(G164), .B2(new_n740), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(G2078), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n719), .A2(G19), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(new_n551), .B2(new_n719), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(G1341), .ZN(new_n828));
  NOR3_X1   g403(.A1(new_n822), .A2(new_n825), .A3(new_n828), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n804), .A2(new_n808), .A3(new_n812), .A4(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(G34), .ZN(new_n831));
  AND2_X1   g406(.A1(new_n831), .A2(KEYINPUT24), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n831), .A2(KEYINPUT24), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n740), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(G160), .B2(new_n740), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(G2084), .ZN(new_n836));
  XOR2_X1   g411(.A(KEYINPUT100), .B(KEYINPUT23), .Z(new_n837));
  NAND2_X1  g412(.A1(new_n719), .A2(G20), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n839), .B1(new_n627), .B2(new_n719), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(G1956), .ZN(new_n841));
  NOR2_X1   g416(.A1(G16), .A2(G21), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n842), .B1(G168), .B2(G16), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT97), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n844), .A2(G1966), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n719), .A2(G4), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n846), .B1(new_n623), .B2(new_n719), .ZN(new_n847));
  INV_X1    g422(.A(G1348), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n844), .A2(G1966), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n845), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  NOR4_X1   g426(.A1(new_n830), .A2(new_n836), .A3(new_n841), .A4(new_n851), .ZN(new_n852));
  AND3_X1   g427(.A1(new_n765), .A2(new_n767), .A3(new_n852), .ZN(G311));
  NAND3_X1  g428(.A1(new_n765), .A2(new_n767), .A3(new_n852), .ZN(G150));
  NAND2_X1  g429(.A1(new_n623), .A2(G559), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT38), .ZN(new_n856));
  INV_X1    g431(.A(G67), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n857), .B1(new_n504), .B2(new_n505), .ZN(new_n858));
  NAND2_X1  g433(.A1(G80), .A2(G543), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  OAI21_X1  g435(.A(KEYINPUT101), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT101), .ZN(new_n862));
  OAI211_X1 g437(.A(new_n862), .B(new_n859), .C1(new_n588), .C2(new_n857), .ZN(new_n863));
  AND3_X1   g438(.A1(new_n861), .A2(new_n863), .A3(G651), .ZN(new_n864));
  INV_X1    g439(.A(G55), .ZN(new_n865));
  INV_X1    g440(.A(G93), .ZN(new_n866));
  OAI22_X1  g441(.A1(new_n526), .A2(new_n865), .B1(new_n866), .B2(new_n532), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n550), .B1(new_n864), .B2(new_n867), .ZN(new_n868));
  AOI22_X1  g443(.A1(new_n538), .A2(G55), .B1(G93), .B2(new_n540), .ZN(new_n869));
  AND2_X1   g444(.A1(new_n544), .A2(new_n548), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n538), .A2(G43), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n861), .A2(new_n863), .A3(G651), .ZN(new_n872));
  NAND4_X1  g447(.A1(new_n869), .A2(new_n870), .A3(new_n871), .A4(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n868), .A2(new_n873), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n856), .B(new_n874), .Z(new_n875));
  OR2_X1    g450(.A1(new_n875), .A2(KEYINPUT39), .ZN(new_n876));
  INV_X1    g451(.A(G860), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n875), .A2(KEYINPUT39), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n877), .B1(new_n869), .B2(new_n872), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT37), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(G145));
  XNOR2_X1  g457(.A(new_n798), .B(G164), .ZN(new_n883));
  OR2_X1    g458(.A1(new_n883), .A2(new_n820), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n820), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT102), .ZN(new_n886));
  OAI211_X1 g461(.A(new_n884), .B(new_n885), .C1(new_n886), .C2(new_n774), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n751), .B(new_n638), .ZN(new_n888));
  OR2_X1    g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n774), .A2(new_n886), .ZN(new_n890));
  AOI22_X1  g465(.A1(new_n482), .A2(G130), .B1(new_n488), .B2(G142), .ZN(new_n891));
  OAI21_X1  g466(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n892));
  INV_X1    g467(.A(G118), .ZN(new_n893));
  AOI22_X1  g468(.A1(new_n892), .A2(KEYINPUT103), .B1(new_n893), .B2(G2105), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n894), .B1(KEYINPUT103), .B2(new_n892), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n891), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n890), .B(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n887), .A2(new_n888), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n889), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n897), .B1(new_n889), .B2(new_n898), .ZN(new_n901));
  OR2_X1    g476(.A1(G160), .A2(new_n649), .ZN(new_n902));
  NAND2_X1  g477(.A1(G160), .A2(new_n649), .ZN(new_n903));
  AND3_X1   g478(.A1(new_n902), .A2(G162), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(G162), .B1(new_n902), .B2(new_n903), .ZN(new_n905));
  OAI22_X1  g480(.A1(new_n900), .A2(new_n901), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n901), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n904), .A2(new_n905), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n907), .A2(new_n908), .A3(new_n899), .ZN(new_n909));
  INV_X1    g484(.A(G37), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n906), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g487(.A(G868), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n913), .B1(new_n864), .B2(new_n867), .ZN(new_n914));
  NAND2_X1  g489(.A1(G166), .A2(G305), .ZN(new_n915));
  NAND2_X1  g490(.A1(G303), .A2(new_n732), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT78), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n601), .A2(KEYINPUT77), .ZN(new_n919));
  INV_X1    g494(.A(G47), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n919), .B1(new_n920), .B2(new_n526), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n918), .B1(new_n921), .B2(new_n602), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n922), .A2(G288), .A3(new_n605), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(G288), .B1(new_n922), .B2(new_n605), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n917), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n721), .B1(new_n606), .B2(new_n607), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n927), .A2(new_n916), .A3(new_n915), .A4(new_n923), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n929), .B1(KEYINPUT105), .B2(KEYINPUT42), .ZN(new_n930));
  NAND2_X1  g505(.A1(KEYINPUT105), .A2(KEYINPUT42), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n930), .B(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(G299), .A2(new_n622), .ZN(new_n933));
  AOI22_X1  g508(.A1(new_n569), .A2(new_n570), .B1(new_n574), .B2(new_n575), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n934), .A2(new_n563), .A3(new_n621), .A4(new_n615), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(KEYINPUT104), .B(KEYINPUT41), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT41), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n933), .A2(new_n941), .A3(new_n935), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  XOR2_X1   g518(.A(new_n633), .B(new_n874), .Z(new_n944));
  MUX2_X1   g519(.A(new_n937), .B(new_n943), .S(new_n944), .Z(new_n945));
  XNOR2_X1  g520(.A(new_n932), .B(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n914), .B1(new_n946), .B2(new_n913), .ZN(G295));
  OAI21_X1  g522(.A(new_n914), .B1(new_n946), .B2(new_n913), .ZN(G331));
  INV_X1    g523(.A(KEYINPUT44), .ZN(new_n949));
  AOI21_X1  g524(.A(G301), .B1(KEYINPUT106), .B2(G168), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT106), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n952), .B1(new_n528), .B2(new_n534), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n868), .A2(new_n873), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n953), .B1(new_n868), .B2(new_n873), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n951), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n953), .ZN(new_n957));
  NOR3_X1   g532(.A1(new_n864), .A2(new_n550), .A3(new_n867), .ZN(new_n958));
  AOI22_X1  g533(.A1(new_n869), .A2(new_n872), .B1(new_n870), .B2(new_n871), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n957), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n868), .A2(new_n873), .A3(new_n953), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n960), .A2(new_n950), .A3(new_n961), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n956), .A2(new_n962), .A3(new_n937), .ZN(new_n963));
  AOI22_X1  g538(.A1(new_n956), .A2(new_n962), .B1(new_n940), .B2(new_n942), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(G37), .B1(new_n965), .B2(new_n929), .ZN(new_n966));
  AND2_X1   g541(.A1(new_n926), .A2(new_n928), .ZN(new_n967));
  NOR2_X1   g542(.A1(G299), .A2(new_n622), .ZN(new_n968));
  AOI22_X1  g543(.A1(new_n934), .A2(new_n563), .B1(new_n615), .B2(new_n621), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n941), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n933), .A2(new_n935), .A3(new_n939), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n972), .B1(new_n962), .B2(new_n956), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n967), .B1(new_n973), .B2(new_n963), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n966), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n949), .B1(new_n975), .B2(KEYINPUT43), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n967), .B1(new_n963), .B2(new_n964), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n956), .A2(new_n962), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(new_n943), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n956), .A2(new_n962), .A3(new_n937), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n979), .A2(new_n929), .A3(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n977), .A2(new_n981), .A3(new_n910), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n976), .B1(KEYINPUT43), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT43), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n974), .A2(new_n984), .A3(new_n910), .A4(new_n981), .ZN(new_n985));
  AOI22_X1  g560(.A1(new_n985), .A2(KEYINPUT107), .B1(new_n982), .B2(KEYINPUT43), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT107), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n966), .A2(new_n987), .A3(new_n984), .A4(new_n974), .ZN(new_n988));
  AOI211_X1 g563(.A(KEYINPUT108), .B(KEYINPUT44), .C1(new_n986), .C2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT108), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n985), .A2(KEYINPUT107), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n991), .A2(new_n988), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n990), .B1(new_n993), .B2(new_n949), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n983), .B1(new_n989), .B2(new_n994), .ZN(G397));
  XNOR2_X1  g570(.A(new_n820), .B(G2067), .ZN(new_n996));
  OAI21_X1  g571(.A(G1996), .B1(new_n792), .B2(new_n797), .ZN(new_n997));
  INV_X1    g572(.A(G1996), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n798), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n996), .A2(new_n997), .A3(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n473), .B1(new_n478), .B2(new_n479), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n474), .A2(new_n466), .ZN(new_n1002));
  OAI21_X1  g577(.A(G2105), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  AND3_X1   g578(.A1(new_n465), .A2(KEYINPUT68), .A3(new_n468), .ZN(new_n1004));
  OAI211_X1 g579(.A(G40), .B(new_n1003), .C1(new_n1004), .C2(new_n469), .ZN(new_n1005));
  XOR2_X1   g580(.A(KEYINPUT109), .B(G1384), .Z(new_n1006));
  NAND2_X1  g581(.A1(new_n497), .A2(new_n500), .ZN(new_n1007));
  AND2_X1   g582(.A1(new_n491), .A2(new_n494), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1006), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NOR3_X1   g584(.A1(new_n1005), .A2(new_n1009), .A3(KEYINPUT45), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1000), .A2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n1011), .B(KEYINPUT110), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1010), .ZN(new_n1013));
  OR2_X1    g588(.A1(new_n752), .A2(new_n755), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n752), .A2(new_n755), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1013), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  OR2_X1    g591(.A1(new_n1012), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G1986), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n608), .B(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1017), .B1(new_n1010), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT111), .ZN(new_n1021));
  AOI21_X1  g596(.A(G1384), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1021), .B1(new_n1022), .B2(KEYINPUT45), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1005), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT45), .ZN(new_n1025));
  OAI211_X1 g600(.A(KEYINPUT111), .B(new_n1025), .C1(G164), .C2(G1384), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1009), .A2(KEYINPUT45), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1023), .A2(new_n1024), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n729), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1030));
  INV_X1    g605(.A(G1384), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1005), .B1(new_n1032), .B2(KEYINPUT50), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT50), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1022), .A2(new_n1034), .ZN(new_n1035));
  XOR2_X1   g610(.A(KEYINPUT112), .B(G2090), .Z(new_n1036));
  NAND3_X1  g611(.A1(new_n1033), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1029), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT113), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(G303), .A2(G8), .ZN(new_n1041));
  XNOR2_X1  g616(.A(new_n1041), .B(KEYINPUT55), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1029), .A2(KEYINPUT113), .A3(new_n1037), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1040), .A2(new_n1043), .A3(new_n1044), .A4(G8), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT49), .ZN(new_n1046));
  INV_X1    g621(.A(G1981), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n591), .A2(new_n595), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT114), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1046), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1048), .A2(new_n1049), .A3(new_n1046), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1051), .B(new_n1052), .C1(new_n1047), .C2(new_n732), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1032), .A2(new_n1005), .ZN(new_n1054));
  INV_X1    g629(.A(G8), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n732), .A2(new_n1047), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1052), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1057), .B1(new_n1058), .B2(new_n1050), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1053), .A2(new_n1056), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(G1976), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1056), .B1(new_n1061), .B2(G288), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT52), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT52), .B1(G288), .B2(new_n1061), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1056), .B(new_n1064), .C1(new_n1061), .C2(G288), .ZN(new_n1065));
  AND3_X1   g640(.A1(new_n1060), .A2(new_n1063), .A3(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(KEYINPUT116), .B1(new_n1022), .B2(new_n1034), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT116), .ZN(new_n1068));
  NOR4_X1   g643(.A1(G164), .A2(new_n1068), .A3(KEYINPUT50), .A4(G1384), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1033), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  AOI22_X1  g646(.A1(new_n1071), .A2(new_n1036), .B1(new_n729), .B2(new_n1028), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1042), .B1(new_n1072), .B2(new_n1055), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1045), .A2(new_n1066), .A3(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1032), .A2(new_n1025), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1022), .A2(KEYINPUT45), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1075), .A2(new_n1024), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(G1966), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(G2084), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1033), .A2(new_n1080), .A3(new_n1035), .ZN(new_n1081));
  AND2_X1   g656(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  NOR2_X1   g657(.A1(G168), .A2(new_n1055), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(KEYINPUT51), .B1(new_n1083), .B2(KEYINPUT122), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1084), .B(new_n1086), .C1(new_n1082), .C2(new_n1055), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1086), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1089));
  OAI211_X1 g664(.A(G8), .B(new_n1088), .C1(new_n1089), .C2(G286), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1085), .B1(new_n1087), .B2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1074), .A2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1005), .B1(KEYINPUT45), .B2(new_n1009), .ZN(new_n1093));
  INV_X1    g668(.A(G2078), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1093), .A2(new_n1094), .A3(new_n1023), .A4(new_n1026), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT53), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1096), .A2(G2078), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1075), .A2(new_n1024), .A3(new_n1098), .A4(new_n1076), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(new_n807), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1097), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(G171), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT123), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT123), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1102), .A2(new_n1105), .A3(G171), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1009), .A2(KEYINPUT45), .ZN(new_n1107));
  NOR3_X1   g682(.A1(new_n1107), .A2(new_n1096), .A3(G2078), .ZN(new_n1108));
  OR2_X1    g683(.A1(new_n1024), .A2(KEYINPUT124), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1024), .A2(KEYINPUT124), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1108), .A2(new_n1109), .A3(new_n1027), .A4(new_n1110), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1111), .A2(new_n1097), .A3(G301), .A4(new_n1101), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1104), .A2(new_n1106), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT54), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1111), .A2(new_n1097), .A3(new_n1101), .ZN(new_n1116));
  AOI21_X1  g691(.A(G301), .B1(new_n1116), .B2(KEYINPUT125), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1117), .B1(KEYINPUT125), .B2(new_n1116), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1102), .A2(G171), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1119), .A2(new_n1114), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1092), .A2(new_n1115), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT57), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n934), .A2(new_n1124), .A3(new_n563), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1035), .A2(new_n1068), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1022), .A2(KEYINPUT116), .A3(new_n1034), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(G1956), .B1(new_n1129), .B2(new_n1033), .ZN(new_n1130));
  XNOR2_X1  g705(.A(KEYINPUT56), .B(G2072), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1093), .A2(new_n1023), .A3(new_n1026), .A4(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1126), .B1(new_n1130), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT117), .ZN(new_n1135));
  AOI21_X1  g710(.A(G1348), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1024), .A2(new_n1022), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1137), .A2(G2067), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1135), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n476), .B(G40), .C1(new_n1022), .C2(new_n1034), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1035), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n848), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(G2067), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1054), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1142), .A2(KEYINPUT117), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1139), .A2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1134), .B1(new_n1146), .B2(new_n622), .ZN(new_n1147));
  INV_X1    g722(.A(G1956), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1070), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1126), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1149), .A2(new_n1150), .A3(new_n1132), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1147), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT119), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(KEYINPUT61), .ZN(new_n1154));
  NOR3_X1   g729(.A1(new_n1130), .A2(new_n1133), .A3(new_n1126), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1150), .B1(new_n1149), .B2(new_n1132), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1154), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  XOR2_X1   g732(.A(KEYINPUT119), .B(KEYINPUT61), .Z(new_n1158));
  NAND3_X1  g733(.A1(new_n1134), .A2(new_n1151), .A3(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g734(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1093), .A2(new_n998), .A3(new_n1023), .A4(new_n1026), .ZN(new_n1161));
  XOR2_X1   g736(.A(KEYINPUT58), .B(G1341), .Z(new_n1162));
  NAND2_X1  g737(.A1(new_n1137), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1160), .B1(new_n1164), .B2(new_n551), .ZN(new_n1165));
  NAND2_X1  g740(.A1(KEYINPUT118), .A2(KEYINPUT59), .ZN(new_n1166));
  AOI211_X1 g741(.A(new_n550), .B(new_n1166), .C1(new_n1161), .C2(new_n1163), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1157), .A2(new_n1159), .A3(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT120), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1146), .A2(KEYINPUT60), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT60), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1139), .A2(new_n1145), .A3(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT121), .ZN(new_n1175));
  AND3_X1   g750(.A1(new_n1174), .A2(new_n1175), .A3(new_n623), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1175), .B1(new_n1174), .B2(new_n623), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1172), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1174), .A2(new_n623), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1179), .A2(KEYINPUT121), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1172), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1174), .A2(new_n1175), .A3(new_n623), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1180), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  NAND4_X1  g758(.A1(new_n1157), .A2(new_n1168), .A3(new_n1159), .A4(KEYINPUT120), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1171), .A2(new_n1178), .A3(new_n1183), .A4(new_n1184), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1122), .B1(new_n1152), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1187));
  INV_X1    g762(.A(new_n1074), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n1091), .A2(KEYINPUT62), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT62), .ZN(new_n1190));
  AOI211_X1 g765(.A(new_n1190), .B(new_n1085), .C1(new_n1087), .C2(new_n1090), .ZN(new_n1191));
  OAI211_X1 g766(.A(new_n1187), .B(new_n1188), .C1(new_n1189), .C2(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT63), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1089), .A2(G8), .A3(G168), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1193), .B1(new_n1074), .B2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1040), .A2(G8), .A3(new_n1044), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1196), .A2(new_n1042), .ZN(new_n1197));
  NOR2_X1   g772(.A1(new_n1194), .A2(new_n1193), .ZN(new_n1198));
  NAND4_X1  g773(.A1(new_n1197), .A2(new_n1045), .A3(new_n1066), .A4(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1195), .A2(new_n1199), .ZN(new_n1200));
  INV_X1    g775(.A(new_n1045), .ZN(new_n1201));
  AND2_X1   g776(.A1(new_n1053), .A2(new_n1059), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n721), .A2(new_n1061), .ZN(new_n1203));
  XNOR2_X1  g778(.A(new_n1203), .B(KEYINPUT115), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1048), .B1(new_n1202), .B2(new_n1204), .ZN(new_n1205));
  AOI22_X1  g780(.A1(new_n1201), .A2(new_n1066), .B1(new_n1056), .B2(new_n1205), .ZN(new_n1206));
  NAND3_X1  g781(.A1(new_n1192), .A2(new_n1200), .A3(new_n1206), .ZN(new_n1207));
  OAI21_X1  g782(.A(new_n1020), .B1(new_n1186), .B2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g783(.A(new_n1013), .B1(new_n996), .B2(new_n798), .ZN(new_n1209));
  XNOR2_X1  g784(.A(new_n1209), .B(KEYINPUT126), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1010), .A2(new_n998), .ZN(new_n1211));
  XOR2_X1   g786(.A(new_n1211), .B(KEYINPUT46), .Z(new_n1212));
  NOR2_X1   g787(.A1(new_n1210), .A2(new_n1212), .ZN(new_n1213));
  XNOR2_X1  g788(.A(KEYINPUT127), .B(KEYINPUT47), .ZN(new_n1214));
  XNOR2_X1  g789(.A(new_n1213), .B(new_n1214), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n820), .A2(new_n1143), .ZN(new_n1216));
  OAI21_X1  g791(.A(new_n1216), .B1(new_n1012), .B2(new_n1015), .ZN(new_n1217));
  AND2_X1   g792(.A1(new_n1217), .A2(new_n1010), .ZN(new_n1218));
  NAND3_X1  g793(.A1(new_n608), .A2(new_n1018), .A3(new_n1010), .ZN(new_n1219));
  XOR2_X1   g794(.A(new_n1219), .B(KEYINPUT48), .Z(new_n1220));
  NOR2_X1   g795(.A1(new_n1017), .A2(new_n1220), .ZN(new_n1221));
  NOR3_X1   g796(.A1(new_n1215), .A2(new_n1218), .A3(new_n1221), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1208), .A2(new_n1222), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g798(.A1(G227), .A2(new_n460), .ZN(new_n1225));
  NAND3_X1  g799(.A1(new_n715), .A2(new_n717), .A3(new_n1225), .ZN(new_n1226));
  AOI21_X1  g800(.A(new_n1226), .B1(new_n672), .B2(new_n674), .ZN(new_n1227));
  AND3_X1   g801(.A1(new_n1227), .A2(new_n911), .A3(new_n993), .ZN(G308));
  NAND3_X1  g802(.A1(new_n1227), .A2(new_n911), .A3(new_n993), .ZN(G225));
endmodule


