

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741;

  NOR2_X1 U375 ( .A1(n741), .A2(n740), .ZN(n555) );
  NOR2_X1 U376 ( .A1(n409), .A2(n536), .ZN(n657) );
  XNOR2_X1 U377 ( .A(n584), .B(n583), .ZN(n383) );
  XNOR2_X1 U378 ( .A(n410), .B(KEYINPUT101), .ZN(n651) );
  AND2_X1 U379 ( .A1(n537), .A2(n542), .ZN(n410) );
  XNOR2_X1 U380 ( .A(n675), .B(KEYINPUT105), .ZN(n586) );
  NOR2_X1 U381 ( .A1(n671), .A2(n531), .ZN(n546) );
  XNOR2_X1 U382 ( .A(n472), .B(n473), .ZN(n537) );
  NOR2_X1 U383 ( .A1(n709), .A2(G902), .ZN(n372) );
  XNOR2_X1 U384 ( .A(n352), .B(n467), .ZN(n469) );
  XNOR2_X1 U385 ( .A(n444), .B(G131), .ZN(n483) );
  NOR2_X1 U386 ( .A1(G953), .A2(G237), .ZN(n486) );
  INV_X1 U387 ( .A(n466), .ZN(n352) );
  XNOR2_X2 U388 ( .A(n375), .B(n712), .ZN(n631) );
  AND2_X2 U389 ( .A1(n552), .A2(n551), .ZN(n553) );
  NAND2_X2 U390 ( .A1(n369), .A2(n366), .ZN(n727) );
  XNOR2_X1 U391 ( .A(n379), .B(n353), .ZN(n378) );
  XNOR2_X1 U392 ( .A(n517), .B(n404), .ZN(n353) );
  INV_X2 U393 ( .A(G953), .ZN(n728) );
  NOR2_X1 U394 ( .A1(n600), .A2(n601), .ZN(n637) );
  XNOR2_X2 U395 ( .A(n450), .B(n359), .ZN(n551) );
  AND2_X2 U396 ( .A1(n547), .A2(n586), .ZN(n550) );
  XNOR2_X2 U397 ( .A(n372), .B(n357), .ZN(n588) );
  INV_X1 U398 ( .A(KEYINPUT67), .ZN(n444) );
  XOR2_X1 U399 ( .A(KEYINPUT4), .B(G146), .Z(n517) );
  AND2_X1 U400 ( .A1(n390), .A2(n397), .ZN(n396) );
  NAND2_X1 U401 ( .A1(n738), .A2(KEYINPUT44), .ZN(n390) );
  XNOR2_X1 U402 ( .A(n507), .B(n506), .ZN(n677) );
  XNOR2_X1 U403 ( .A(n633), .B(n632), .ZN(n634) );
  XNOR2_X1 U404 ( .A(n378), .B(n376), .ZN(n375) );
  XNOR2_X1 U405 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U406 ( .A(n405), .B(G110), .ZN(n519) );
  XNOR2_X1 U407 ( .A(n553), .B(KEYINPUT109), .ZN(n557) );
  XNOR2_X1 U408 ( .A(n725), .B(n490), .ZN(n617) );
  XNOR2_X2 U409 ( .A(n432), .B(KEYINPUT22), .ZN(n585) );
  NOR2_X2 U410 ( .A1(n605), .A2(n423), .ZN(n432) );
  XNOR2_X1 U411 ( .A(n374), .B(G140), .ZN(n726) );
  XNOR2_X1 U412 ( .A(n377), .B(n518), .ZN(n376) );
  OR2_X2 U413 ( .A1(n703), .A2(G902), .ZN(n450) );
  XOR2_X1 U414 ( .A(G122), .B(G107), .Z(n520) );
  XNOR2_X1 U415 ( .A(n425), .B(n517), .ZN(n485) );
  XNOR2_X1 U416 ( .A(n483), .B(n426), .ZN(n425) );
  INV_X1 U417 ( .A(G137), .ZN(n426) );
  XNOR2_X1 U418 ( .A(n481), .B(n480), .ZN(n542) );
  XNOR2_X1 U419 ( .A(KEYINPUT100), .B(G478), .ZN(n480) );
  INV_X1 U420 ( .A(n610), .ZN(n399) );
  XNOR2_X1 U421 ( .A(KEYINPUT5), .B(KEYINPUT94), .ZN(n487) );
  XOR2_X1 U422 ( .A(G113), .B(KEYINPUT95), .Z(n488) );
  INV_X1 U423 ( .A(KEYINPUT48), .ZN(n370) );
  XNOR2_X1 U424 ( .A(n442), .B(n441), .ZN(n523) );
  XNOR2_X1 U425 ( .A(G116), .B(KEYINPUT3), .ZN(n441) );
  XNOR2_X1 U426 ( .A(n443), .B(n451), .ZN(n442) );
  INV_X1 U427 ( .A(G119), .ZN(n451) );
  XNOR2_X1 U428 ( .A(n525), .B(n519), .ZN(n379) );
  XOR2_X1 U429 ( .A(KEYINPUT89), .B(KEYINPUT90), .Z(n525) );
  NAND2_X1 U430 ( .A1(G898), .A2(G953), .ZN(n579) );
  INV_X1 U431 ( .A(KEYINPUT19), .ZN(n386) );
  OR2_X2 U432 ( .A1(n435), .A2(n437), .ZN(n675) );
  NOR2_X1 U433 ( .A1(n617), .A2(n436), .ZN(n435) );
  NAND2_X1 U434 ( .A1(G472), .A2(n500), .ZN(n436) );
  XNOR2_X1 U435 ( .A(n726), .B(n470), .ZN(n494) );
  INV_X1 U436 ( .A(G146), .ZN(n470) );
  INV_X1 U437 ( .A(KEYINPUT39), .ZN(n420) );
  NOR2_X1 U438 ( .A1(n577), .A2(n412), .ZN(n411) );
  NAND2_X1 U439 ( .A1(n580), .A2(n424), .ZN(n423) );
  XNOR2_X1 U440 ( .A(n475), .B(n474), .ZN(n476) );
  AND2_X2 U441 ( .A1(n616), .A2(n615), .ZN(n707) );
  XNOR2_X1 U442 ( .A(n725), .B(n408), .ZN(n703) );
  XNOR2_X1 U443 ( .A(n509), .B(n365), .ZN(n408) );
  XNOR2_X1 U444 ( .A(n427), .B(n519), .ZN(n509) );
  NOR2_X1 U445 ( .A1(G952), .A2(n728), .ZN(n711) );
  XNOR2_X1 U446 ( .A(n544), .B(KEYINPUT41), .ZN(n697) );
  NOR2_X1 U447 ( .A1(n666), .A2(n665), .ZN(n544) );
  XNOR2_X1 U448 ( .A(G101), .B(KEYINPUT69), .ZN(n443) );
  OR2_X1 U449 ( .A1(G237), .A2(G902), .ZN(n526) );
  NAND2_X1 U450 ( .A1(n440), .A2(G902), .ZN(n438) );
  NAND2_X1 U451 ( .A1(n398), .A2(n396), .ZN(n395) );
  AND2_X1 U452 ( .A1(n394), .A2(n393), .ZN(n392) );
  NAND2_X1 U453 ( .A1(n637), .A2(KEYINPUT84), .ZN(n394) );
  XNOR2_X1 U454 ( .A(G125), .B(KEYINPUT10), .ZN(n374) );
  XNOR2_X1 U455 ( .A(G143), .B(G122), .ZN(n464) );
  XOR2_X1 U456 ( .A(KEYINPUT12), .B(KEYINPUT98), .Z(n465) );
  XOR2_X1 U457 ( .A(KEYINPUT97), .B(KEYINPUT11), .Z(n463) );
  INV_X1 U458 ( .A(KEYINPUT74), .ZN(n433) );
  XNOR2_X1 U459 ( .A(G125), .B(n453), .ZN(n404) );
  INV_X1 U460 ( .A(KEYINPUT75), .ZN(n453) );
  XNOR2_X1 U461 ( .A(n459), .B(n524), .ZN(n377) );
  XNOR2_X1 U462 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n524) );
  AND2_X1 U463 ( .A1(G224), .A2(n728), .ZN(n459) );
  XNOR2_X1 U464 ( .A(n388), .B(G143), .ZN(n518) );
  XNOR2_X1 U465 ( .A(G128), .B(KEYINPUT78), .ZN(n388) );
  XNOR2_X1 U466 ( .A(n556), .B(n429), .ZN(n400) );
  INV_X1 U467 ( .A(KEYINPUT38), .ZN(n429) );
  INV_X1 U468 ( .A(n601), .ZN(n577) );
  XNOR2_X1 U469 ( .A(n551), .B(n355), .ZN(n676) );
  XNOR2_X1 U470 ( .A(n417), .B(n523), .ZN(n490) );
  XNOR2_X1 U471 ( .A(n489), .B(n457), .ZN(n417) );
  XNOR2_X1 U472 ( .A(n371), .B(n370), .ZN(n369) );
  XNOR2_X1 U473 ( .A(n382), .B(n520), .ZN(n381) );
  XNOR2_X1 U474 ( .A(n521), .B(n522), .ZN(n382) );
  XOR2_X1 U475 ( .A(KEYINPUT72), .B(KEYINPUT16), .Z(n522) );
  XNOR2_X1 U476 ( .A(n414), .B(n413), .ZN(n493) );
  INV_X1 U477 ( .A(KEYINPUT8), .ZN(n413) );
  NAND2_X1 U478 ( .A1(n728), .A2(G234), .ZN(n414) );
  XNOR2_X1 U479 ( .A(n495), .B(KEYINPUT92), .ZN(n419) );
  XNOR2_X1 U480 ( .A(G119), .B(G110), .ZN(n495) );
  XNOR2_X1 U481 ( .A(G137), .B(G128), .ZN(n497) );
  XOR2_X1 U482 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n475) );
  INV_X1 U483 ( .A(KEYINPUT99), .ZN(n474) );
  XNOR2_X1 U484 ( .A(n518), .B(n479), .ZN(n484) );
  INV_X1 U485 ( .A(G134), .ZN(n479) );
  INV_X1 U486 ( .A(KEYINPUT70), .ZN(n405) );
  XNOR2_X1 U487 ( .A(n508), .B(n360), .ZN(n427) );
  XOR2_X1 U488 ( .A(G107), .B(G104), .Z(n508) );
  XNOR2_X1 U489 ( .A(n452), .B(KEYINPUT110), .ZN(n666) );
  NAND2_X1 U490 ( .A1(n400), .A2(n662), .ZN(n452) );
  BUF_X1 U491 ( .A(n676), .Z(n409) );
  NOR2_X1 U492 ( .A1(n677), .A2(n389), .ZN(n607) );
  INV_X1 U493 ( .A(KEYINPUT0), .ZN(n385) );
  NAND2_X1 U494 ( .A1(n361), .A2(n579), .ZN(n428) );
  XNOR2_X1 U495 ( .A(n625), .B(n458), .ZN(n626) );
  XNOR2_X1 U496 ( .A(n554), .B(KEYINPUT42), .ZN(n741) );
  AND2_X1 U497 ( .A1(n461), .A2(n582), .ZN(n431) );
  XNOR2_X1 U498 ( .A(n418), .B(KEYINPUT31), .ZN(n654) );
  NOR2_X1 U499 ( .A1(n605), .A2(n682), .ZN(n418) );
  XNOR2_X1 U500 ( .A(n704), .B(n422), .ZN(n706) );
  XNOR2_X1 U501 ( .A(n705), .B(KEYINPUT120), .ZN(n422) );
  XNOR2_X1 U502 ( .A(n703), .B(n702), .ZN(n455) );
  AND2_X1 U503 ( .A1(n516), .A2(n367), .ZN(n354) );
  INV_X1 U504 ( .A(G472), .ZN(n440) );
  XOR2_X1 U505 ( .A(KEYINPUT1), .B(KEYINPUT64), .Z(n355) );
  XOR2_X1 U506 ( .A(G116), .B(n520), .Z(n356) );
  XOR2_X1 U507 ( .A(n502), .B(KEYINPUT25), .Z(n357) );
  XOR2_X1 U508 ( .A(n419), .B(n496), .Z(n358) );
  XNOR2_X1 U509 ( .A(KEYINPUT68), .B(G469), .ZN(n359) );
  XOR2_X1 U510 ( .A(G101), .B(G140), .Z(n360) );
  AND2_X1 U511 ( .A1(n689), .A2(n513), .ZN(n361) );
  AND2_X1 U512 ( .A1(n539), .A2(n648), .ZN(n362) );
  AND2_X1 U513 ( .A1(n607), .A2(n373), .ZN(n363) );
  AND2_X1 U514 ( .A1(n570), .A2(n362), .ZN(n364) );
  AND2_X1 U515 ( .A1(G227), .A2(n728), .ZN(n365) );
  AND2_X1 U516 ( .A1(n434), .A2(n661), .ZN(n366) );
  AND2_X1 U517 ( .A1(n607), .A2(n545), .ZN(n367) );
  AND2_X1 U518 ( .A1(n556), .A2(n354), .ZN(n368) );
  INV_X1 U519 ( .A(n671), .ZN(n424) );
  XOR2_X1 U520 ( .A(G902), .B(KEYINPUT15), .Z(n612) );
  NAND2_X1 U521 ( .A1(n364), .A2(n571), .ZN(n371) );
  XNOR2_X1 U522 ( .A(n499), .B(n498), .ZN(n709) );
  AND2_X1 U523 ( .A1(n400), .A2(n545), .ZN(n373) );
  XNOR2_X2 U524 ( .A(n523), .B(n381), .ZN(n712) );
  NAND2_X1 U525 ( .A1(n644), .A2(n383), .ZN(n596) );
  XNOR2_X1 U526 ( .A(n383), .B(n739), .ZN(G21) );
  XNOR2_X2 U527 ( .A(n384), .B(n385), .ZN(n605) );
  NOR2_X2 U528 ( .A1(n578), .A2(n428), .ZN(n384) );
  XNOR2_X2 U529 ( .A(n387), .B(n386), .ZN(n578) );
  NAND2_X1 U530 ( .A1(n556), .A2(n662), .ZN(n387) );
  INV_X1 U531 ( .A(n551), .ZN(n389) );
  NAND2_X1 U532 ( .A1(n390), .A2(n610), .ZN(n391) );
  NAND2_X1 U533 ( .A1(n391), .A2(KEYINPUT84), .ZN(n393) );
  NAND2_X1 U534 ( .A1(n395), .A2(n392), .ZN(n445) );
  INV_X1 U535 ( .A(KEYINPUT84), .ZN(n397) );
  NOR2_X1 U536 ( .A1(n637), .A2(n399), .ZN(n398) );
  NOR2_X1 U537 ( .A1(n400), .A2(n662), .ZN(n663) );
  INV_X1 U538 ( .A(n614), .ZN(n719) );
  NAND2_X1 U539 ( .A1(n401), .A2(n613), .ZN(n616) );
  XNOR2_X1 U540 ( .A(n402), .B(KEYINPUT82), .ZN(n401) );
  NAND2_X1 U541 ( .A1(n403), .A2(n430), .ZN(n402) );
  NOR2_X1 U542 ( .A1(n614), .A2(n576), .ZN(n403) );
  NAND2_X1 U543 ( .A1(n707), .A2(G210), .ZN(n406) );
  XNOR2_X1 U544 ( .A(n406), .B(n634), .ZN(n635) );
  XNOR2_X1 U545 ( .A(n421), .B(n420), .ZN(n540) );
  NAND2_X1 U546 ( .A1(n407), .A2(n592), .ZN(n593) );
  XNOR2_X1 U547 ( .A(n591), .B(KEYINPUT34), .ZN(n407) );
  NOR2_X1 U548 ( .A1(n446), .A2(n445), .ZN(n611) );
  XNOR2_X1 U549 ( .A(n594), .B(n449), .ZN(n448) );
  AND2_X1 U550 ( .A1(n533), .A2(n411), .ZN(n572) );
  INV_X1 U551 ( .A(n546), .ZN(n412) );
  XNOR2_X1 U552 ( .A(n415), .B(n478), .ZN(n705) );
  XNOR2_X1 U553 ( .A(n484), .B(n356), .ZN(n415) );
  NAND2_X1 U554 ( .A1(n585), .A2(n409), .ZN(n598) );
  NAND2_X1 U555 ( .A1(n439), .A2(n438), .ZN(n437) );
  BUF_X1 U556 ( .A(n588), .Z(n416) );
  XNOR2_X1 U557 ( .A(n727), .B(n433), .ZN(n430) );
  NAND2_X1 U558 ( .A1(n363), .A2(n516), .ZN(n421) );
  INV_X1 U559 ( .A(n598), .ZN(n599) );
  XNOR2_X2 U560 ( .A(n675), .B(KEYINPUT6), .ZN(n601) );
  NAND2_X1 U561 ( .A1(n587), .A2(n416), .ZN(n644) );
  XNOR2_X1 U562 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U563 ( .A(n611), .B(KEYINPUT45), .ZN(n614) );
  NOR2_X2 U564 ( .A1(n605), .A2(n698), .ZN(n591) );
  NOR2_X2 U565 ( .A1(n677), .A2(n676), .ZN(n602) );
  XNOR2_X2 U566 ( .A(n593), .B(KEYINPUT35), .ZN(n738) );
  NAND2_X1 U567 ( .A1(n585), .A2(n431), .ZN(n584) );
  INV_X1 U568 ( .A(n660), .ZN(n434) );
  NAND2_X1 U569 ( .A1(n617), .A2(n440), .ZN(n439) );
  NAND2_X1 U570 ( .A1(n447), .A2(n597), .ZN(n446) );
  NOR2_X2 U571 ( .A1(n612), .A2(n631), .ZN(n530) );
  NAND2_X1 U572 ( .A1(n595), .A2(n448), .ZN(n447) );
  INV_X1 U573 ( .A(KEYINPUT65), .ZN(n449) );
  NOR2_X1 U574 ( .A1(n454), .A2(n711), .ZN(G54) );
  XNOR2_X1 U575 ( .A(n456), .B(n455), .ZN(n454) );
  NAND2_X1 U576 ( .A1(n707), .A2(G469), .ZN(n456) );
  XOR2_X2 U577 ( .A(G113), .B(G104), .Z(n521) );
  AND2_X1 U578 ( .A1(G210), .A2(n486), .ZN(n457) );
  XNOR2_X1 U579 ( .A(KEYINPUT59), .B(KEYINPUT87), .ZN(n458) );
  AND2_X1 U580 ( .A1(G221), .A2(n493), .ZN(n460) );
  XNOR2_X1 U581 ( .A(KEYINPUT104), .B(n581), .ZN(n461) );
  AND2_X1 U582 ( .A1(n567), .A2(n566), .ZN(n568) );
  AND2_X1 U583 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U584 ( .A(KEYINPUT36), .B(KEYINPUT86), .ZN(n534) );
  INV_X1 U585 ( .A(KEYINPUT66), .ZN(n506) );
  XNOR2_X1 U586 ( .A(KEYINPUT33), .B(KEYINPUT71), .ZN(n589) );
  XNOR2_X1 U587 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U588 ( .A(n618), .B(KEYINPUT62), .ZN(n619) );
  XNOR2_X1 U589 ( .A(n460), .B(n494), .ZN(n499) );
  INV_X1 U590 ( .A(KEYINPUT63), .ZN(n622) );
  XNOR2_X1 U591 ( .A(KEYINPUT32), .B(KEYINPUT76), .ZN(n583) );
  XNOR2_X1 U592 ( .A(n622), .B(KEYINPUT88), .ZN(n623) );
  XNOR2_X1 U593 ( .A(n541), .B(KEYINPUT40), .ZN(n740) );
  INV_X1 U594 ( .A(n612), .ZN(n576) );
  XNOR2_X1 U595 ( .A(KEYINPUT13), .B(G475), .ZN(n473) );
  NAND2_X1 U596 ( .A1(G214), .A2(n486), .ZN(n462) );
  XNOR2_X1 U597 ( .A(n463), .B(n462), .ZN(n467) );
  XNOR2_X1 U598 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U599 ( .A(n483), .B(n521), .ZN(n468) );
  XNOR2_X1 U600 ( .A(n469), .B(n468), .ZN(n471) );
  XOR2_X1 U601 ( .A(n494), .B(n471), .Z(n625) );
  NOR2_X1 U602 ( .A1(G902), .A2(n625), .ZN(n472) );
  NAND2_X1 U603 ( .A1(G217), .A2(n493), .ZN(n477) );
  NOR2_X1 U604 ( .A1(G902), .A2(n705), .ZN(n481) );
  NOR2_X1 U605 ( .A1(n537), .A2(n542), .ZN(n482) );
  XOR2_X1 U606 ( .A(KEYINPUT102), .B(n482), .Z(n655) );
  INV_X1 U607 ( .A(KEYINPUT30), .ZN(n492) );
  XNOR2_X2 U608 ( .A(n484), .B(n485), .ZN(n725) );
  XNOR2_X1 U609 ( .A(n488), .B(n487), .ZN(n489) );
  NAND2_X1 U610 ( .A1(G214), .A2(n526), .ZN(n662) );
  NAND2_X1 U611 ( .A1(n586), .A2(n662), .ZN(n491) );
  XNOR2_X1 U612 ( .A(n492), .B(n491), .ZN(n516) );
  XOR2_X1 U613 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n496) );
  XNOR2_X1 U614 ( .A(n358), .B(n497), .ZN(n498) );
  INV_X1 U615 ( .A(G902), .ZN(n500) );
  NAND2_X1 U616 ( .A1(n576), .A2(G234), .ZN(n501) );
  XNOR2_X1 U617 ( .A(n501), .B(KEYINPUT20), .ZN(n503) );
  NAND2_X1 U618 ( .A1(G217), .A2(n503), .ZN(n502) );
  XOR2_X1 U619 ( .A(KEYINPUT93), .B(KEYINPUT21), .Z(n505) );
  NAND2_X1 U620 ( .A1(n503), .A2(G221), .ZN(n504) );
  XNOR2_X1 U621 ( .A(n505), .B(n504), .ZN(n671) );
  NOR2_X1 U622 ( .A1(n588), .A2(n671), .ZN(n507) );
  NAND2_X1 U623 ( .A1(G234), .A2(G237), .ZN(n510) );
  XNOR2_X1 U624 ( .A(n510), .B(KEYINPUT14), .ZN(n689) );
  NOR2_X1 U625 ( .A1(G902), .A2(n728), .ZN(n512) );
  NOR2_X1 U626 ( .A1(G953), .A2(G952), .ZN(n511) );
  NOR2_X1 U627 ( .A1(n512), .A2(n511), .ZN(n513) );
  NAND2_X1 U628 ( .A1(G953), .A2(G900), .ZN(n514) );
  NAND2_X1 U629 ( .A1(n361), .A2(n514), .ZN(n515) );
  XNOR2_X1 U630 ( .A(KEYINPUT79), .B(n515), .ZN(n545) );
  NAND2_X1 U631 ( .A1(G210), .A2(n526), .ZN(n528) );
  INV_X1 U632 ( .A(KEYINPUT91), .ZN(n527) );
  XNOR2_X2 U633 ( .A(n530), .B(n529), .ZN(n556) );
  NOR2_X1 U634 ( .A1(n655), .A2(n540), .ZN(n660) );
  INV_X1 U635 ( .A(n588), .ZN(n531) );
  NAND2_X1 U636 ( .A1(n545), .A2(n662), .ZN(n532) );
  NOR2_X1 U637 ( .A1(n651), .A2(n532), .ZN(n533) );
  NAND2_X1 U638 ( .A1(n572), .A2(n556), .ZN(n535) );
  XNOR2_X1 U639 ( .A(n657), .B(KEYINPUT83), .ZN(n539) );
  INV_X1 U640 ( .A(n556), .ZN(n574) );
  XNOR2_X1 U641 ( .A(KEYINPUT106), .B(n368), .ZN(n538) );
  INV_X1 U642 ( .A(n537), .ZN(n543) );
  NOR2_X1 U643 ( .A1(n542), .A2(n543), .ZN(n592) );
  NAND2_X1 U644 ( .A1(n538), .A2(n592), .ZN(n648) );
  NOR2_X1 U645 ( .A1(n540), .A2(n651), .ZN(n541) );
  NAND2_X1 U646 ( .A1(n543), .A2(n542), .ZN(n665) );
  AND2_X1 U647 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U648 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n548) );
  XNOR2_X1 U649 ( .A(KEYINPUT28), .B(n548), .ZN(n549) );
  XNOR2_X1 U650 ( .A(n550), .B(n549), .ZN(n552) );
  NOR2_X1 U651 ( .A1(n697), .A2(n557), .ZN(n554) );
  XNOR2_X1 U652 ( .A(n555), .B(KEYINPUT46), .ZN(n571) );
  INV_X1 U653 ( .A(n651), .ZN(n558) );
  NOR2_X2 U654 ( .A1(n578), .A2(n557), .ZN(n564) );
  NAND2_X1 U655 ( .A1(n558), .A2(n564), .ZN(n649) );
  INV_X1 U656 ( .A(n655), .ZN(n559) );
  NAND2_X1 U657 ( .A1(n564), .A2(n559), .ZN(n645) );
  NAND2_X1 U658 ( .A1(n649), .A2(n645), .ZN(n561) );
  NOR2_X1 U659 ( .A1(KEYINPUT47), .A2(KEYINPUT73), .ZN(n560) );
  NAND2_X1 U660 ( .A1(n561), .A2(n560), .ZN(n569) );
  NAND2_X1 U661 ( .A1(n655), .A2(n651), .ZN(n608) );
  INV_X1 U662 ( .A(n608), .ZN(n667) );
  NOR2_X1 U663 ( .A1(n667), .A2(KEYINPUT73), .ZN(n562) );
  NAND2_X1 U664 ( .A1(n562), .A2(n564), .ZN(n563) );
  NAND2_X1 U665 ( .A1(n563), .A2(KEYINPUT47), .ZN(n567) );
  AND2_X1 U666 ( .A1(n667), .A2(KEYINPUT73), .ZN(n565) );
  NAND2_X1 U667 ( .A1(n565), .A2(n564), .ZN(n566) );
  NAND2_X1 U668 ( .A1(n409), .A2(n572), .ZN(n573) );
  XNOR2_X1 U669 ( .A(KEYINPUT43), .B(n573), .ZN(n575) );
  NAND2_X1 U670 ( .A1(n575), .A2(n574), .ZN(n661) );
  XNOR2_X1 U671 ( .A(n601), .B(KEYINPUT77), .ZN(n582) );
  INV_X1 U672 ( .A(n665), .ZN(n580) );
  XNOR2_X1 U673 ( .A(n416), .B(KEYINPUT103), .ZN(n672) );
  NOR2_X1 U674 ( .A1(n672), .A2(n409), .ZN(n581) );
  NOR2_X1 U675 ( .A1(n586), .A2(n598), .ZN(n587) );
  XNOR2_X1 U676 ( .A(n596), .B(KEYINPUT85), .ZN(n595) );
  NAND2_X1 U677 ( .A1(n602), .A2(n601), .ZN(n590) );
  XNOR2_X2 U678 ( .A(n590), .B(n589), .ZN(n698) );
  NOR2_X1 U679 ( .A1(n738), .A2(KEYINPUT44), .ZN(n594) );
  NAND2_X1 U680 ( .A1(n596), .A2(KEYINPUT44), .ZN(n597) );
  NAND2_X1 U681 ( .A1(n599), .A2(n672), .ZN(n600) );
  INV_X1 U682 ( .A(n675), .ZN(n604) );
  NAND2_X1 U683 ( .A1(n602), .A2(n604), .ZN(n603) );
  XNOR2_X1 U684 ( .A(n603), .B(KEYINPUT96), .ZN(n682) );
  NOR2_X1 U685 ( .A1(n605), .A2(n604), .ZN(n606) );
  NAND2_X1 U686 ( .A1(n607), .A2(n606), .ZN(n641) );
  NAND2_X1 U687 ( .A1(n654), .A2(n641), .ZN(n609) );
  NAND2_X1 U688 ( .A1(n609), .A2(n608), .ZN(n610) );
  NAND2_X1 U689 ( .A1(KEYINPUT2), .A2(n612), .ZN(n613) );
  NOR2_X1 U690 ( .A1(n614), .A2(n727), .ZN(n693) );
  NAND2_X1 U691 ( .A1(n693), .A2(KEYINPUT2), .ZN(n615) );
  NAND2_X1 U692 ( .A1(n707), .A2(G472), .ZN(n620) );
  XOR2_X1 U693 ( .A(n617), .B(KEYINPUT111), .Z(n618) );
  XNOR2_X1 U694 ( .A(n620), .B(n619), .ZN(n621) );
  NOR2_X2 U695 ( .A1(n621), .A2(n711), .ZN(n624) );
  XNOR2_X1 U696 ( .A(n624), .B(n623), .ZN(G57) );
  NAND2_X1 U697 ( .A1(n707), .A2(G475), .ZN(n627) );
  XNOR2_X1 U698 ( .A(n627), .B(n626), .ZN(n628) );
  NOR2_X2 U699 ( .A1(n628), .A2(n711), .ZN(n630) );
  XOR2_X1 U700 ( .A(KEYINPUT60), .B(KEYINPUT119), .Z(n629) );
  XNOR2_X1 U701 ( .A(n630), .B(n629), .ZN(G60) );
  XOR2_X1 U702 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n633) );
  XNOR2_X1 U703 ( .A(n631), .B(KEYINPUT80), .ZN(n632) );
  NOR2_X2 U704 ( .A1(n635), .A2(n711), .ZN(n636) );
  XNOR2_X1 U705 ( .A(n636), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U706 ( .A(G101), .B(n637), .Z(G3) );
  NOR2_X1 U707 ( .A1(n651), .A2(n641), .ZN(n638) );
  XOR2_X1 U708 ( .A(G104), .B(n638), .Z(G6) );
  XOR2_X1 U709 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n640) );
  XNOR2_X1 U710 ( .A(G107), .B(KEYINPUT112), .ZN(n639) );
  XNOR2_X1 U711 ( .A(n640), .B(n639), .ZN(n643) );
  NOR2_X1 U712 ( .A1(n655), .A2(n641), .ZN(n642) );
  XOR2_X1 U713 ( .A(n643), .B(n642), .Z(G9) );
  XNOR2_X1 U714 ( .A(G110), .B(n644), .ZN(G12) );
  XNOR2_X1 U715 ( .A(KEYINPUT29), .B(KEYINPUT113), .ZN(n646) );
  XNOR2_X1 U716 ( .A(n646), .B(n645), .ZN(n647) );
  XNOR2_X1 U717 ( .A(G128), .B(n647), .ZN(G30) );
  XNOR2_X1 U718 ( .A(G143), .B(n648), .ZN(G45) );
  XNOR2_X1 U719 ( .A(G146), .B(KEYINPUT114), .ZN(n650) );
  XNOR2_X1 U720 ( .A(n650), .B(n649), .ZN(G48) );
  NOR2_X1 U721 ( .A1(n651), .A2(n654), .ZN(n653) );
  XNOR2_X1 U722 ( .A(G113), .B(KEYINPUT115), .ZN(n652) );
  XNOR2_X1 U723 ( .A(n653), .B(n652), .ZN(G15) );
  NOR2_X1 U724 ( .A1(n655), .A2(n654), .ZN(n656) );
  XOR2_X1 U725 ( .A(G116), .B(n656), .Z(G18) );
  XNOR2_X1 U726 ( .A(n657), .B(KEYINPUT116), .ZN(n658) );
  XNOR2_X1 U727 ( .A(n658), .B(KEYINPUT37), .ZN(n659) );
  XNOR2_X1 U728 ( .A(G125), .B(n659), .ZN(G27) );
  XOR2_X1 U729 ( .A(G134), .B(n660), .Z(G36) );
  XNOR2_X1 U730 ( .A(G140), .B(n661), .ZN(G42) );
  XNOR2_X1 U731 ( .A(n663), .B(KEYINPUT118), .ZN(n664) );
  NOR2_X1 U732 ( .A1(n665), .A2(n664), .ZN(n669) );
  NOR2_X1 U733 ( .A1(n667), .A2(n666), .ZN(n668) );
  NOR2_X1 U734 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U735 ( .A1(n670), .A2(n698), .ZN(n687) );
  NOR2_X1 U736 ( .A1(n424), .A2(n672), .ZN(n673) );
  XNOR2_X1 U737 ( .A(n673), .B(KEYINPUT49), .ZN(n674) );
  NAND2_X1 U738 ( .A1(n675), .A2(n674), .ZN(n680) );
  NAND2_X1 U739 ( .A1(n677), .A2(n409), .ZN(n678) );
  XOR2_X1 U740 ( .A(KEYINPUT50), .B(n678), .Z(n679) );
  NOR2_X1 U741 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U742 ( .A(KEYINPUT117), .B(n681), .ZN(n683) );
  NAND2_X1 U743 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U744 ( .A(KEYINPUT51), .B(n684), .ZN(n685) );
  NOR2_X1 U745 ( .A1(n697), .A2(n685), .ZN(n686) );
  NOR2_X1 U746 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U747 ( .A(KEYINPUT52), .B(n688), .ZN(n691) );
  NAND2_X1 U748 ( .A1(G952), .A2(n689), .ZN(n690) );
  NOR2_X1 U749 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U750 ( .A1(G953), .A2(n692), .ZN(n696) );
  NOR2_X1 U751 ( .A1(n693), .A2(KEYINPUT81), .ZN(n694) );
  XOR2_X1 U752 ( .A(KEYINPUT2), .B(n694), .Z(n695) );
  NAND2_X1 U753 ( .A1(n696), .A2(n695), .ZN(n700) );
  NOR2_X1 U754 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U755 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U756 ( .A(KEYINPUT53), .B(n701), .ZN(G75) );
  XOR2_X1 U757 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n702) );
  NAND2_X1 U758 ( .A1(n707), .A2(G478), .ZN(n704) );
  NOR2_X1 U759 ( .A1(n711), .A2(n706), .ZN(G63) );
  NAND2_X1 U760 ( .A1(G217), .A2(n707), .ZN(n708) );
  XNOR2_X1 U761 ( .A(n709), .B(n708), .ZN(n710) );
  NOR2_X1 U762 ( .A1(n711), .A2(n710), .ZN(G66) );
  NOR2_X1 U763 ( .A1(G898), .A2(n728), .ZN(n714) );
  XOR2_X1 U764 ( .A(G110), .B(n712), .Z(n713) );
  NOR2_X1 U765 ( .A1(n714), .A2(n713), .ZN(n715) );
  XOR2_X1 U766 ( .A(KEYINPUT123), .B(n715), .Z(n724) );
  NAND2_X1 U767 ( .A1(G953), .A2(G224), .ZN(n716) );
  XNOR2_X1 U768 ( .A(KEYINPUT61), .B(n716), .ZN(n717) );
  NAND2_X1 U769 ( .A1(n717), .A2(G898), .ZN(n718) );
  XNOR2_X1 U770 ( .A(KEYINPUT121), .B(n718), .ZN(n722) );
  NAND2_X1 U771 ( .A1(n719), .A2(n728), .ZN(n720) );
  XOR2_X1 U772 ( .A(n720), .B(KEYINPUT122), .Z(n721) );
  NOR2_X1 U773 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U774 ( .A(n724), .B(n723), .Z(G69) );
  XNOR2_X1 U775 ( .A(n726), .B(n725), .ZN(n730) );
  XNOR2_X1 U776 ( .A(n727), .B(n730), .ZN(n729) );
  NAND2_X1 U777 ( .A1(n729), .A2(n728), .ZN(n736) );
  XNOR2_X1 U778 ( .A(n730), .B(G227), .ZN(n731) );
  XNOR2_X1 U779 ( .A(n731), .B(KEYINPUT124), .ZN(n732) );
  NAND2_X1 U780 ( .A1(n732), .A2(G900), .ZN(n733) );
  NAND2_X1 U781 ( .A1(G953), .A2(n733), .ZN(n734) );
  XOR2_X1 U782 ( .A(KEYINPUT125), .B(n734), .Z(n735) );
  NAND2_X1 U783 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U784 ( .A(KEYINPUT126), .B(n737), .ZN(G72) );
  XOR2_X1 U785 ( .A(G122), .B(n738), .Z(G24) );
  XOR2_X1 U786 ( .A(G119), .B(KEYINPUT127), .Z(n739) );
  XOR2_X1 U787 ( .A(n740), .B(G131), .Z(G33) );
  XOR2_X1 U788 ( .A(n741), .B(G137), .Z(G39) );
endmodule

