//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 1 1 0 0 1 0 0 0 0 1 1 0 0 1 0 1 0 1 1 0 1 0 1 1 1 1 0 1 1 0 1 1 0 1 1 1 0 0 0 1 0 1 1 1 0 0 0 0 1 0 1 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n847, new_n848, new_n850,
    new_n851, new_n852, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970;
  INV_X1    g000(.A(G141gat), .ZN(new_n202));
  OAI21_X1  g001(.A(KEYINPUT78), .B1(new_n202), .B2(G148gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT78), .ZN(new_n204));
  INV_X1    g003(.A(G148gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n204), .A2(new_n205), .A3(G141gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n202), .A2(G148gat), .ZN(new_n207));
  NAND4_X1  g006(.A1(new_n203), .A2(new_n206), .A3(KEYINPUT79), .A4(new_n207), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n203), .A2(new_n206), .A3(new_n207), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT79), .ZN(new_n210));
  NAND2_X1  g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT2), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AOI22_X1  g013(.A1(new_n209), .A2(new_n210), .B1(new_n211), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n205), .A2(G141gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n207), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT77), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT77), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n207), .A2(new_n216), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n211), .A2(KEYINPUT2), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n218), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT76), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n223), .B1(G155gat), .B2(G162gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n211), .A2(KEYINPUT76), .ZN(new_n225));
  NOR3_X1   g024(.A1(new_n224), .A2(new_n225), .A3(new_n212), .ZN(new_n226));
  AOI22_X1  g025(.A1(new_n208), .A2(new_n215), .B1(new_n222), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT29), .ZN(new_n228));
  XOR2_X1   g027(.A(G211gat), .B(G218gat), .Z(new_n229));
  AND2_X1   g028(.A1(G197gat), .A2(G204gat), .ZN(new_n230));
  NOR2_X1   g029(.A1(G197gat), .A2(G204gat), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  AOI21_X1  g031(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n233));
  OAI21_X1  g032(.A(KEYINPUT73), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(G197gat), .B(G204gat), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT73), .ZN(new_n236));
  INV_X1    g035(.A(new_n233), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n235), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n229), .B1(new_n234), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(G211gat), .A2(G218gat), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT22), .ZN(new_n241));
  INV_X1    g040(.A(G197gat), .ZN(new_n242));
  INV_X1    g041(.A(G204gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(G197gat), .A2(G204gat), .ZN(new_n245));
  AOI221_X4 g044(.A(KEYINPUT73), .B1(new_n240), .B2(new_n241), .C1(new_n244), .C2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n229), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n228), .B1(new_n239), .B2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n227), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n236), .B1(new_n235), .B2(new_n237), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n247), .B1(new_n246), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n238), .A2(new_n229), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n209), .A2(new_n210), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n214), .A2(new_n211), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n256), .A2(new_n208), .A3(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(G141gat), .B(G148gat), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n221), .B1(new_n259), .B2(new_n219), .ZN(new_n260));
  INV_X1    g059(.A(new_n220), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n226), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n258), .A2(new_n262), .A3(new_n250), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n255), .B1(new_n263), .B2(new_n228), .ZN(new_n264));
  OAI21_X1  g063(.A(KEYINPUT83), .B1(new_n251), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(G228gat), .A2(G233gat), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(KEYINPUT84), .B(G22gat), .ZN(new_n269));
  OAI211_X1 g068(.A(KEYINPUT83), .B(new_n266), .C1(new_n251), .C2(new_n264), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n268), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT85), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n268), .A2(KEYINPUT85), .A3(new_n269), .A4(new_n270), .ZN(new_n274));
  INV_X1    g073(.A(new_n269), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n258), .A2(new_n262), .ZN(new_n276));
  AOI21_X1  g075(.A(KEYINPUT29), .B1(new_n253), .B2(new_n254), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n276), .B1(new_n277), .B2(KEYINPUT3), .ZN(new_n278));
  AOI21_X1  g077(.A(KEYINPUT29), .B1(new_n227), .B2(new_n250), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n278), .B1(new_n279), .B2(new_n255), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n266), .B1(new_n280), .B2(KEYINPUT83), .ZN(new_n281));
  INV_X1    g080(.A(new_n270), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n275), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n273), .A2(new_n274), .A3(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(G78gat), .B(G106gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(KEYINPUT31), .B(G50gat), .ZN(new_n286));
  XOR2_X1   g085(.A(new_n285), .B(new_n286), .Z(new_n287));
  NAND2_X1  g086(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n287), .ZN(new_n289));
  AND2_X1   g088(.A1(new_n271), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g089(.A(G22gat), .B1(new_n281), .B2(new_n282), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT34), .ZN(new_n294));
  INV_X1    g093(.A(G120gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(G113gat), .ZN(new_n296));
  INV_X1    g095(.A(G113gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(G120gat), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT68), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n296), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT1), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n295), .A2(KEYINPUT68), .A3(G113gat), .ZN(new_n302));
  AND3_X1   g101(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  NOR2_X1   g102(.A1(G127gat), .A2(G134gat), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(G127gat), .A2(G134gat), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n305), .A2(KEYINPUT69), .A3(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT69), .ZN(new_n308));
  INV_X1    g107(.A(new_n306), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n308), .B1(new_n309), .B2(new_n304), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  AND2_X1   g110(.A1(KEYINPUT67), .A2(G134gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(KEYINPUT67), .A2(G134gat), .ZN(new_n313));
  OAI21_X1  g112(.A(G127gat), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n296), .A2(new_n298), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n304), .B1(new_n315), .B2(new_n301), .ZN(new_n316));
  AOI22_X1  g115(.A1(new_n303), .A2(new_n311), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(G183gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(KEYINPUT27), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT27), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(G183gat), .ZN(new_n321));
  INV_X1    g120(.A(G190gat), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n319), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NOR2_X1   g122(.A1(KEYINPUT65), .A2(KEYINPUT28), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(KEYINPUT27), .B(G183gat), .ZN(new_n326));
  INV_X1    g125(.A(new_n324), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n326), .A2(new_n322), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(G169gat), .A2(G176gat), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT26), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  OAI211_X1 g131(.A(new_n332), .B(KEYINPUT66), .C1(G169gat), .C2(G176gat), .ZN(new_n333));
  NOR2_X1   g132(.A1(G169gat), .A2(G176gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(new_n331), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT66), .ZN(new_n336));
  AOI21_X1  g135(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n336), .B1(new_n337), .B2(new_n334), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n333), .A2(new_n335), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(G183gat), .A2(G190gat), .ZN(new_n340));
  AND3_X1   g139(.A1(new_n329), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT24), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n318), .A2(new_n322), .ZN(new_n344));
  NAND3_X1  g143(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(G169gat), .ZN(new_n347));
  INV_X1    g146(.A(G176gat), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n347), .A2(new_n348), .A3(KEYINPUT23), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT23), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n350), .B1(G169gat), .B2(G176gat), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n346), .A2(new_n349), .A3(new_n330), .A4(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT25), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n340), .A2(KEYINPUT64), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT64), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n355), .A2(G183gat), .A3(G190gat), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n354), .A2(new_n356), .A3(new_n342), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n357), .A2(new_n344), .A3(new_n345), .ZN(new_n358));
  AND4_X1   g157(.A1(KEYINPUT25), .A2(new_n349), .A3(new_n351), .A4(new_n330), .ZN(new_n359));
  AOI22_X1  g158(.A1(new_n352), .A2(new_n353), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n317), .B1(new_n341), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n358), .A2(new_n359), .ZN(new_n362));
  INV_X1    g161(.A(new_n346), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n349), .A2(new_n351), .A3(new_n330), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n353), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n316), .A2(new_n314), .ZN(new_n367));
  INV_X1    g166(.A(new_n311), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n301), .B(new_n302), .C1(new_n315), .C2(KEYINPUT68), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n367), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n329), .A2(new_n339), .A3(new_n340), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n366), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n361), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(G227gat), .ZN(new_n374));
  INV_X1    g173(.A(G233gat), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n294), .B1(new_n373), .B2(new_n377), .ZN(new_n378));
  AOI211_X1 g177(.A(KEYINPUT34), .B(new_n376), .C1(new_n361), .C2(new_n372), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT32), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n361), .A2(new_n376), .A3(new_n372), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(KEYINPUT70), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT70), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n361), .A2(new_n385), .A3(new_n372), .A4(new_n376), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n382), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT33), .B1(new_n384), .B2(new_n386), .ZN(new_n388));
  XNOR2_X1  g187(.A(KEYINPUT71), .B(G71gat), .ZN(new_n389));
  INV_X1    g188(.A(G99gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n389), .B(new_n390), .ZN(new_n391));
  XOR2_X1   g190(.A(G15gat), .B(G43gat), .Z(new_n392));
  XOR2_X1   g191(.A(new_n391), .B(new_n392), .Z(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NOR3_X1   g193(.A1(new_n387), .A2(new_n388), .A3(new_n394), .ZN(new_n395));
  AOI221_X4 g194(.A(new_n382), .B1(KEYINPUT33), .B2(new_n393), .C1(new_n384), .C2(new_n386), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n381), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(KEYINPUT72), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n384), .A2(new_n386), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(KEYINPUT32), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT33), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n400), .A2(new_n402), .A3(new_n393), .ZN(new_n403));
  INV_X1    g202(.A(new_n396), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n380), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT72), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n403), .A2(new_n404), .A3(new_n380), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n293), .A2(new_n398), .A3(new_n407), .A4(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n255), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT29), .B1(new_n366), .B2(new_n371), .ZN(new_n411));
  NAND2_X1  g210(.A1(G226gat), .A2(G233gat), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n412), .B1(new_n366), .B2(new_n371), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n410), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  XOR2_X1   g215(.A(G8gat), .B(G36gat), .Z(new_n417));
  XNOR2_X1  g216(.A(new_n417), .B(KEYINPUT74), .ZN(new_n418));
  XNOR2_X1  g217(.A(G64gat), .B(G92gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n418), .B(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n415), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n421), .B(new_n255), .C1(new_n413), .C2(new_n411), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n416), .A2(new_n420), .A3(new_n422), .ZN(new_n423));
  AND2_X1   g222(.A1(new_n423), .A2(KEYINPUT30), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n423), .A2(KEYINPUT30), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n416), .A2(new_n422), .ZN(new_n426));
  INV_X1    g225(.A(new_n420), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT75), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT75), .ZN(new_n429));
  AOI211_X1 g228(.A(new_n429), .B(new_n420), .C1(new_n416), .C2(new_n422), .ZN(new_n430));
  OAI22_X1  g229(.A1(new_n424), .A2(new_n425), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(G1gat), .B(G29gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n433), .B(KEYINPUT0), .ZN(new_n434));
  XNOR2_X1  g233(.A(G57gat), .B(G85gat), .ZN(new_n435));
  XOR2_X1   g234(.A(new_n434), .B(new_n435), .Z(new_n436));
  NAND2_X1  g235(.A1(new_n276), .A2(KEYINPUT3), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n437), .A2(new_n263), .A3(new_n370), .ZN(new_n438));
  NAND2_X1  g237(.A1(G225gat), .A2(G233gat), .ZN(new_n439));
  AND2_X1   g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  XOR2_X1   g239(.A(KEYINPUT80), .B(KEYINPUT5), .Z(new_n441));
  NAND3_X1  g240(.A1(new_n317), .A2(new_n262), .A3(new_n258), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n442), .A2(KEYINPUT82), .A3(KEYINPUT4), .ZN(new_n443));
  OAI21_X1  g242(.A(KEYINPUT4), .B1(new_n276), .B2(new_n370), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT4), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n227), .A2(new_n445), .A3(new_n317), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT82), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n444), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n440), .A2(new_n441), .A3(new_n443), .A4(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n444), .A2(new_n446), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n450), .A2(new_n439), .A3(new_n438), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n276), .A2(new_n370), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(new_n442), .ZN(new_n453));
  INV_X1    g252(.A(new_n439), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n441), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n451), .A2(KEYINPUT81), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(KEYINPUT81), .B1(new_n451), .B2(new_n455), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n436), .B(new_n449), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT6), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n451), .A2(new_n455), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT81), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n451), .A2(KEYINPUT81), .A3(new_n455), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n436), .B1(new_n465), .B2(new_n449), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n460), .A2(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n449), .B1(new_n456), .B2(new_n457), .ZN(new_n468));
  INV_X1    g267(.A(new_n436), .ZN(new_n469));
  AND3_X1   g268(.A1(new_n468), .A2(KEYINPUT6), .A3(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n432), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT35), .B1(new_n409), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n460), .A2(new_n466), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n468), .A2(new_n469), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n474), .A2(new_n459), .A3(new_n458), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n431), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  AOI22_X1  g275(.A1(new_n284), .A2(new_n287), .B1(new_n291), .B2(new_n290), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n477), .A2(KEYINPUT35), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n397), .A2(new_n408), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT86), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n397), .A2(KEYINPUT86), .A3(new_n408), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n476), .A2(new_n478), .A3(new_n481), .A4(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n472), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n471), .A2(new_n477), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n420), .B1(new_n426), .B2(KEYINPUT37), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT38), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT37), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n416), .A2(new_n488), .A3(new_n422), .ZN(new_n489));
  AND3_X1   g288(.A1(new_n486), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  AOI22_X1  g289(.A1(new_n486), .A2(new_n489), .B1(new_n487), .B2(new_n423), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n492), .A2(new_n473), .A3(new_n475), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT40), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n448), .A2(new_n438), .A3(new_n443), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(new_n454), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n453), .A2(new_n454), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT39), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AND2_X1   g298(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n495), .A2(new_n498), .A3(new_n454), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(new_n436), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n494), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n496), .A2(new_n499), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n504), .A2(KEYINPUT40), .A3(new_n436), .A4(new_n501), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n431), .A2(new_n474), .A3(new_n503), .A4(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n493), .A2(new_n293), .A3(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n408), .B1(new_n405), .B2(new_n406), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n397), .A2(KEYINPUT72), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT36), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  OR2_X1    g309(.A1(new_n479), .A2(KEYINPUT36), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n485), .A2(new_n507), .A3(new_n510), .A4(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n484), .A2(new_n512), .ZN(new_n513));
  XOR2_X1   g312(.A(G43gat), .B(G50gat), .Z(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT88), .ZN(new_n515));
  XNOR2_X1  g314(.A(G43gat), .B(G50gat), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT88), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n515), .A2(KEYINPUT15), .A3(new_n518), .ZN(new_n519));
  NOR2_X1   g318(.A1(G29gat), .A2(G36gat), .ZN(new_n520));
  XOR2_X1   g319(.A(new_n520), .B(KEYINPUT14), .Z(new_n521));
  NOR2_X1   g320(.A1(new_n521), .A2(KEYINPUT89), .ZN(new_n522));
  XNOR2_X1  g321(.A(KEYINPUT90), .B(G36gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(G29gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n520), .B(KEYINPUT14), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT89), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n519), .B1(new_n522), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n515), .A2(KEYINPUT15), .A3(new_n518), .ZN(new_n529));
  OR2_X1    g328(.A1(new_n516), .A2(KEYINPUT15), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n529), .A2(new_n521), .A3(new_n524), .A4(new_n530), .ZN(new_n531));
  AND2_X1   g330(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n532), .A2(KEYINPUT91), .ZN(new_n533));
  AND3_X1   g332(.A1(new_n528), .A2(KEYINPUT91), .A3(new_n531), .ZN(new_n534));
  OR2_X1    g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT17), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(G1gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT16), .ZN(new_n539));
  XOR2_X1   g338(.A(G15gat), .B(G22gat), .Z(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(KEYINPUT92), .ZN(new_n541));
  MUX2_X1   g340(.A(new_n539), .B(new_n538), .S(new_n541), .Z(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(G8gat), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n532), .A2(KEYINPUT17), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n537), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(G229gat), .A2(G233gat), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT93), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n535), .A2(new_n543), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n548), .B1(new_n535), .B2(new_n543), .ZN(new_n551));
  OAI211_X1 g350(.A(new_n546), .B(new_n547), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT18), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n551), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(new_n549), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n556), .A2(KEYINPUT18), .A3(new_n547), .A4(new_n546), .ZN(new_n557));
  OAI22_X1  g356(.A1(new_n550), .A2(new_n551), .B1(new_n535), .B2(new_n543), .ZN(new_n558));
  XOR2_X1   g357(.A(new_n547), .B(KEYINPUT13), .Z(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n554), .A2(new_n557), .A3(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(G113gat), .B(G141gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(KEYINPUT87), .B(G197gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  XOR2_X1   g363(.A(KEYINPUT11), .B(G169gat), .Z(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(KEYINPUT12), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n561), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n554), .A2(new_n557), .A3(new_n560), .A4(new_n567), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AND3_X1   g370(.A1(new_n513), .A2(KEYINPUT94), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(KEYINPUT94), .B1(new_n513), .B2(new_n571), .ZN(new_n573));
  OR2_X1    g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n575));
  XOR2_X1   g374(.A(new_n575), .B(KEYINPUT97), .Z(new_n576));
  XNOR2_X1  g375(.A(G134gat), .B(G162gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(G85gat), .A2(G92gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(KEYINPUT7), .ZN(new_n581));
  NAND2_X1  g380(.A1(G99gat), .A2(G106gat), .ZN(new_n582));
  INV_X1    g381(.A(G85gat), .ZN(new_n583));
  INV_X1    g382(.A(G92gat), .ZN(new_n584));
  AOI22_X1  g383(.A1(KEYINPUT8), .A2(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(G99gat), .B(G106gat), .ZN(new_n587));
  XOR2_X1   g386(.A(new_n586), .B(new_n587), .Z(new_n588));
  NAND3_X1  g387(.A1(new_n537), .A2(new_n545), .A3(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n588), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n535), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n592));
  AOI21_X1  g391(.A(KEYINPUT98), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT98), .ZN(new_n594));
  INV_X1    g393(.A(new_n592), .ZN(new_n595));
  AOI211_X1 g394(.A(new_n594), .B(new_n595), .C1(new_n535), .C2(new_n590), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n589), .B1(new_n593), .B2(new_n596), .ZN(new_n597));
  XOR2_X1   g396(.A(G190gat), .B(G218gat), .Z(new_n598));
  AND2_X1   g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n597), .A2(new_n598), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n579), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  OR2_X1    g400(.A1(new_n597), .A2(new_n598), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n597), .A2(new_n598), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n602), .A2(new_n578), .A3(new_n603), .ZN(new_n604));
  AND2_X1   g403(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  XOR2_X1   g404(.A(G57gat), .B(G64gat), .Z(new_n606));
  INV_X1    g405(.A(KEYINPUT9), .ZN(new_n607));
  INV_X1    g406(.A(G71gat), .ZN(new_n608));
  INV_X1    g407(.A(G78gat), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g410(.A(G71gat), .B(G78gat), .Z(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT21), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(G231gat), .A2(G233gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(G127gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n613), .A2(new_n614), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n543), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n619), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(KEYINPUT95), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(G155gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(G183gat), .B(G211gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT96), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n625), .B(new_n627), .ZN(new_n628));
  XOR2_X1   g427(.A(new_n622), .B(new_n628), .Z(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  OR2_X1    g429(.A1(new_n588), .A2(new_n613), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n588), .A2(new_n613), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(G230gat), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n634), .A2(new_n375), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n636), .B(KEYINPUT99), .Z(new_n637));
  INV_X1    g436(.A(KEYINPUT10), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n631), .A2(new_n638), .A3(new_n632), .ZN(new_n639));
  OR3_X1    g438(.A1(new_n588), .A2(new_n613), .A3(new_n638), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n635), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n637), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g442(.A(G120gat), .B(G148gat), .Z(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(KEYINPUT100), .ZN(new_n645));
  XNOR2_X1  g444(.A(G176gat), .B(G204gat), .ZN(new_n646));
  XOR2_X1   g445(.A(new_n645), .B(new_n646), .Z(new_n647));
  NAND2_X1  g446(.A1(new_n643), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n647), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n637), .A2(new_n649), .A3(new_n642), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n605), .A2(new_n630), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n574), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n467), .A2(new_n470), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(new_n538), .ZN(G1324gat));
  INV_X1    g458(.A(G8gat), .ZN(new_n660));
  INV_X1    g459(.A(new_n655), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n660), .B1(new_n661), .B2(new_n431), .ZN(new_n662));
  XNOR2_X1  g461(.A(KEYINPUT101), .B(KEYINPUT16), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(G8gat), .ZN(new_n664));
  NOR3_X1   g463(.A1(new_n655), .A2(new_n432), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(KEYINPUT42), .B1(new_n662), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n666), .B1(KEYINPUT42), .B2(new_n665), .ZN(G1325gat));
  AND2_X1   g466(.A1(new_n510), .A2(new_n511), .ZN(new_n668));
  OAI21_X1  g467(.A(G15gat), .B1(new_n655), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n481), .A2(new_n482), .ZN(new_n670));
  OR2_X1    g469(.A1(new_n670), .A2(G15gat), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n669), .B1(new_n655), .B2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT102), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n672), .B(new_n673), .ZN(G1326gat));
  NOR2_X1   g473(.A1(new_n655), .A2(new_n293), .ZN(new_n675));
  XOR2_X1   g474(.A(KEYINPUT43), .B(G22gat), .Z(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(G1327gat));
  NAND2_X1  g476(.A1(new_n629), .A2(new_n652), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n605), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n574), .A2(new_n679), .ZN(new_n680));
  OR3_X1    g479(.A1(new_n680), .A2(G29gat), .A3(new_n657), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT45), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n684));
  AND2_X1   g483(.A1(new_n293), .A2(new_n506), .ZN(new_n685));
  AOI22_X1  g484(.A1(new_n685), .A2(new_n493), .B1(new_n471), .B2(new_n477), .ZN(new_n686));
  AOI22_X1  g485(.A1(new_n668), .A2(new_n686), .B1(new_n472), .B2(new_n483), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n684), .B1(new_n687), .B2(new_n605), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n601), .A2(new_n604), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n513), .A2(KEYINPUT44), .A3(new_n689), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n571), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n692), .A2(new_n678), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(G29gat), .B1(new_n694), .B2(new_n657), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n681), .A2(new_n682), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n683), .A2(new_n695), .A3(new_n696), .ZN(G1328gat));
  NOR3_X1   g496(.A1(new_n680), .A2(new_n432), .A3(new_n523), .ZN(new_n698));
  XOR2_X1   g497(.A(KEYINPUT103), .B(KEYINPUT46), .Z(new_n699));
  OR2_X1    g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n523), .B1(new_n694), .B2(new_n432), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n698), .A2(new_n699), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n700), .A2(new_n701), .A3(new_n702), .ZN(G1329gat));
  NOR2_X1   g502(.A1(new_n680), .A2(new_n670), .ZN(new_n704));
  INV_X1    g503(.A(new_n668), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(G43gat), .ZN(new_n706));
  OAI22_X1  g505(.A1(new_n704), .A2(G43gat), .B1(new_n694), .B2(new_n706), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g507(.A1(new_n293), .A2(G50gat), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n574), .A2(new_n679), .A3(new_n709), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n688), .A2(new_n690), .A3(new_n477), .A4(new_n693), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(G50gat), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n710), .A2(KEYINPUT48), .A3(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT105), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n711), .A2(KEYINPUT105), .A3(G50gat), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n715), .A2(new_n710), .A3(new_n716), .ZN(new_n717));
  XOR2_X1   g516(.A(KEYINPUT104), .B(KEYINPUT48), .Z(new_n718));
  AND3_X1   g517(.A1(new_n717), .A2(KEYINPUT106), .A3(new_n718), .ZN(new_n719));
  AOI21_X1  g518(.A(KEYINPUT106), .B1(new_n717), .B2(new_n718), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n713), .B1(new_n719), .B2(new_n720), .ZN(G1331gat));
  NOR4_X1   g520(.A1(new_n689), .A2(new_n571), .A3(new_n629), .A4(new_n652), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n513), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n656), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g525(.A1(new_n724), .A2(KEYINPUT107), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT107), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n723), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n730), .A2(new_n432), .ZN(new_n731));
  NOR2_X1   g530(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n732));
  AND2_X1   g531(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n731), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n734), .B1(new_n731), .B2(new_n732), .ZN(G1333gat));
  NAND4_X1  g534(.A1(new_n727), .A2(G71gat), .A3(new_n705), .A4(new_n729), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n608), .B1(new_n723), .B2(new_n670), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT50), .ZN(G1334gat));
  XNOR2_X1  g538(.A(KEYINPUT108), .B(G78gat), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(KEYINPUT109), .B1(new_n730), .B2(new_n293), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n730), .A2(KEYINPUT109), .A3(new_n293), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n741), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n744), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n746), .A2(new_n742), .A3(new_n740), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(G1335gat));
  NOR2_X1   g547(.A1(new_n571), .A2(new_n630), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n513), .A2(new_n689), .A3(new_n749), .ZN(new_n750));
  XOR2_X1   g549(.A(new_n750), .B(KEYINPUT51), .Z(new_n751));
  AND2_X1   g550(.A1(new_n751), .A2(new_n651), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n752), .A2(new_n583), .A3(new_n656), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n569), .A2(new_n629), .A3(new_n570), .A4(new_n651), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(KEYINPUT110), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n688), .A2(new_n690), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(KEYINPUT111), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT111), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n688), .A2(new_n690), .A3(new_n755), .A4(new_n758), .ZN(new_n759));
  AND3_X1   g558(.A1(new_n757), .A2(new_n656), .A3(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n753), .B1(new_n583), .B2(new_n760), .ZN(G1336gat));
  NAND3_X1  g560(.A1(new_n691), .A2(new_n431), .A3(new_n755), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT113), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n584), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n764), .B1(new_n763), .B2(new_n762), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n652), .A2(G92gat), .A3(new_n432), .ZN(new_n766));
  AOI21_X1  g565(.A(KEYINPUT52), .B1(new_n751), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT52), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n757), .A2(new_n431), .A3(new_n759), .ZN(new_n770));
  AND3_X1   g569(.A1(new_n750), .A2(KEYINPUT112), .A3(KEYINPUT51), .ZN(new_n771));
  AOI21_X1  g570(.A(KEYINPUT51), .B1(new_n750), .B2(KEYINPUT112), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI22_X1  g572(.A1(new_n770), .A2(G92gat), .B1(new_n773), .B2(new_n766), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n768), .B1(new_n769), .B2(new_n774), .ZN(G1337gat));
  NAND4_X1  g574(.A1(new_n752), .A2(new_n390), .A3(new_n482), .A4(new_n481), .ZN(new_n776));
  AND3_X1   g575(.A1(new_n757), .A2(new_n705), .A3(new_n759), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n776), .B1(new_n390), .B2(new_n777), .ZN(G1338gat));
  NOR3_X1   g577(.A1(new_n652), .A2(G106gat), .A3(new_n293), .ZN(new_n779));
  AOI21_X1  g578(.A(KEYINPUT53), .B1(new_n751), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n691), .A2(new_n477), .A3(new_n755), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(KEYINPUT115), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(G106gat), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n781), .A2(KEYINPUT115), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n780), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n757), .A2(new_n477), .A3(new_n759), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(G106gat), .ZN(new_n787));
  INV_X1    g586(.A(new_n779), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n771), .A2(new_n772), .A3(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(KEYINPUT114), .B1(new_n791), .B2(KEYINPUT53), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n789), .B1(new_n786), .B2(G106gat), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT114), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT53), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n785), .B1(new_n792), .B2(new_n796), .ZN(G1339gat));
  NAND2_X1  g596(.A1(new_n656), .A2(new_n432), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n798), .A2(new_n670), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n639), .A2(new_n635), .A3(new_n640), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n642), .A2(KEYINPUT54), .A3(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT54), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n649), .B1(new_n641), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n801), .A2(KEYINPUT55), .A3(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(KEYINPUT55), .B1(new_n801), .B2(new_n803), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n805), .A2(KEYINPUT116), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT116), .ZN(new_n807));
  AOI211_X1 g606(.A(new_n807), .B(KEYINPUT55), .C1(new_n801), .C2(new_n803), .ZN(new_n808));
  OAI211_X1 g607(.A(new_n650), .B(new_n804), .C1(new_n806), .C2(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n809), .B1(new_n569), .B2(new_n570), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n558), .A2(new_n559), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n547), .B1(new_n556), .B2(new_n546), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n566), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n813), .A2(new_n570), .A3(new_n651), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(KEYINPUT117), .B1(new_n810), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n806), .A2(new_n808), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n650), .A2(new_n804), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n570), .ZN(new_n820));
  AOI22_X1  g619(.A1(new_n552), .A2(new_n553), .B1(new_n558), .B2(new_n559), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n567), .B1(new_n821), .B2(new_n557), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n819), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT117), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n823), .A2(new_n824), .A3(new_n814), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n816), .A2(new_n825), .A3(new_n605), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n689), .A2(new_n570), .A3(new_n813), .A4(new_n819), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n630), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n653), .A2(new_n571), .ZN(new_n829));
  OAI211_X1 g628(.A(new_n293), .B(new_n799), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(G113gat), .B1(new_n830), .B2(new_n692), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n826), .A2(new_n827), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(new_n629), .ZN(new_n833));
  INV_X1    g632(.A(new_n829), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n657), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n409), .A2(new_n431), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n571), .A2(new_n297), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n831), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(KEYINPUT118), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT118), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n831), .B(new_n841), .C1(new_n837), .C2(new_n838), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n840), .A2(new_n842), .ZN(G1340gat));
  NOR3_X1   g642(.A1(new_n830), .A2(new_n295), .A3(new_n652), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n835), .A2(new_n651), .A3(new_n836), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n844), .B1(new_n845), .B2(new_n295), .ZN(G1341gat));
  OAI21_X1  g645(.A(G127gat), .B1(new_n830), .B2(new_n629), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n630), .A2(new_n618), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n847), .B1(new_n837), .B2(new_n848), .ZN(G1342gat));
  OR3_X1    g648(.A1(new_n605), .A2(new_n313), .A3(new_n312), .ZN(new_n850));
  OR3_X1    g649(.A1(new_n837), .A2(KEYINPUT56), .A3(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(G134gat), .B1(new_n830), .B2(new_n605), .ZN(new_n852));
  OAI21_X1  g651(.A(KEYINPUT56), .B1(new_n837), .B2(new_n850), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(G1343gat));
  NAND3_X1  g653(.A1(new_n668), .A2(new_n656), .A3(new_n432), .ZN(new_n855));
  OR2_X1    g654(.A1(new_n818), .A2(new_n805), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n856), .B1(new_n569), .B2(new_n570), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n605), .B1(new_n857), .B2(new_n815), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n630), .B1(new_n858), .B2(new_n827), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n477), .B1(new_n859), .B2(new_n829), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n855), .B1(new_n860), .B2(KEYINPUT57), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n293), .A2(KEYINPUT57), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n862), .B1(new_n828), .B2(new_n829), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n861), .A2(new_n863), .A3(new_n571), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(G141gat), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n705), .A2(new_n293), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n867), .A2(new_n431), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n835), .A2(new_n202), .A3(new_n571), .A4(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n865), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(KEYINPUT58), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT58), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n865), .A2(new_n869), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n871), .A2(new_n873), .ZN(G1344gat));
  NAND2_X1  g673(.A1(new_n205), .A2(KEYINPUT59), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n833), .A2(new_n834), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n876), .A2(new_n656), .A3(new_n868), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n875), .B1(new_n878), .B2(new_n651), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT59), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n861), .A2(new_n863), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n880), .B1(new_n881), .B2(new_n652), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT57), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n293), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n884), .B1(new_n828), .B2(new_n829), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n860), .A2(new_n883), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT119), .ZN(new_n888));
  OR2_X1    g687(.A1(new_n855), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n855), .A2(new_n888), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n652), .A2(new_n880), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n887), .A2(new_n889), .A3(new_n890), .A4(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n882), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n879), .B1(new_n893), .B2(G148gat), .ZN(G1345gat));
  INV_X1    g693(.A(G155gat), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n881), .A2(new_n895), .A3(new_n629), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n877), .A2(new_n629), .ZN(new_n897));
  AOI21_X1  g696(.A(G155gat), .B1(new_n897), .B2(KEYINPUT120), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT120), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n899), .B1(new_n877), .B2(new_n629), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n896), .B1(new_n898), .B2(new_n900), .ZN(G1346gat));
  OR3_X1    g700(.A1(new_n877), .A2(G162gat), .A3(new_n605), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT121), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n903), .B1(new_n881), .B2(new_n605), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(G162gat), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n881), .A2(new_n903), .A3(new_n605), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n902), .B1(new_n905), .B2(new_n906), .ZN(G1347gat));
  NAND2_X1  g706(.A1(new_n657), .A2(new_n431), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(KEYINPUT122), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n909), .A2(new_n670), .ZN(new_n910));
  OAI211_X1 g709(.A(new_n293), .B(new_n910), .C1(new_n828), .C2(new_n829), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n911), .A2(new_n347), .A3(new_n692), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n409), .A2(new_n432), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n876), .A2(new_n657), .A3(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(new_n571), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n912), .B1(new_n916), .B2(new_n347), .ZN(G1348gat));
  OAI21_X1  g716(.A(G176gat), .B1(new_n911), .B2(new_n652), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n651), .A2(new_n348), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n918), .B1(new_n914), .B2(new_n919), .ZN(G1349gat));
  INV_X1    g719(.A(KEYINPUT123), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n921), .A2(KEYINPUT60), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n921), .A2(KEYINPUT60), .ZN(new_n923));
  OAI21_X1  g722(.A(G183gat), .B1(new_n911), .B2(new_n629), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n630), .A2(new_n326), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n876), .A2(new_n657), .A3(new_n913), .A4(new_n925), .ZN(new_n926));
  AOI211_X1 g725(.A(new_n922), .B(new_n923), .C1(new_n924), .C2(new_n926), .ZN(new_n927));
  AND4_X1   g726(.A1(new_n921), .A2(new_n924), .A3(KEYINPUT60), .A4(new_n926), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n927), .A2(new_n928), .ZN(G1350gat));
  OAI21_X1  g728(.A(G190gat), .B1(new_n911), .B2(new_n605), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT61), .ZN(new_n931));
  OR2_X1    g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n930), .A2(new_n931), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n605), .A2(G190gat), .ZN(new_n934));
  AOI21_X1  g733(.A(KEYINPUT124), .B1(new_n915), .B2(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT124), .ZN(new_n936));
  NOR4_X1   g735(.A1(new_n914), .A2(new_n936), .A3(G190gat), .A4(new_n605), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n932), .B(new_n933), .C1(new_n935), .C2(new_n937), .ZN(G1351gat));
  NOR2_X1   g737(.A1(new_n867), .A2(new_n432), .ZN(new_n939));
  OAI211_X1 g738(.A(new_n657), .B(new_n939), .C1(new_n828), .C2(new_n829), .ZN(new_n940));
  INV_X1    g739(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(G197gat), .B1(new_n941), .B2(new_n571), .ZN(new_n942));
  OR2_X1    g741(.A1(new_n909), .A2(new_n705), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n943), .B1(new_n885), .B2(new_n886), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n692), .A2(new_n242), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n942), .B1(new_n944), .B2(new_n945), .ZN(G1352gat));
  INV_X1    g745(.A(new_n944), .ZN(new_n947));
  OAI21_X1  g746(.A(G204gat), .B1(new_n947), .B2(new_n652), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n940), .A2(G204gat), .A3(new_n652), .ZN(new_n949));
  XOR2_X1   g748(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n950));
  OR2_X1    g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n949), .A2(new_n950), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n948), .A2(new_n951), .A3(new_n952), .ZN(G1353gat));
  INV_X1    g752(.A(G211gat), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n941), .A2(new_n954), .A3(new_n630), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT63), .ZN(new_n956));
  AOI211_X1 g755(.A(new_n956), .B(new_n954), .C1(new_n944), .C2(new_n630), .ZN(new_n957));
  INV_X1    g756(.A(new_n943), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n887), .A2(new_n630), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g758(.A(KEYINPUT63), .B1(new_n959), .B2(G211gat), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n955), .B1(new_n957), .B2(new_n960), .ZN(G1354gat));
  NAND2_X1  g760(.A1(new_n947), .A2(KEYINPUT127), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n689), .A2(G218gat), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT127), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n963), .B1(new_n944), .B2(new_n964), .ZN(new_n965));
  INV_X1    g764(.A(G218gat), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n966), .B1(new_n940), .B2(new_n605), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT126), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI211_X1 g768(.A(KEYINPUT126), .B(new_n966), .C1(new_n940), .C2(new_n605), .ZN(new_n970));
  AOI22_X1  g769(.A1(new_n962), .A2(new_n965), .B1(new_n969), .B2(new_n970), .ZN(G1355gat));
endmodule


