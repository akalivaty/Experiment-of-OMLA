//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 1 1 1 0 1 0 1 1 0 0 0 1 0 0 0 0 1 1 1 1 1 0 0 1 1 0 0 1 0 0 0 0 0 0 1 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:00 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1276, new_n1277, new_n1278, new_n1279;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR3_X1   g0007(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT0), .Z(new_n210));
  AOI22_X1  g0010(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n211));
  INV_X1    g0011(.A(G116), .ZN(new_n212));
  INV_X1    g0012(.A(G270), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n215));
  INV_X1    g0015(.A(G50), .ZN(new_n216));
  INV_X1    g0016(.A(G226), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI211_X1 g0020(.A(new_n214), .B(new_n220), .C1(G97), .C2(G257), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n221), .B1(G1), .B2(G20), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT1), .Z(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n224), .A2(new_n207), .ZN(new_n225));
  OAI21_X1  g0025(.A(G50), .B1(G58), .B2(G68), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  AOI211_X1 g0027(.A(new_n210), .B(new_n223), .C1(new_n225), .C2(new_n227), .ZN(G361));
  XNOR2_X1  g0028(.A(G250), .B(G257), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(new_n213), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT65), .B(G264), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G226), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G238), .B(G244), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n233), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G68), .B(G77), .Z(new_n240));
  XNOR2_X1  g0040(.A(G50), .B(G58), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(new_n224), .ZN(new_n248));
  AOI21_X1  g0048(.A(new_n248), .B1(new_n206), .B2(G20), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n250), .A2(new_n216), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n253));
  NOR2_X1   g0053(.A1(G58), .A2(G68), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n207), .B1(new_n254), .B2(new_n216), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G20), .A2(G33), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G150), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AND2_X1   g0059(.A1(KEYINPUT69), .A2(KEYINPUT8), .ZN(new_n260));
  NOR2_X1   g0060(.A1(KEYINPUT69), .A2(KEYINPUT8), .ZN(new_n261));
  OAI21_X1  g0061(.A(G58), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT70), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G58), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(KEYINPUT8), .ZN(new_n266));
  OR2_X1    g0066(.A1(new_n266), .A2(KEYINPUT68), .ZN(new_n267));
  OAI211_X1 g0067(.A(KEYINPUT70), .B(G58), .C1(new_n260), .C2(new_n261), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n266), .A2(KEYINPUT68), .ZN(new_n269));
  NAND4_X1  g0069(.A1(new_n264), .A2(new_n267), .A3(new_n268), .A4(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G33), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n271), .A2(G20), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(KEYINPUT71), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n207), .A2(G33), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT71), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  AOI211_X1 g0077(.A(new_n255), .B(new_n259), .C1(new_n270), .C2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n248), .ZN(new_n279));
  OAI221_X1 g0079(.A(new_n252), .B1(G50), .B2(new_n253), .C1(new_n278), .C2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT9), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT67), .ZN(new_n283));
  NAND2_X1  g0083(.A1(G33), .A2(G41), .ZN(new_n284));
  AND4_X1   g0084(.A1(new_n283), .A2(new_n284), .A3(G1), .A4(G13), .ZN(new_n285));
  AND2_X1   g0085(.A1(G1), .A2(G13), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n283), .B1(new_n286), .B2(new_n284), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  XNOR2_X1  g0088(.A(KEYINPUT3), .B(G33), .ZN(new_n289));
  INV_X1    g0089(.A(G1698), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G222), .ZN(new_n291));
  XNOR2_X1  g0091(.A(KEYINPUT66), .B(G223), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n289), .B(new_n291), .C1(new_n292), .C2(new_n290), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n288), .B(new_n293), .C1(G77), .C2(new_n289), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n295));
  INV_X1    g0095(.A(G274), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n286), .A2(new_n284), .ZN(new_n299));
  AND2_X1   g0099(.A1(new_n299), .A2(new_n295), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G226), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n294), .A2(new_n298), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G200), .ZN(new_n303));
  INV_X1    g0103(.A(G190), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n303), .B1(new_n304), .B2(new_n302), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n282), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT72), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n280), .A2(new_n307), .A3(new_n281), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n307), .B1(new_n280), .B2(new_n281), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n306), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT73), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT10), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n277), .A2(G77), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT74), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n207), .A2(G68), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n315), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G77), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n320), .B1(new_n273), .B2(new_n276), .ZN(new_n321));
  OAI21_X1  g0121(.A(KEYINPUT74), .B1(new_n321), .B2(new_n317), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n256), .A2(G50), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n319), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n248), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(KEYINPUT11), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT11), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n324), .A2(new_n327), .A3(new_n248), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n326), .A2(new_n328), .B1(G68), .B2(new_n249), .ZN(new_n329));
  INV_X1    g0129(.A(new_n253), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n330), .A2(KEYINPUT75), .A3(new_n218), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(KEYINPUT12), .ZN(new_n332));
  AOI21_X1  g0132(.A(KEYINPUT75), .B1(new_n330), .B2(new_n218), .ZN(new_n333));
  XOR2_X1   g0133(.A(new_n332), .B(new_n333), .Z(new_n334));
  NAND2_X1  g0134(.A1(new_n300), .A2(G238), .ZN(new_n335));
  INV_X1    g0135(.A(new_n288), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n271), .A2(new_n202), .ZN(new_n337));
  NOR2_X1   g0137(.A1(G226), .A2(G1698), .ZN(new_n338));
  INV_X1    g0138(.A(G232), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n338), .B1(new_n339), .B2(G1698), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n337), .B1(new_n340), .B2(new_n289), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n335), .B(new_n298), .C1(new_n336), .C2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(KEYINPUT13), .ZN(new_n343));
  AND2_X1   g0143(.A1(new_n340), .A2(new_n289), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n288), .B1(new_n344), .B2(new_n337), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT13), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n345), .A2(new_n346), .A3(new_n298), .A4(new_n335), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n343), .A2(new_n347), .A3(G190), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n343), .A2(new_n347), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(G200), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n329), .A2(new_n334), .A3(new_n348), .A4(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(G238), .A2(G1698), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n289), .B(new_n352), .C1(new_n339), .C2(G1698), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n288), .B(new_n353), .C1(G107), .C2(new_n289), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n300), .A2(G244), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n354), .A2(new_n298), .A3(new_n355), .ZN(new_n356));
  OR2_X1    g0156(.A1(new_n356), .A2(G179), .ZN(new_n357));
  NAND2_X1  g0157(.A1(G20), .A2(G77), .ZN(new_n358));
  XNOR2_X1  g0158(.A(KEYINPUT15), .B(G87), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT8), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(G58), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n266), .A2(new_n361), .ZN(new_n362));
  OAI221_X1 g0162(.A(new_n358), .B1(new_n359), .B2(new_n274), .C1(new_n362), .C2(new_n257), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n363), .A2(new_n248), .B1(new_n320), .B2(new_n330), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n249), .A2(G77), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(G169), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n356), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n357), .A2(new_n366), .A3(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT14), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n370), .B1(new_n349), .B2(G169), .ZN(new_n371));
  AOI211_X1 g0171(.A(KEYINPUT14), .B(new_n367), .C1(new_n343), .C2(new_n347), .ZN(new_n372));
  INV_X1    g0172(.A(G179), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n349), .A2(new_n373), .ZN(new_n374));
  NOR3_X1   g0174(.A1(new_n371), .A2(new_n372), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n249), .A2(G68), .ZN(new_n376));
  INV_X1    g0176(.A(new_n328), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n327), .B1(new_n324), .B2(new_n248), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n376), .B(new_n334), .C1(new_n377), .C2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n351), .B(new_n369), .C1(new_n375), .C2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n310), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n308), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n312), .A2(new_n313), .ZN(new_n385));
  NAND2_X1  g0185(.A1(KEYINPUT73), .A2(KEYINPUT10), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n384), .A2(new_n385), .A3(new_n386), .A4(new_n306), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n302), .A2(new_n367), .ZN(new_n388));
  OR2_X1    g0188(.A1(new_n302), .A2(G179), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n280), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n314), .A2(new_n382), .A3(new_n387), .A4(new_n390), .ZN(new_n391));
  XNOR2_X1  g0191(.A(G58), .B(G68), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n392), .A2(G20), .B1(G159), .B2(new_n256), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n271), .A2(KEYINPUT3), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT3), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(G33), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n397), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT76), .ZN(new_n400));
  AND3_X1   g0200(.A1(new_n394), .A2(new_n396), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n400), .B1(new_n394), .B2(new_n396), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n207), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT7), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n399), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  OAI211_X1 g0205(.A(KEYINPUT16), .B(new_n393), .C1(new_n405), .C2(new_n218), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT16), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n404), .B1(new_n289), .B2(G20), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n218), .B1(new_n408), .B2(new_n398), .ZN(new_n409));
  INV_X1    g0209(.A(new_n393), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n407), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n406), .A2(new_n411), .A3(new_n248), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n270), .A2(new_n250), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n413), .B1(new_n330), .B2(new_n270), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  OR2_X1    g0215(.A1(G223), .A2(G1698), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n217), .A2(G1698), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n394), .A2(new_n416), .A3(new_n396), .A4(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(G33), .A2(G87), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n288), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n300), .A2(G232), .ZN(new_n422));
  AND4_X1   g0222(.A1(G179), .A2(new_n421), .A3(new_n422), .A4(new_n298), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n297), .B1(new_n420), .B2(new_n288), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n367), .B1(new_n424), .B2(new_n422), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(KEYINPUT18), .B1(new_n415), .B2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT18), .ZN(new_n429));
  AOI211_X1 g0229(.A(new_n429), .B(new_n426), .C1(new_n412), .C2(new_n414), .ZN(new_n430));
  OR2_X1    g0230(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n424), .A2(new_n304), .A3(new_n422), .ZN(new_n432));
  AND3_X1   g0232(.A1(new_n421), .A2(new_n422), .A3(new_n298), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n432), .B1(new_n433), .B2(G200), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n412), .A2(new_n414), .A3(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT17), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AND3_X1   g0237(.A1(new_n412), .A2(new_n414), .A3(new_n434), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(KEYINPUT17), .ZN(new_n439));
  INV_X1    g0239(.A(new_n366), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n356), .A2(G200), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n440), .B(new_n441), .C1(new_n304), .C2(new_n356), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n431), .A2(new_n437), .A3(new_n439), .A4(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n391), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(G45), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n445), .A2(G1), .ZN(new_n446));
  AND2_X1   g0246(.A1(KEYINPUT5), .A2(G41), .ZN(new_n447));
  NOR2_X1   g0247(.A1(KEYINPUT5), .A2(G41), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n449), .A2(G270), .A3(new_n299), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT81), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT81), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n449), .A2(new_n452), .A3(G270), .A4(new_n299), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n446), .B(G274), .C1(new_n448), .C2(new_n447), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  OR2_X1    g0256(.A1(G257), .A2(G1698), .ZN(new_n457));
  INV_X1    g0257(.A(G264), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(G1698), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n394), .A2(new_n457), .A3(new_n396), .A4(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(G303), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n460), .B1(new_n461), .B2(new_n289), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n456), .B1(new_n462), .B2(new_n288), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT82), .ZN(new_n464));
  AND3_X1   g0264(.A1(new_n454), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n464), .B1(new_n454), .B2(new_n463), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n330), .A2(new_n212), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n206), .A2(G33), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n279), .A2(G116), .A3(new_n253), .A4(new_n468), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n247), .A2(new_n224), .B1(G20), .B2(new_n212), .ZN(new_n470));
  NAND2_X1  g0270(.A1(G33), .A2(G283), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n471), .B(new_n207), .C1(G33), .C2(new_n202), .ZN(new_n472));
  AND3_X1   g0272(.A1(new_n470), .A2(KEYINPUT20), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(KEYINPUT20), .B1(new_n470), .B2(new_n472), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n467), .B(new_n469), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(G169), .ZN(new_n476));
  NOR3_X1   g0276(.A1(new_n465), .A2(new_n466), .A3(new_n476), .ZN(new_n477));
  OAI21_X1  g0277(.A(KEYINPUT21), .B1(new_n477), .B2(KEYINPUT83), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT83), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT21), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n454), .A2(new_n463), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT82), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n454), .A2(new_n463), .A3(new_n464), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n479), .B(new_n480), .C1(new_n484), .C2(new_n476), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n454), .A2(new_n463), .A3(G179), .ZN(new_n486));
  INV_X1    g0286(.A(new_n475), .ZN(new_n487));
  OR2_X1    g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(G190), .B1(new_n465), .B2(new_n466), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n482), .A2(G200), .A3(new_n483), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n489), .A2(new_n490), .A3(new_n487), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n478), .A2(new_n485), .A3(new_n488), .A4(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT24), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n394), .A2(new_n396), .A3(new_n207), .A4(G87), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(KEYINPUT22), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT22), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n289), .A2(new_n496), .A3(new_n207), .A4(G87), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n272), .A2(G116), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n203), .A2(G20), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT23), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(KEYINPUT23), .B1(new_n203), .B2(G20), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  AND4_X1   g0305(.A1(new_n493), .A2(new_n498), .A3(new_n499), .A4(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n504), .B1(new_n495), .B2(new_n497), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n493), .B1(new_n507), .B2(new_n499), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n248), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(G13), .ZN(new_n510));
  NOR3_X1   g0310(.A1(new_n500), .A2(G1), .A3(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT25), .ZN(new_n512));
  OR2_X1    g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AND3_X1   g0313(.A1(new_n279), .A2(new_n253), .A3(new_n468), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n514), .A2(G107), .B1(new_n512), .B2(new_n511), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n509), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n449), .A2(G264), .A3(new_n299), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n394), .A2(new_n396), .A3(G257), .A4(G1698), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT84), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT84), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n289), .A2(new_n520), .A3(G257), .A4(G1698), .ZN(new_n521));
  NAND2_X1  g0321(.A1(G33), .A2(G294), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n289), .A2(G250), .A3(new_n290), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n519), .A2(new_n521), .A3(new_n522), .A4(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n517), .B1(new_n524), .B2(new_n288), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n525), .A2(G179), .A3(new_n455), .ZN(new_n526));
  AOI211_X1 g0326(.A(new_n456), .B(new_n517), .C1(new_n524), .C2(new_n288), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n526), .B1(new_n367), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n516), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n524), .A2(new_n288), .ZN(new_n530));
  INV_X1    g0330(.A(new_n517), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n530), .A2(new_n304), .A3(new_n455), .A4(new_n531), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n532), .B1(new_n527), .B2(G200), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n533), .A2(new_n513), .A3(new_n509), .A4(new_n515), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n253), .A2(G97), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n514), .A2(G97), .ZN(new_n537));
  NAND2_X1  g0337(.A1(G97), .A2(G107), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(G97), .A2(G107), .ZN(new_n540));
  OAI21_X1  g0340(.A(KEYINPUT78), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT78), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n204), .A2(new_n542), .A3(new_n538), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT6), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n541), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n203), .A2(KEYINPUT6), .A3(G97), .ZN(new_n546));
  XNOR2_X1  g0346(.A(new_n546), .B(KEYINPUT77), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n207), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n203), .B1(new_n408), .B2(new_n398), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n257), .A2(new_n320), .ZN(new_n550));
  NOR3_X1   g0350(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n536), .B(new_n537), .C1(new_n551), .C2(new_n279), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n394), .A2(new_n396), .A3(G244), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT4), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n553), .A2(new_n554), .B1(G33), .B2(G283), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n554), .A2(G1698), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n289), .A2(G244), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n554), .B1(new_n289), .B2(G250), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n555), .B(new_n557), .C1(new_n290), .C2(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n456), .B1(new_n559), .B2(new_n288), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n449), .A2(G257), .A3(new_n299), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n367), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n553), .A2(new_n554), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n563), .A2(new_n557), .A3(new_n471), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n289), .A2(G250), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n290), .B1(new_n565), .B2(KEYINPUT4), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n288), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n567), .A2(G179), .A3(new_n455), .A4(new_n561), .ZN(new_n568));
  INV_X1    g0368(.A(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n552), .B1(new_n562), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n545), .A2(new_n547), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(G20), .ZN(new_n572));
  INV_X1    g0372(.A(new_n549), .ZN(new_n573));
  INV_X1    g0373(.A(new_n550), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n535), .B1(new_n575), .B2(new_n248), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n567), .A2(new_n455), .A3(new_n561), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(G200), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n567), .A2(G190), .A3(new_n455), .A4(new_n561), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n576), .A2(new_n578), .A3(new_n537), .A4(new_n579), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n529), .A2(new_n534), .A3(new_n570), .A4(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n289), .A2(new_n207), .A3(G68), .ZN(new_n582));
  INV_X1    g0382(.A(G87), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n583), .A2(new_n202), .A3(new_n203), .ZN(new_n584));
  OAI211_X1 g0384(.A(KEYINPUT19), .B(new_n584), .C1(new_n337), .C2(G20), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n274), .A2(new_n202), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n582), .B(new_n585), .C1(KEYINPUT19), .C2(new_n586), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n587), .A2(new_n248), .B1(new_n330), .B2(new_n359), .ZN(new_n588));
  INV_X1    g0388(.A(new_n359), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n514), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n219), .A2(new_n290), .ZN(new_n591));
  INV_X1    g0391(.A(G244), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(G1698), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n394), .A2(new_n591), .A3(new_n396), .A4(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n594), .B1(new_n271), .B2(new_n212), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n288), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT79), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n597), .B(G250), .C1(new_n445), .C2(G1), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n206), .A2(G45), .ZN(new_n599));
  AOI21_X1  g0399(.A(G274), .B1(KEYINPUT79), .B2(G250), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n299), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(KEYINPUT80), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT80), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n601), .A2(new_n604), .A3(new_n299), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n596), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n588), .A2(new_n590), .B1(new_n606), .B2(new_n367), .ZN(new_n607));
  AND3_X1   g0407(.A1(new_n596), .A2(new_n603), .A3(new_n605), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n373), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n608), .A2(G190), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n514), .A2(G87), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n606), .A2(G200), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n611), .A2(new_n588), .A3(new_n612), .A4(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  NOR3_X1   g0415(.A1(new_n492), .A2(new_n581), .A3(new_n615), .ZN(new_n616));
  AND2_X1   g0416(.A1(new_n444), .A2(new_n616), .ZN(G372));
  INV_X1    g0417(.A(new_n610), .ZN(new_n618));
  AND4_X1   g0418(.A1(new_n534), .A2(new_n570), .A3(new_n580), .A4(new_n614), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n478), .A2(new_n529), .A3(new_n485), .A4(new_n488), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g0421(.A(KEYINPUT85), .B1(new_n562), .B2(new_n569), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT85), .ZN(new_n623));
  INV_X1    g0423(.A(new_n577), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n623), .B(new_n568), .C1(new_n624), .C2(new_n367), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n622), .A2(new_n625), .A3(new_n552), .A4(new_n614), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT26), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n570), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n629), .A2(KEYINPUT26), .A3(new_n614), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n621), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n444), .A2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n390), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n375), .A2(new_n380), .ZN(new_n635));
  INV_X1    g0435(.A(new_n369), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n635), .B1(new_n351), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n439), .A2(new_n437), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n431), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n314), .A2(new_n387), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n634), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n633), .A2(new_n641), .ZN(G369));
  NOR2_X1   g0442(.A1(new_n510), .A2(G20), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n206), .ZN(new_n644));
  OR2_X1    g0444(.A1(new_n644), .A2(KEYINPUT27), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(KEYINPUT27), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n645), .A2(G213), .A3(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  XNOR2_X1  g0448(.A(KEYINPUT86), .B(G343), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n478), .A2(new_n485), .ZN(new_n652));
  AOI211_X1 g0452(.A(new_n487), .B(new_n651), .C1(new_n652), .C2(new_n486), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n492), .B1(new_n475), .B2(new_n650), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n529), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n650), .ZN(new_n658));
  XNOR2_X1  g0458(.A(new_n658), .B(KEYINPUT87), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n516), .A2(new_n650), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n529), .A2(new_n660), .A3(new_n534), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n656), .A2(G330), .A3(new_n662), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n650), .B1(new_n652), .B2(new_n488), .ZN(new_n664));
  AOI22_X1  g0464(.A1(new_n662), .A2(new_n664), .B1(new_n657), .B2(new_n651), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n663), .A2(new_n665), .ZN(G399));
  INV_X1    g0466(.A(new_n208), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n667), .A2(G41), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(G1), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n584), .A2(G116), .ZN(new_n671));
  OAI22_X1  g0471(.A1(new_n670), .A2(new_n671), .B1(new_n226), .B2(new_n669), .ZN(new_n672));
  XNOR2_X1  g0472(.A(new_n672), .B(KEYINPUT28), .ZN(new_n673));
  INV_X1    g0473(.A(G330), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT30), .ZN(new_n675));
  AND3_X1   g0475(.A1(new_n608), .A2(KEYINPUT88), .A3(new_n525), .ZN(new_n676));
  AOI21_X1  g0476(.A(KEYINPUT88), .B1(new_n608), .B2(new_n525), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n624), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n486), .B(KEYINPUT89), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n675), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NOR3_X1   g0480(.A1(new_n527), .A2(G179), .A3(new_n608), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n681), .A2(new_n577), .A3(new_n482), .A4(new_n483), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n608), .A2(new_n525), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT88), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n608), .A2(new_n525), .A3(KEYINPUT88), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT89), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n486), .B(new_n688), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n687), .A2(KEYINPUT30), .A3(new_n689), .A4(new_n624), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n680), .A2(new_n682), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(new_n650), .ZN(new_n692));
  NOR4_X1   g0492(.A1(new_n492), .A2(new_n581), .A3(new_n615), .A4(new_n650), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT31), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n692), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n691), .A2(KEYINPUT31), .A3(new_n650), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n674), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT29), .ZN(new_n698));
  INV_X1    g0498(.A(new_n615), .ZN(new_n699));
  OAI211_X1 g0499(.A(new_n552), .B(new_n627), .C1(new_n562), .C2(new_n569), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  AOI22_X1  g0501(.A1(KEYINPUT26), .A2(new_n626), .B1(new_n699), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n621), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n698), .B1(new_n703), .B2(new_n651), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n650), .B1(new_n621), .B2(new_n631), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n705), .A2(new_n698), .ZN(new_n706));
  NOR3_X1   g0506(.A1(new_n697), .A2(new_n704), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n673), .B1(new_n707), .B2(G1), .ZN(G364));
  AOI21_X1  g0508(.A(new_n670), .B1(G45), .B2(new_n643), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n709), .B1(new_n656), .B2(G330), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(G330), .B2(new_n656), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n224), .B1(G20), .B2(new_n367), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(G200), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(G179), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n715), .A2(G20), .A3(G190), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n715), .A2(G20), .A3(new_n304), .ZN(new_n717));
  XNOR2_X1  g0517(.A(new_n717), .B(KEYINPUT94), .ZN(new_n718));
  INV_X1    g0518(.A(G283), .ZN(new_n719));
  OAI221_X1 g0519(.A(new_n397), .B1(new_n461), .B2(new_n716), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(G179), .A2(G200), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n721), .A2(G20), .A3(new_n304), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n720), .B1(G329), .B2(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n207), .A2(new_n373), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(G190), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(new_n714), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(G326), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n726), .A2(G200), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n207), .B1(new_n721), .B2(G190), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  AOI22_X1  g0531(.A1(new_n729), .A2(G322), .B1(G294), .B2(new_n731), .ZN(new_n732));
  AND3_X1   g0532(.A1(new_n724), .A2(new_n728), .A3(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(G311), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n725), .A2(new_n304), .A3(new_n714), .ZN(new_n735));
  OR2_X1    g0535(.A1(new_n735), .A2(KEYINPUT91), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(KEYINPUT91), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n725), .A2(new_n304), .A3(G200), .ZN(new_n740));
  OR2_X1    g0540(.A1(new_n740), .A2(KEYINPUT95), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(KEYINPUT95), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  XOR2_X1   g0544(.A(KEYINPUT33), .B(G317), .Z(new_n745));
  OAI221_X1 g0545(.A(new_n733), .B1(new_n734), .B2(new_n739), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  AOI22_X1  g0546(.A1(new_n738), .A2(G77), .B1(G50), .B2(new_n727), .ZN(new_n747));
  INV_X1    g0547(.A(new_n729), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n747), .B1(new_n265), .B2(new_n748), .ZN(new_n749));
  XNOR2_X1  g0549(.A(new_n749), .B(KEYINPUT92), .ZN(new_n750));
  INV_X1    g0550(.A(new_n716), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G87), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(new_n289), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT93), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n731), .A2(G97), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n755), .B1(new_n744), .B2(new_n218), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n718), .A2(new_n203), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n754), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(G159), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n722), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n760), .B(KEYINPUT32), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n750), .A2(new_n758), .A3(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n713), .B1(new_n746), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n401), .A2(new_n402), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n667), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n227), .A2(new_n445), .ZN(new_n766));
  OAI211_X1 g0566(.A(new_n765), .B(new_n766), .C1(new_n242), .C2(new_n445), .ZN(new_n767));
  NAND3_X1  g0567(.A1(G355), .A2(new_n289), .A3(new_n208), .ZN(new_n768));
  OAI211_X1 g0568(.A(new_n767), .B(new_n768), .C1(G116), .C2(new_n208), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  OR2_X1    g0570(.A1(new_n770), .A2(KEYINPUT90), .ZN(new_n771));
  NOR2_X1   g0571(.A1(G13), .A2(G33), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(G20), .ZN(new_n774));
  AOI211_X1 g0574(.A(new_n774), .B(new_n712), .C1(new_n770), .C2(KEYINPUT90), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n763), .B1(new_n771), .B2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n774), .ZN(new_n777));
  OAI211_X1 g0577(.A(new_n776), .B(new_n709), .C1(new_n656), .C2(new_n777), .ZN(new_n778));
  AND2_X1   g0578(.A1(new_n711), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(G396));
  NOR2_X1   g0580(.A1(new_n712), .A2(new_n772), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n743), .A2(G150), .B1(G137), .B2(new_n727), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT97), .ZN(new_n784));
  INV_X1    g0584(.A(G143), .ZN(new_n785));
  OAI221_X1 g0585(.A(new_n784), .B1(new_n785), .B2(new_n748), .C1(new_n759), .C2(new_n739), .ZN(new_n786));
  INV_X1    g0586(.A(KEYINPUT34), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n723), .A2(G132), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n786), .A2(new_n787), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n764), .B1(new_n216), .B2(new_n716), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n718), .A2(new_n218), .ZN(new_n792));
  AOI211_X1 g0592(.A(new_n791), .B(new_n792), .C1(G58), .C2(new_n731), .ZN(new_n793));
  NAND4_X1  g0593(.A1(new_n788), .A2(new_n789), .A3(new_n790), .A4(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n727), .ZN(new_n795));
  INV_X1    g0595(.A(G294), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n755), .B1(new_n795), .B2(new_n461), .C1(new_n796), .C2(new_n748), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n718), .A2(new_n583), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n397), .B1(new_n722), .B2(new_n734), .ZN(new_n799));
  NOR3_X1   g0599(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  AOI22_X1  g0600(.A1(G116), .A2(new_n738), .B1(new_n743), .B2(G283), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n800), .B(new_n801), .C1(new_n203), .C2(new_n716), .ZN(new_n802));
  XOR2_X1   g0602(.A(new_n802), .B(KEYINPUT96), .Z(new_n803));
  AND2_X1   g0603(.A1(new_n794), .A2(new_n803), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n709), .B1(G77), .B2(new_n782), .C1(new_n804), .C2(new_n713), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT98), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n442), .B1(new_n440), .B2(new_n651), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(new_n369), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n369), .A2(new_n650), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n806), .B1(new_n773), .B2(new_n812), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n705), .B(new_n812), .ZN(new_n814));
  XOR2_X1   g0614(.A(new_n814), .B(new_n697), .Z(new_n815));
  OAI21_X1  g0615(.A(new_n813), .B1(new_n709), .B2(new_n815), .ZN(G384));
  NAND3_X1  g0616(.A1(new_n424), .A2(G179), .A3(new_n422), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n817), .B(new_n647), .C1(new_n433), .C2(new_n367), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n393), .B1(new_n405), .B2(new_n218), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n407), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n821), .A2(new_n248), .A3(new_n406), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n819), .B1(new_n822), .B2(new_n414), .ZN(new_n823));
  OAI21_X1  g0623(.A(KEYINPUT37), .B1(new_n823), .B2(new_n438), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(KEYINPUT102), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n415), .A2(new_n818), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT37), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n826), .A2(new_n827), .A3(new_n435), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT102), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n829), .B(KEYINPUT37), .C1(new_n823), .C2(new_n438), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n825), .A2(new_n828), .A3(new_n830), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n439), .B(new_n437), .C1(new_n428), .C2(new_n430), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n822), .A2(new_n414), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n832), .A2(new_n648), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT38), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n831), .A2(new_n834), .A3(KEYINPUT38), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n696), .A2(KEYINPUT106), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT106), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n691), .A2(new_n841), .A3(KEYINPUT31), .A4(new_n650), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n695), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n351), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n379), .B(new_n650), .C1(new_n635), .C2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n379), .A2(new_n650), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n351), .B(new_n846), .C1(new_n375), .C2(new_n380), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n849), .A2(new_n811), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n839), .A2(new_n843), .A3(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT40), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AND3_X1   g0653(.A1(new_n832), .A2(new_n415), .A3(new_n648), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n412), .A2(new_n414), .B1(new_n426), .B2(new_n647), .ZN(new_n855));
  OAI21_X1  g0655(.A(KEYINPUT37), .B1(new_n438), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n856), .A2(new_n828), .A3(KEYINPUT104), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT104), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n826), .A2(new_n858), .A3(new_n827), .A4(new_n435), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n836), .B1(new_n854), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(new_n838), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n862), .A2(new_n850), .A3(new_n843), .A4(KEYINPUT40), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n853), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n843), .A2(new_n444), .ZN(new_n865));
  XOR2_X1   g0665(.A(new_n864), .B(new_n865), .Z(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(G330), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT101), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n809), .B1(new_n705), .B2(new_n812), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n868), .B1(new_n869), .B2(new_n849), .ZN(new_n870));
  AOI211_X1 g0670(.A(new_n650), .B(new_n811), .C1(new_n621), .C2(new_n631), .ZN(new_n871));
  OAI211_X1 g0671(.A(KEYINPUT101), .B(new_n848), .C1(new_n871), .C2(new_n809), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n870), .A2(new_n839), .A3(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT39), .ZN(new_n874));
  AND3_X1   g0674(.A1(new_n831), .A2(new_n834), .A3(KEYINPUT38), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n857), .A2(new_n859), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n832), .A2(new_n415), .A3(new_n648), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT38), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n874), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n837), .A2(KEYINPUT39), .A3(new_n838), .ZN(new_n880));
  NOR3_X1   g0680(.A1(new_n375), .A2(new_n380), .A3(new_n650), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT103), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n881), .A2(new_n882), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n879), .A2(new_n880), .A3(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n431), .A2(new_n648), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n873), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT105), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n873), .A2(new_n887), .A3(KEYINPUT105), .A4(new_n889), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n867), .B(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n444), .B1(new_n706), .B2(new_n704), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n641), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n895), .B(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n898), .B1(new_n206), .B2(new_n643), .ZN(new_n899));
  OAI211_X1 g0699(.A(G116), .B(new_n225), .C1(new_n571), .C2(KEYINPUT35), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n900), .B(KEYINPUT99), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n571), .A2(KEYINPUT35), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n903), .B(KEYINPUT36), .ZN(new_n904));
  OAI21_X1  g0704(.A(G77), .B1(new_n265), .B2(new_n218), .ZN(new_n905));
  OAI22_X1  g0705(.A1(new_n905), .A2(new_n226), .B1(G50), .B2(new_n218), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n906), .A2(G1), .A3(new_n510), .ZN(new_n907));
  XOR2_X1   g0707(.A(new_n907), .B(KEYINPUT100), .Z(new_n908));
  NAND3_X1  g0708(.A1(new_n899), .A2(new_n904), .A3(new_n908), .ZN(G367));
  NAND2_X1  g0709(.A1(new_n588), .A2(new_n612), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n650), .ZN(new_n911));
  AOI21_X1  g0711(.A(KEYINPUT107), .B1(new_n699), .B2(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n610), .A2(new_n911), .ZN(new_n913));
  MUX2_X1   g0713(.A(new_n912), .B(KEYINPUT107), .S(new_n913), .Z(new_n914));
  INV_X1    g0714(.A(KEYINPUT43), .ZN(new_n915));
  OR2_X1    g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n622), .A2(new_n552), .A3(new_n625), .A4(new_n650), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n552), .A2(new_n650), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n570), .A2(new_n580), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n662), .A2(new_n664), .A3(new_n920), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n921), .B(KEYINPUT42), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n920), .B(KEYINPUT108), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n657), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n650), .B1(new_n924), .B2(new_n570), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n916), .B1(new_n922), .B2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n663), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n926), .A2(new_n927), .A3(new_n923), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n914), .A2(new_n915), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n927), .A2(new_n923), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n930), .B(new_n916), .C1(new_n922), .C2(new_n925), .ZN(new_n931));
  AND3_X1   g0731(.A1(new_n928), .A2(new_n929), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n929), .B1(new_n928), .B2(new_n931), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n668), .B(KEYINPUT41), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n661), .B(new_n659), .C1(new_n655), .C2(new_n674), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n663), .A2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n664), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n663), .A2(new_n937), .A3(new_n664), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n942), .A2(KEYINPUT110), .A3(new_n707), .ZN(new_n943));
  INV_X1    g0743(.A(new_n665), .ZN(new_n944));
  INV_X1    g0744(.A(new_n920), .ZN(new_n945));
  NAND2_X1  g0745(.A1(KEYINPUT109), .A2(KEYINPUT44), .ZN(new_n946));
  OR2_X1    g0746(.A1(KEYINPUT109), .A2(KEYINPUT44), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n944), .A2(new_n945), .A3(new_n946), .A4(new_n947), .ZN(new_n948));
  OAI211_X1 g0748(.A(KEYINPUT109), .B(KEYINPUT44), .C1(new_n665), .C2(new_n920), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n662), .A2(new_n664), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n657), .A2(new_n651), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n951), .A2(new_n952), .A3(new_n920), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT45), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n927), .B1(new_n950), .B2(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n940), .A2(new_n707), .A3(new_n941), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT110), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT45), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n953), .B(new_n959), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n960), .A2(new_n663), .A3(new_n949), .A4(new_n948), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n943), .A2(new_n955), .A3(new_n958), .A4(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n936), .B1(new_n962), .B2(new_n707), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n206), .B1(new_n643), .B2(G45), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n934), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n914), .A2(new_n774), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n774), .A2(new_n712), .ZN(new_n968));
  INV_X1    g0768(.A(new_n765), .ZN(new_n969));
  OAI221_X1 g0769(.A(new_n968), .B1(new_n208), .B2(new_n359), .C1(new_n233), .C2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n709), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n289), .B1(new_n717), .B2(new_n320), .C1(new_n265), .C2(new_n716), .ZN(new_n972));
  OAI22_X1  g0772(.A1(new_n795), .A2(new_n785), .B1(new_n730), .B2(new_n218), .ZN(new_n973));
  AOI211_X1 g0773(.A(new_n972), .B(new_n973), .C1(G137), .C2(new_n723), .ZN(new_n974));
  AOI22_X1  g0774(.A1(G50), .A2(new_n738), .B1(new_n743), .B2(G159), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n974), .B(new_n975), .C1(new_n258), .C2(new_n748), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n748), .A2(new_n461), .B1(new_n730), .B2(new_n203), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(G311), .B2(new_n727), .ZN(new_n978));
  AOI22_X1  g0778(.A1(G283), .A2(new_n738), .B1(new_n743), .B2(G294), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n716), .A2(new_n212), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT46), .Z(new_n981));
  AOI21_X1  g0781(.A(new_n764), .B1(G317), .B2(new_n723), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n978), .A2(new_n979), .A3(new_n981), .A4(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n717), .A2(new_n202), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n976), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT47), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n971), .B1(new_n986), .B2(new_n712), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n967), .A2(new_n970), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n966), .A2(new_n988), .ZN(G387));
  NAND2_X1  g0789(.A1(new_n943), .A2(new_n958), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n990), .B(new_n668), .C1(new_n707), .C2(new_n942), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n738), .A2(G303), .B1(G322), .B2(new_n727), .ZN(new_n992));
  INV_X1    g0792(.A(G317), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n992), .B1(new_n734), .B2(new_n744), .C1(new_n993), .C2(new_n748), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT114), .Z(new_n995));
  AOI22_X1  g0795(.A1(new_n995), .A2(KEYINPUT48), .B1(G283), .B2(new_n731), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n996), .B1(KEYINPUT48), .B2(new_n995), .C1(new_n796), .C2(new_n716), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT49), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n723), .A2(G326), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n997), .A2(new_n998), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n717), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n764), .B1(G116), .B2(new_n1002), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .A4(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n718), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n1005), .A2(G97), .B1(G150), .B2(new_n723), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n751), .A2(G77), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1006), .A2(new_n764), .A3(new_n1007), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n1008), .B(KEYINPUT112), .Z(new_n1009));
  AOI22_X1  g0809(.A1(new_n729), .A2(G50), .B1(new_n589), .B2(new_n731), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n1011), .A2(KEYINPUT113), .B1(G159), .B2(new_n727), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(KEYINPUT113), .B2(new_n1011), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(new_n270), .B2(new_n743), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1009), .B(new_n1014), .C1(new_n218), .C2(new_n739), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1004), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n712), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n662), .A2(new_n777), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n362), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(new_n216), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n1020), .A2(KEYINPUT50), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n671), .B1(new_n1020), .B2(KEYINPUT50), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(G68), .A2(G77), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1021), .A2(new_n1022), .A3(new_n445), .A4(new_n1023), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1024), .B(new_n765), .C1(new_n238), .C2(new_n445), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n671), .A2(new_n208), .A3(new_n289), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(G107), .B2(new_n208), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT111), .Z(new_n1028));
  NAND2_X1  g0828(.A1(new_n1025), .A2(new_n1028), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n971), .B(new_n1018), .C1(new_n968), .C2(new_n1029), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n965), .A2(new_n942), .B1(new_n1017), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n991), .A2(new_n1031), .ZN(G393));
  NAND2_X1  g0832(.A1(new_n955), .A2(new_n961), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n990), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1034), .A2(new_n668), .A3(new_n962), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n955), .A2(new_n961), .A3(new_n965), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n748), .A2(new_n759), .B1(new_n795), .B2(new_n258), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT51), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  AND2_X1   g0839(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n1039), .B(new_n1040), .C1(new_n1019), .C2(new_n738), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n764), .B1(new_n218), .B2(new_n716), .C1(new_n785), .C2(new_n722), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n798), .B(new_n1042), .C1(G77), .C2(new_n731), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1041), .B(new_n1043), .C1(new_n216), .C2(new_n744), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n739), .A2(new_n796), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n289), .B1(new_n723), .B2(G322), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n212), .B2(new_n730), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n1047), .B(new_n757), .C1(G283), .C2(new_n751), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n748), .A2(new_n734), .B1(new_n795), .B2(new_n993), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT52), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n1049), .A2(new_n1050), .B1(G303), .B2(new_n743), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1048), .B(new_n1051), .C1(new_n1050), .C2(new_n1049), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1044), .B1(new_n1045), .B2(new_n1052), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT115), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n971), .B1(new_n1054), .B2(new_n712), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n968), .B1(new_n202), .B2(new_n208), .C1(new_n969), .C2(new_n245), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1055), .B(new_n1056), .C1(new_n777), .C2(new_n923), .ZN(new_n1057));
  AND2_X1   g0857(.A1(new_n1036), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1035), .A2(new_n1058), .ZN(G390));
  OAI21_X1  g0859(.A(new_n885), .B1(new_n869), .B2(new_n849), .ZN(new_n1060));
  AOI21_X1  g0860(.A(KEYINPUT38), .B1(new_n831), .B2(new_n834), .ZN(new_n1061));
  NOR3_X1   g0861(.A1(new_n875), .A2(new_n1061), .A3(new_n874), .ZN(new_n1062));
  AOI21_X1  g0862(.A(KEYINPUT39), .B1(new_n861), .B2(new_n838), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1060), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  AND3_X1   g0864(.A1(new_n703), .A2(new_n651), .A3(new_n808), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n848), .B1(new_n1065), .B2(new_n809), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1066), .A2(new_n862), .A3(new_n885), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n694), .B1(new_n616), .B2(new_n651), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n692), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n696), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n811), .A2(new_n674), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1070), .A2(new_n848), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(new_n1073));
  AND3_X1   g0873(.A1(new_n1064), .A2(new_n1067), .A3(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n840), .A2(new_n842), .ZN(new_n1075));
  AND4_X1   g0875(.A1(new_n488), .A2(new_n478), .A3(new_n485), .A4(new_n491), .ZN(new_n1076));
  AND4_X1   g0876(.A1(new_n529), .A2(new_n534), .A3(new_n570), .A4(new_n580), .ZN(new_n1077));
  NAND4_X1  g0877(.A1(new_n1076), .A2(new_n1077), .A3(new_n699), .A4(new_n651), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n1078), .A2(KEYINPUT31), .B1(new_n650), .B2(new_n691), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n848), .B(new_n1071), .C1(new_n1075), .C2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1082));
  OR2_X1    g0882(.A1(new_n1074), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(new_n965), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n773), .B1(new_n879), .B2(new_n880), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n792), .B1(G294), .B2(new_n723), .ZN(new_n1086));
  XOR2_X1   g0886(.A(new_n1086), .B(KEYINPUT116), .Z(new_n1087));
  AOI22_X1  g0887(.A1(new_n729), .A2(G116), .B1(new_n727), .B2(G283), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n1088), .B1(new_n320), .B2(new_n730), .C1(new_n739), .C2(new_n202), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(G107), .B2(new_n743), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1087), .A2(new_n397), .A3(new_n752), .A4(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(G132), .ZN(new_n1092));
  INV_X1    g0892(.A(G128), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n748), .A2(new_n1092), .B1(new_n795), .B2(new_n1093), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n397), .B(new_n1094), .C1(G50), .C2(new_n1002), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n723), .A2(G125), .ZN(new_n1096));
  XOR2_X1   g0896(.A(KEYINPUT54), .B(G143), .Z(new_n1097));
  AOI22_X1  g0897(.A1(G137), .A2(new_n743), .B1(new_n738), .B2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n716), .A2(new_n258), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT53), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n1099), .A2(new_n1100), .B1(new_n759), .B2(new_n730), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(new_n1100), .B2(new_n1099), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1095), .A2(new_n1096), .A3(new_n1098), .A4(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n713), .B1(new_n1091), .B2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n270), .A2(new_n782), .ZN(new_n1105));
  OR4_X1    g0905(.A1(new_n971), .A2(new_n1085), .A3(new_n1104), .A4(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1084), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n843), .A2(G330), .A3(new_n444), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1108), .A2(new_n896), .A3(new_n641), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n869), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n848), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1110), .B1(new_n1081), .B2(new_n1111), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1065), .A2(new_n809), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1071), .ZN(new_n1114));
  AND2_X1   g0914(.A1(new_n840), .A2(new_n842), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1114), .B1(new_n1115), .B2(new_n695), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1072), .B(new_n1113), .C1(new_n1116), .C2(new_n848), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1109), .B1(new_n1112), .B2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1118), .B1(new_n1074), .B2(new_n1082), .ZN(new_n1119));
  AND2_X1   g0919(.A1(new_n1119), .A2(new_n668), .ZN(new_n1120));
  OR2_X1    g0920(.A1(new_n1083), .A2(new_n1118), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1107), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(G378));
  NAND2_X1  g0923(.A1(new_n640), .A2(new_n390), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT55), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n280), .A2(new_n648), .ZN(new_n1126));
  XOR2_X1   g0926(.A(new_n1126), .B(KEYINPUT56), .Z(new_n1127));
  XNOR2_X1  g0927(.A(new_n1125), .B(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n853), .A2(G330), .A3(new_n863), .ZN(new_n1130));
  AND3_X1   g0930(.A1(new_n892), .A2(new_n893), .A3(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1130), .B1(new_n892), .B2(new_n893), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1129), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1130), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n894), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n892), .A2(new_n893), .A3(new_n1130), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1135), .A2(new_n1128), .A3(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1133), .A2(new_n1137), .A3(new_n965), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n751), .A2(new_n1097), .B1(new_n731), .B2(G150), .ZN(new_n1139));
  INV_X1    g0939(.A(G125), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1139), .B1(new_n1140), .B2(new_n795), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(G137), .B2(new_n738), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n1142), .B1(new_n1093), .B2(new_n748), .C1(new_n1092), .C2(new_n744), .ZN(new_n1143));
  XOR2_X1   g0943(.A(new_n1143), .B(KEYINPUT59), .Z(new_n1144));
  AOI21_X1  g0944(.A(G41), .B1(new_n1002), .B2(G159), .ZN(new_n1145));
  XOR2_X1   g0945(.A(KEYINPUT117), .B(G124), .Z(new_n1146));
  AOI21_X1  g0946(.A(G33), .B1(new_n723), .B2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1144), .A2(new_n1145), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1002), .A2(G58), .ZN(new_n1149));
  INV_X1    g0949(.A(G41), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1007), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n764), .B1(G68), .B2(new_n731), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1152), .B1(new_n203), .B2(new_n748), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n1151), .B(new_n1153), .C1(G283), .C2(new_n723), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(G97), .A2(new_n743), .B1(new_n738), .B2(new_n589), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1154), .B(new_n1155), .C1(new_n212), .C2(new_n795), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1156), .B(KEYINPUT58), .ZN(new_n1157));
  AOI21_X1  g0957(.A(G41), .B1(new_n764), .B2(G33), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1148), .B(new_n1157), .C1(G50), .C2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n971), .B1(new_n1159), .B2(new_n712), .ZN(new_n1160));
  OAI221_X1 g0960(.A(new_n1160), .B1(G50), .B2(new_n782), .C1(new_n1129), .C2(new_n773), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1138), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1109), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1119), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(KEYINPUT118), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT118), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1119), .A2(new_n1167), .A3(new_n1164), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1133), .A2(new_n1137), .A3(new_n1166), .A4(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT57), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n668), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n1133), .A2(new_n1137), .ZN(new_n1172));
  AND3_X1   g0972(.A1(new_n1119), .A2(new_n1167), .A3(new_n1164), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1167), .B1(new_n1119), .B2(new_n1164), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(KEYINPUT57), .B1(new_n1172), .B2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1163), .B1(new_n1171), .B2(new_n1176), .ZN(G375));
  AND3_X1   g0977(.A1(new_n1112), .A2(new_n1109), .A3(new_n1117), .ZN(new_n1178));
  NOR3_X1   g0978(.A1(new_n1178), .A2(new_n1118), .A3(new_n936), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1179), .B(KEYINPUT119), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1112), .A2(new_n1117), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n965), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n849), .A2(new_n772), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n764), .B1(new_n795), .B2(new_n1092), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n1149), .B1(new_n1093), .B2(new_n722), .C1(new_n759), .C2(new_n716), .ZN(new_n1185));
  AOI211_X1 g0985(.A(new_n1184), .B(new_n1185), .C1(G137), .C2(new_n729), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(G150), .A2(new_n738), .B1(new_n743), .B2(new_n1097), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1186), .B(new_n1187), .C1(new_n216), .C2(new_n730), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n397), .B1(new_n722), .B2(new_n461), .C1(new_n795), .C2(new_n796), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(G77), .B2(new_n1005), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(G107), .A2(new_n738), .B1(new_n743), .B2(G116), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1190), .B(new_n1191), .C1(new_n202), .C2(new_n716), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n729), .A2(G283), .B1(new_n589), .B2(new_n731), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n1193), .B(KEYINPUT121), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1188), .B1(new_n1192), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(new_n712), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n709), .B1(G68), .B2(new_n782), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT120), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1183), .A2(new_n1196), .A3(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1182), .A2(KEYINPUT122), .A3(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT122), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n964), .B1(new_n1112), .B2(new_n1117), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1199), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1201), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1200), .A2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1180), .A2(new_n1205), .ZN(G381));
  NAND3_X1  g1006(.A1(new_n1122), .A2(new_n1138), .A3(new_n1161), .ZN(new_n1207));
  AND4_X1   g1007(.A1(new_n1137), .A2(new_n1133), .A3(new_n1166), .A4(new_n1168), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n669), .B1(new_n1208), .B2(KEYINPUT57), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1207), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n991), .A2(new_n779), .A3(new_n1031), .ZN(new_n1212));
  NOR4_X1   g1012(.A1(G387), .A2(G384), .A3(G390), .A4(new_n1212), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1211), .A2(new_n1213), .A3(new_n1205), .A4(new_n1180), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(new_n1214), .B(KEYINPUT123), .ZN(G407));
  INV_X1    g1015(.A(G213), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n649), .A2(new_n1216), .ZN(new_n1217));
  XOR2_X1   g1017(.A(new_n1217), .B(KEYINPUT124), .Z(new_n1218));
  XOR2_X1   g1018(.A(new_n1218), .B(KEYINPUT125), .Z(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1211), .A2(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(G407), .A2(G213), .A3(new_n1221), .ZN(G409));
  AOI21_X1  g1022(.A(G390), .B1(new_n966), .B2(new_n988), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(G393), .A2(G396), .ZN(new_n1225));
  AND3_X1   g1025(.A1(new_n1225), .A2(KEYINPUT127), .A3(new_n1212), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n966), .A2(new_n988), .A3(G390), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1224), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  AND3_X1   g1028(.A1(new_n966), .A2(new_n988), .A3(G390), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1225), .A2(new_n1212), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1223), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1228), .B1(new_n1231), .B2(new_n1226), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1175), .A2(KEYINPUT57), .A3(new_n1137), .A4(new_n1133), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1210), .A2(new_n668), .A3(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1122), .B1(new_n1234), .B2(new_n1163), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1169), .A2(new_n936), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1207), .A2(new_n1236), .ZN(new_n1237));
  NOR3_X1   g1037(.A1(new_n1235), .A2(new_n1220), .A3(new_n1237), .ZN(new_n1238));
  OAI21_X1  g1038(.A(KEYINPUT60), .B1(new_n1178), .B2(new_n1118), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT60), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1240), .B1(new_n1181), .B2(new_n1164), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1239), .A2(new_n668), .A3(new_n1241), .ZN(new_n1242));
  AND3_X1   g1042(.A1(new_n1242), .A2(G384), .A3(new_n1205), .ZN(new_n1243));
  AOI21_X1  g1043(.A(G384), .B1(new_n1242), .B2(new_n1205), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT63), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1232), .B1(new_n1238), .B2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT61), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1218), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1237), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1162), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n1251), .B(new_n1252), .C1(new_n1253), .C2(new_n1122), .ZN(new_n1254));
  OAI211_X1 g1054(.A(G2897), .B(new_n1220), .C1(new_n1243), .C2(new_n1244), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1218), .A2(G2897), .ZN(new_n1256));
  AOI21_X1  g1056(.A(KEYINPUT126), .B1(new_n1245), .B2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT126), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1256), .ZN(new_n1259));
  NOR4_X1   g1059(.A1(new_n1243), .A2(new_n1244), .A3(new_n1258), .A4(new_n1259), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1255), .B1(new_n1257), .B2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1247), .B1(new_n1254), .B2(new_n1262), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1254), .A2(new_n1246), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1249), .B(new_n1250), .C1(new_n1263), .C2(new_n1264), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1219), .B(new_n1252), .C1(new_n1253), .C2(new_n1122), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT62), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1261), .A2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1266), .A2(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1237), .B1(G375), .B2(G378), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1270), .A2(new_n1267), .A3(new_n1251), .A4(new_n1245), .ZN(new_n1271));
  AOI21_X1  g1071(.A(KEYINPUT61), .B1(new_n1246), .B2(KEYINPUT62), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1269), .A2(new_n1271), .A3(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(new_n1232), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1265), .A2(new_n1274), .ZN(G405));
  OR3_X1    g1075(.A1(new_n1235), .A2(new_n1211), .A3(new_n1245), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1245), .B1(new_n1235), .B2(new_n1211), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1232), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(new_n1278), .B(new_n1279), .ZN(G402));
endmodule


