//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 0 0 1 0 1 1 0 1 0 0 0 1 1 0 1 0 0 1 1 1 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 1 1 1 1 1 1 1 0 0 1 0 0 0 1 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n744,
    new_n745, new_n746, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n850, new_n852, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n982, new_n983;
  INV_X1    g000(.A(KEYINPUT10), .ZN(new_n202));
  XOR2_X1   g001(.A(G99gat), .B(G106gat), .Z(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT97), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n205), .A2(KEYINPUT7), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(KEYINPUT7), .ZN(new_n207));
  AND2_X1   g006(.A1(G85gat), .A2(G92gat), .ZN(new_n208));
  AND3_X1   g007(.A1(new_n207), .A2(new_n208), .A3(KEYINPUT98), .ZN(new_n209));
  AOI21_X1  g008(.A(KEYINPUT98), .B1(new_n207), .B2(new_n208), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n206), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT7), .ZN(new_n212));
  OAI211_X1 g011(.A(G85gat), .B(G92gat), .C1(new_n212), .C2(KEYINPUT97), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT98), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n206), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n207), .A2(new_n208), .A3(KEYINPUT98), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n211), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(G99gat), .A2(G106gat), .ZN(new_n220));
  INV_X1    g019(.A(G85gat), .ZN(new_n221));
  INV_X1    g020(.A(G92gat), .ZN(new_n222));
  AOI22_X1  g021(.A1(KEYINPUT8), .A2(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n204), .B1(new_n219), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(new_n223), .ZN(new_n225));
  AOI211_X1 g024(.A(new_n203), .B(new_n225), .C1(new_n211), .C2(new_n218), .ZN(new_n226));
  XOR2_X1   g025(.A(G71gat), .B(G78gat), .Z(new_n227));
  INV_X1    g026(.A(KEYINPUT9), .ZN(new_n228));
  XNOR2_X1  g027(.A(G57gat), .B(G64gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n227), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT93), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n227), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT94), .ZN(new_n234));
  INV_X1    g033(.A(G64gat), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n234), .B1(new_n235), .B2(G57gat), .ZN(new_n236));
  INV_X1    g035(.A(G57gat), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n237), .A2(KEYINPUT94), .A3(G64gat), .ZN(new_n238));
  OAI211_X1 g037(.A(new_n236), .B(new_n238), .C1(new_n237), .C2(G64gat), .ZN(new_n239));
  INV_X1    g038(.A(G71gat), .ZN(new_n240));
  INV_X1    g039(.A(G78gat), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n228), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT95), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT95), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n244), .B(new_n228), .C1(new_n240), .C2(new_n241), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n233), .A2(new_n239), .A3(new_n243), .A4(new_n245), .ZN(new_n246));
  OAI211_X1 g045(.A(new_n227), .B(KEYINPUT93), .C1(new_n228), .C2(new_n229), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n232), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  NOR3_X1   g047(.A1(new_n224), .A2(new_n226), .A3(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT100), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n202), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(G230gat), .A2(G233gat), .ZN(new_n252));
  INV_X1    g051(.A(new_n248), .ZN(new_n253));
  NOR3_X1   g052(.A1(new_n209), .A2(new_n210), .A3(new_n206), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n216), .B1(new_n215), .B2(new_n217), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n223), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(new_n203), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n219), .A2(new_n204), .A3(new_n223), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n253), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n257), .A2(new_n258), .ZN(new_n261));
  OAI211_X1 g060(.A(KEYINPUT100), .B(KEYINPUT10), .C1(new_n261), .C2(new_n248), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n251), .A2(new_n252), .A3(new_n260), .A4(new_n262), .ZN(new_n263));
  OAI211_X1 g062(.A(G230gat), .B(G233gat), .C1(new_n259), .C2(new_n249), .ZN(new_n264));
  XNOR2_X1  g063(.A(G120gat), .B(G148gat), .ZN(new_n265));
  INV_X1    g064(.A(G176gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n265), .B(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(G204gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n267), .B(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n263), .A2(new_n264), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(KEYINPUT102), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n252), .B(KEYINPUT101), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n251), .A2(new_n260), .A3(new_n273), .A4(new_n262), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n270), .B1(new_n274), .B2(new_n264), .ZN(new_n275));
  OR2_X1    g074(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT102), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  NOR2_X1   g079(.A1(G29gat), .A2(G36gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT14), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT14), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n283), .B1(G29gat), .B2(G36gat), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n282), .B1(new_n284), .B2(new_n281), .ZN(new_n285));
  XNOR2_X1  g084(.A(G43gat), .B(G50gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT15), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(KEYINPUT90), .B(G50gat), .ZN(new_n289));
  INV_X1    g088(.A(G43gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT15), .B1(G43gat), .B2(G50gat), .ZN(new_n292));
  AOI22_X1  g091(.A1(new_n291), .A2(new_n292), .B1(KEYINPUT15), .B2(new_n286), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n288), .B1(new_n293), .B2(new_n285), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT17), .ZN(new_n295));
  XNOR2_X1  g094(.A(G15gat), .B(G22gat), .ZN(new_n296));
  INV_X1    g095(.A(G1gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(KEYINPUT16), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n296), .A2(G1gat), .ZN(new_n301));
  NOR3_X1   g100(.A1(new_n300), .A2(new_n301), .A3(G8gat), .ZN(new_n302));
  INV_X1    g101(.A(G8gat), .ZN(new_n303));
  OR2_X1    g102(.A1(new_n296), .A2(G1gat), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n303), .B1(new_n304), .B2(new_n299), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT17), .ZN(new_n307));
  OAI211_X1 g106(.A(new_n307), .B(new_n288), .C1(new_n293), .C2(new_n285), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n295), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  OAI221_X1 g108(.A(new_n288), .B1(new_n293), .B2(new_n285), .C1(new_n302), .C2(new_n305), .ZN(new_n310));
  NAND2_X1  g109(.A1(G229gat), .A2(G233gat), .ZN(new_n311));
  XOR2_X1   g110(.A(new_n311), .B(KEYINPUT91), .Z(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n309), .A2(new_n310), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(KEYINPUT92), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT18), .ZN(new_n316));
  INV_X1    g115(.A(new_n294), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n317), .B(new_n306), .ZN(new_n318));
  XOR2_X1   g117(.A(new_n312), .B(KEYINPUT13), .Z(new_n319));
  NOR2_X1   g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT18), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n314), .A2(KEYINPUT92), .A3(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n316), .A2(new_n321), .A3(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(G113gat), .B(G141gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n325), .B(G197gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n326), .B(KEYINPUT11), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n327), .B(G169gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n328), .B(KEYINPUT12), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n324), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT12), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n328), .B(new_n331), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n332), .A2(new_n316), .A3(new_n321), .A4(new_n323), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n280), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(G169gat), .ZN(new_n337));
  OAI21_X1  g136(.A(KEYINPUT67), .B1(new_n337), .B2(new_n266), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT67), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n339), .A2(G169gat), .A3(G176gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n342));
  OR3_X1    g141(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(G183gat), .A2(G190gat), .ZN(new_n345));
  INV_X1    g144(.A(G190gat), .ZN(new_n346));
  AND2_X1   g145(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n347));
  NOR2_X1   g146(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n348));
  OAI211_X1 g147(.A(KEYINPUT28), .B(new_n346), .C1(new_n347), .C2(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n349), .B(KEYINPUT71), .ZN(new_n350));
  INV_X1    g149(.A(new_n348), .ZN(new_n351));
  XNOR2_X1  g150(.A(KEYINPUT70), .B(G183gat), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT27), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n351), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(KEYINPUT28), .B1(new_n354), .B2(new_n346), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n344), .B(new_n345), .C1(new_n350), .C2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT23), .ZN(new_n357));
  NOR3_X1   g156(.A1(new_n357), .A2(G169gat), .A3(G176gat), .ZN(new_n358));
  AOI21_X1  g157(.A(KEYINPUT23), .B1(new_n337), .B2(new_n266), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT66), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n361), .B(KEYINPUT24), .C1(G183gat), .C2(G190gat), .ZN(new_n362));
  INV_X1    g161(.A(new_n345), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT24), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT66), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n362), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  OR2_X1    g165(.A1(G183gat), .A2(G190gat), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n367), .A2(new_n361), .A3(KEYINPUT24), .A4(new_n345), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n360), .A2(new_n366), .A3(new_n341), .A4(new_n368), .ZN(new_n369));
  XOR2_X1   g168(.A(KEYINPUT65), .B(KEYINPUT25), .Z(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n363), .B1(KEYINPUT69), .B2(KEYINPUT24), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT69), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n345), .A2(new_n373), .A3(new_n364), .ZN(new_n374));
  XOR2_X1   g173(.A(KEYINPUT70), .B(G183gat), .Z(new_n375));
  OAI211_X1 g174(.A(new_n372), .B(new_n374), .C1(new_n375), .C2(G190gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT25), .ZN(new_n377));
  AND3_X1   g176(.A1(new_n338), .A2(KEYINPUT68), .A3(new_n340), .ZN(new_n378));
  AOI21_X1  g177(.A(KEYINPUT68), .B1(new_n338), .B2(new_n340), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n360), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n371), .B1(new_n377), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n356), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(G120gat), .ZN(new_n383));
  AND2_X1   g182(.A1(new_n383), .A2(G113gat), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n383), .A2(G113gat), .ZN(new_n385));
  OAI21_X1  g184(.A(KEYINPUT73), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(G113gat), .B(G120gat), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT73), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT1), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n386), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(G127gat), .ZN(new_n392));
  OR3_X1    g191(.A1(new_n392), .A2(KEYINPUT72), .A3(G134gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(G127gat), .B(G134gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT72), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n391), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n394), .B(new_n390), .C1(new_n384), .C2(new_n385), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n382), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(G227gat), .A2(G233gat), .ZN(new_n401));
  XOR2_X1   g200(.A(new_n401), .B(KEYINPUT64), .Z(new_n402));
  NAND3_X1  g201(.A1(new_n356), .A2(new_n381), .A3(new_n398), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n400), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(KEYINPUT32), .ZN(new_n405));
  XNOR2_X1  g204(.A(G15gat), .B(G43gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n406), .B(G71gat), .ZN(new_n407));
  INV_X1    g206(.A(G99gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n407), .B(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT74), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT33), .ZN(new_n411));
  AND3_X1   g210(.A1(new_n404), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n410), .B1(new_n404), .B2(new_n411), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n405), .B(new_n409), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n409), .A2(KEYINPUT33), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n404), .A2(KEYINPUT32), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(KEYINPUT75), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT75), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n404), .A2(new_n418), .A3(KEYINPUT32), .A4(new_n415), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n414), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n400), .A2(new_n403), .ZN(new_n422));
  INV_X1    g221(.A(new_n402), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT34), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n425), .B1(new_n423), .B2(KEYINPUT76), .ZN(new_n426));
  AND2_X1   g225(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n424), .A2(new_n426), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n421), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n414), .A2(new_n429), .A3(new_n420), .ZN(new_n432));
  XNOR2_X1  g231(.A(G8gat), .B(G36gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n433), .B(new_n235), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n434), .B(new_n222), .ZN(new_n435));
  XNOR2_X1  g234(.A(G197gat), .B(G204gat), .ZN(new_n436));
  NOR2_X1   g235(.A1(G211gat), .A2(G218gat), .ZN(new_n437));
  AND2_X1   g236(.A1(new_n437), .A2(KEYINPUT22), .ZN(new_n438));
  INV_X1    g237(.A(G211gat), .ZN(new_n439));
  INV_X1    g238(.A(G218gat), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n436), .B1(new_n438), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT77), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n442), .B(new_n443), .ZN(new_n444));
  AOI211_X1 g243(.A(new_n437), .B(new_n441), .C1(new_n436), .C2(KEYINPUT22), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT29), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n382), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(G226gat), .ZN(new_n450));
  INV_X1    g249(.A(G233gat), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n449), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n453), .B1(new_n356), .B2(new_n381), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n447), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n452), .B1(new_n382), .B2(new_n448), .ZN(new_n458));
  NOR3_X1   g257(.A1(new_n458), .A2(new_n446), .A3(new_n455), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n435), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n454), .A2(new_n447), .A3(new_n456), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n446), .B1(new_n458), .B2(new_n455), .ZN(new_n462));
  INV_X1    g261(.A(new_n435), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n460), .A2(KEYINPUT30), .A3(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT30), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n461), .A2(new_n462), .A3(new_n466), .A4(new_n463), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  XOR2_X1   g267(.A(G78gat), .B(G106gat), .Z(new_n469));
  NAND2_X1  g268(.A1(G228gat), .A2(G233gat), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n469), .B(new_n470), .ZN(new_n471));
  XNOR2_X1  g270(.A(KEYINPUT31), .B(G50gat), .ZN(new_n472));
  XOR2_X1   g271(.A(new_n471), .B(new_n472), .Z(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT3), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n475), .B1(new_n446), .B2(KEYINPUT29), .ZN(new_n476));
  XNOR2_X1  g275(.A(KEYINPUT78), .B(KEYINPUT2), .ZN(new_n477));
  NAND2_X1  g276(.A1(G155gat), .A2(G162gat), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(KEYINPUT79), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(G141gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(G148gat), .ZN(new_n482));
  INV_X1    g281(.A(G148gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(G141gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT79), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT2), .ZN(new_n487));
  AND2_X1   g286(.A1(new_n487), .A2(KEYINPUT78), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n487), .A2(KEYINPUT78), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n486), .B(new_n478), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n480), .A2(new_n485), .A3(new_n490), .ZN(new_n491));
  NOR2_X1   g290(.A1(G155gat), .A2(G162gat), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n479), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  AND2_X1   g293(.A1(KEYINPUT80), .A2(G148gat), .ZN(new_n495));
  NOR2_X1   g294(.A1(KEYINPUT80), .A2(G148gat), .ZN(new_n496));
  OAI21_X1  g295(.A(G141gat), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n492), .A2(new_n487), .ZN(new_n498));
  AOI22_X1  g297(.A1(new_n497), .A2(new_n482), .B1(new_n478), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n494), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n476), .A2(new_n501), .ZN(new_n502));
  XOR2_X1   g301(.A(KEYINPUT85), .B(G22gat), .Z(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n499), .B1(new_n491), .B2(new_n493), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(new_n475), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n447), .B1(new_n448), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n502), .A2(new_n504), .A3(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n504), .B1(new_n508), .B2(new_n502), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n474), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n511), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n513), .A2(new_n509), .A3(new_n473), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  AND4_X1   g314(.A1(new_n431), .A2(new_n432), .A3(new_n468), .A4(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT87), .ZN(new_n517));
  NAND2_X1  g316(.A1(G225gat), .A2(G233gat), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n399), .A2(new_n505), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n505), .A2(new_n396), .A3(new_n397), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n519), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT5), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n501), .A2(KEYINPUT3), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n525), .A2(new_n398), .A3(new_n506), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT81), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT81), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n525), .A2(new_n528), .A3(new_n398), .A4(new_n506), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n519), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT4), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n399), .A2(KEYINPUT82), .A3(new_n531), .A4(new_n505), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n505), .A2(new_n531), .A3(new_n396), .A4(new_n397), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT82), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n521), .A2(KEYINPUT4), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n532), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n524), .B1(new_n530), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n519), .A2(KEYINPUT5), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  AOI221_X4 g339(.A(new_n540), .B1(new_n536), .B2(new_n533), .C1(new_n527), .C2(new_n529), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n517), .B1(new_n538), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n505), .A2(new_n475), .ZN(new_n543));
  AOI211_X1 g342(.A(KEYINPUT3), .B(new_n499), .C1(new_n491), .C2(new_n493), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n528), .B1(new_n545), .B2(new_n398), .ZN(new_n546));
  AND4_X1   g345(.A1(new_n528), .A2(new_n525), .A3(new_n398), .A4(new_n506), .ZN(new_n547));
  OAI211_X1 g346(.A(new_n518), .B(new_n537), .C1(new_n546), .C2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n524), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AOI22_X1  g349(.A1(new_n527), .A2(new_n529), .B1(new_n536), .B2(new_n533), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(new_n539), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n550), .A2(new_n552), .A3(KEYINPUT87), .ZN(new_n553));
  XNOR2_X1  g352(.A(G1gat), .B(G29gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(KEYINPUT0), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(G57gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(new_n221), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n542), .A2(new_n553), .A3(new_n558), .ZN(new_n559));
  XOR2_X1   g358(.A(KEYINPUT83), .B(KEYINPUT6), .Z(new_n560));
  AOI22_X1  g359(.A1(new_n548), .A2(new_n549), .B1(new_n551), .B2(new_n539), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n560), .B1(new_n561), .B2(new_n557), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n560), .ZN(new_n564));
  NOR3_X1   g363(.A1(new_n561), .A2(new_n557), .A3(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  XOR2_X1   g366(.A(KEYINPUT88), .B(KEYINPUT35), .Z(new_n568));
  NAND3_X1  g367(.A1(new_n516), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT89), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n561), .A2(new_n557), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n550), .A2(new_n552), .A3(new_n557), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(new_n564), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n572), .B1(new_n574), .B2(KEYINPUT84), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT84), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n562), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n565), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n431), .A2(new_n432), .A3(new_n515), .A4(new_n468), .ZN(new_n579));
  OAI21_X1  g378(.A(KEYINPUT35), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n516), .A2(new_n567), .A3(KEYINPUT89), .A4(new_n568), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n571), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n565), .B1(new_n559), .B2(new_n562), .ZN(new_n583));
  AND3_X1   g382(.A1(new_n461), .A2(new_n462), .A3(KEYINPUT37), .ZN(new_n584));
  AOI21_X1  g383(.A(KEYINPUT37), .B1(new_n461), .B2(new_n462), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n435), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(KEYINPUT38), .ZN(new_n587));
  OR2_X1    g386(.A1(new_n586), .A2(KEYINPUT38), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n583), .A2(new_n464), .A3(new_n587), .A4(new_n588), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n465), .A2(new_n467), .ZN(new_n590));
  AND2_X1   g389(.A1(new_n590), .A2(new_n559), .ZN(new_n591));
  OR3_X1    g390(.A1(new_n520), .A2(new_n522), .A3(new_n519), .ZN(new_n592));
  OAI211_X1 g391(.A(KEYINPUT39), .B(new_n592), .C1(new_n551), .C2(new_n518), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n536), .A2(new_n533), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n594), .B1(new_n546), .B2(new_n547), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT39), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n595), .A2(new_n596), .A3(new_n519), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT86), .ZN(new_n598));
  AND3_X1   g397(.A1(new_n597), .A2(new_n598), .A3(new_n557), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n598), .B1(new_n597), .B2(new_n557), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n593), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT40), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI211_X1 g402(.A(KEYINPUT40), .B(new_n593), .C1(new_n599), .C2(new_n600), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n591), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n589), .A2(new_n605), .A3(new_n515), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n431), .A2(new_n432), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT36), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n515), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n610), .B1(new_n578), .B2(new_n590), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n606), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n582), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT21), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n306), .B1(new_n614), .B2(new_n248), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT19), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT20), .ZN(new_n617));
  OR2_X1    g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n616), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G127gat), .B(G155gat), .ZN(new_n621));
  XOR2_X1   g420(.A(new_n621), .B(KEYINPUT96), .Z(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n622), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n618), .A2(new_n619), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n248), .A2(new_n614), .ZN(new_n626));
  XOR2_X1   g425(.A(G183gat), .B(G211gat), .Z(new_n627));
  NAND2_X1  g426(.A1(G231gat), .A2(G233gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n626), .B(new_n629), .ZN(new_n630));
  AND3_X1   g429(.A1(new_n623), .A2(new_n625), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n630), .B1(new_n623), .B2(new_n625), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(G190gat), .B(G218gat), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n261), .A2(new_n295), .A3(new_n308), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n257), .A2(new_n317), .A3(new_n258), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT99), .ZN(new_n638));
  NAND3_X1  g437(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n639));
  AND3_X1   g438(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n638), .B1(new_n637), .B2(new_n639), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n636), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(G134gat), .B(G162gat), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n643), .ZN(new_n647));
  OAI211_X1 g446(.A(new_n636), .B(new_n647), .C1(new_n640), .C2(new_n641), .ZN(new_n648));
  AND3_X1   g447(.A1(new_n644), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n646), .B1(new_n644), .B2(new_n648), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n635), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n644), .A2(new_n648), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(new_n645), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n644), .A2(new_n646), .A3(new_n648), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n653), .A2(new_n634), .A3(new_n654), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n651), .A2(new_n655), .ZN(new_n656));
  AND4_X1   g455(.A1(new_n336), .A2(new_n613), .A3(new_n633), .A4(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(new_n578), .ZN(new_n658));
  XOR2_X1   g457(.A(KEYINPUT103), .B(G1gat), .Z(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(G1324gat));
  INV_X1    g459(.A(KEYINPUT104), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT42), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n657), .A2(new_n590), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(G8gat), .ZN(new_n664));
  NOR2_X1   g463(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n657), .A2(new_n590), .A3(new_n666), .A4(new_n667), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n662), .B1(new_n664), .B2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n668), .A2(new_n662), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n661), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n671), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n669), .A2(new_n673), .A3(KEYINPUT104), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n672), .A2(new_n674), .ZN(G1325gat));
  INV_X1    g474(.A(new_n607), .ZN(new_n676));
  AOI21_X1  g475(.A(G15gat), .B1(new_n657), .B2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n609), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n678), .A2(G15gat), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n677), .B1(new_n657), .B2(new_n679), .ZN(G1326gat));
  NAND2_X1  g479(.A1(new_n657), .A2(new_n610), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT43), .B(G22gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(G1327gat));
  NAND2_X1  g482(.A1(new_n651), .A2(new_n655), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n613), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n578), .ZN(new_n686));
  INV_X1    g485(.A(new_n633), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n336), .A2(new_n687), .ZN(new_n688));
  NOR4_X1   g487(.A1(new_n685), .A2(G29gat), .A3(new_n686), .A4(new_n688), .ZN(new_n689));
  XOR2_X1   g488(.A(new_n689), .B(KEYINPUT45), .Z(new_n690));
  NAND2_X1  g489(.A1(new_n685), .A2(KEYINPUT44), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n656), .B1(new_n582), .B2(new_n612), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n688), .B1(new_n691), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(new_n578), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(G29gat), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n690), .A2(new_n697), .ZN(G1328gat));
  INV_X1    g497(.A(G36gat), .ZN(new_n699));
  INV_X1    g498(.A(new_n688), .ZN(new_n700));
  NAND4_X1  g499(.A1(new_n692), .A2(new_n699), .A3(new_n590), .A4(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT105), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n701), .B1(new_n702), .B2(KEYINPUT46), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(KEYINPUT46), .ZN(new_n704));
  XOR2_X1   g503(.A(new_n703), .B(new_n704), .Z(new_n705));
  NAND2_X1  g504(.A1(new_n695), .A2(new_n590), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n705), .B1(new_n699), .B2(new_n707), .ZN(G1329gat));
  INV_X1    g507(.A(KEYINPUT47), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n290), .B1(new_n695), .B2(new_n678), .ZN(new_n710));
  NOR4_X1   g509(.A1(new_n685), .A2(G43gat), .A3(new_n607), .A4(new_n688), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n709), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n695), .A2(KEYINPUT106), .A3(new_n678), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n693), .B1(new_n613), .B2(new_n684), .ZN(new_n714));
  AOI211_X1 g513(.A(KEYINPUT44), .B(new_n656), .C1(new_n582), .C2(new_n612), .ZN(new_n715));
  OAI211_X1 g514(.A(new_n678), .B(new_n700), .C1(new_n714), .C2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT106), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n713), .A2(new_n718), .A3(G43gat), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT107), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n711), .A2(new_n709), .ZN(new_n721));
  AND3_X1   g520(.A1(new_n719), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n720), .B1(new_n719), .B2(new_n721), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n712), .B1(new_n722), .B2(new_n723), .ZN(G1330gat));
  INV_X1    g523(.A(new_n289), .ZN(new_n725));
  NOR4_X1   g524(.A1(new_n685), .A2(new_n725), .A3(new_n515), .A4(new_n688), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n695), .A2(new_n610), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n726), .B1(new_n727), .B2(new_n725), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT48), .ZN(G1331gat));
  NAND3_X1  g528(.A1(new_n656), .A2(new_n633), .A3(new_n335), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n730), .B1(new_n582), .B2(new_n612), .ZN(new_n731));
  AND2_X1   g530(.A1(new_n731), .A2(new_n280), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(new_n578), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g533(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n732), .A2(new_n590), .A3(new_n735), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(KEYINPUT108), .ZN(new_n737));
  NOR2_X1   g536(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n738));
  XOR2_X1   g537(.A(new_n737), .B(new_n738), .Z(G1333gat));
  AOI21_X1  g538(.A(G71gat), .B1(new_n732), .B2(new_n676), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n609), .A2(new_n240), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n740), .B1(new_n732), .B2(new_n741), .ZN(new_n742));
  XOR2_X1   g541(.A(new_n742), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g542(.A1(new_n280), .A2(new_n610), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n731), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g546(.A1(new_n633), .A2(new_n334), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n749), .B1(new_n691), .B2(new_n694), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n750), .A2(KEYINPUT109), .A3(new_n578), .A4(new_n280), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT109), .ZN(new_n752));
  OAI211_X1 g551(.A(new_n280), .B(new_n748), .C1(new_n714), .C2(new_n715), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n752), .B1(new_n753), .B2(new_n686), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n751), .A2(new_n754), .A3(G85gat), .ZN(new_n755));
  AND4_X1   g554(.A1(KEYINPUT51), .A2(new_n613), .A3(new_n684), .A4(new_n748), .ZN(new_n756));
  AOI21_X1  g555(.A(KEYINPUT51), .B1(new_n692), .B2(new_n748), .ZN(new_n757));
  OAI21_X1  g556(.A(KEYINPUT110), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT51), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n759), .B1(new_n685), .B2(new_n749), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT110), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n758), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n763), .A2(new_n221), .A3(new_n578), .A4(new_n280), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n755), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(KEYINPUT111), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT111), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n755), .A2(new_n764), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n766), .A2(new_n768), .ZN(G1336gat));
  NAND3_X1  g568(.A1(new_n750), .A2(new_n280), .A3(new_n590), .ZN(new_n770));
  AOI21_X1  g569(.A(KEYINPUT52), .B1(new_n770), .B2(G92gat), .ZN(new_n771));
  INV_X1    g570(.A(new_n763), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n280), .A2(new_n222), .A3(new_n590), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n771), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n692), .A2(KEYINPUT51), .A3(new_n748), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n773), .B1(new_n760), .B2(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n776), .B1(new_n770), .B2(G92gat), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n774), .B1(new_n777), .B2(new_n778), .ZN(G1337gat));
  OAI21_X1  g578(.A(G99gat), .B1(new_n753), .B2(new_n609), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n761), .B1(new_n760), .B2(new_n775), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n757), .A2(KEYINPUT110), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n408), .B(new_n280), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n780), .B1(new_n783), .B2(new_n607), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(KEYINPUT112), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT112), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n786), .B(new_n780), .C1(new_n783), .C2(new_n607), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(new_n787), .ZN(G1338gat));
  OR3_X1    g587(.A1(new_n753), .A2(KEYINPUT114), .A3(new_n515), .ZN(new_n789));
  OAI21_X1  g588(.A(KEYINPUT114), .B1(new_n753), .B2(new_n515), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n789), .A2(G106gat), .A3(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n792));
  OR2_X1    g591(.A1(new_n792), .A2(KEYINPUT113), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n744), .A2(G106gat), .ZN(new_n794));
  AOI22_X1  g593(.A1(new_n763), .A2(new_n794), .B1(KEYINPUT113), .B2(new_n792), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n791), .A2(new_n793), .A3(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(G106gat), .B1(new_n753), .B2(new_n515), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n794), .B1(new_n756), .B2(new_n757), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(KEYINPUT53), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n796), .A2(new_n800), .ZN(G1339gat));
  NAND2_X1  g600(.A1(new_n318), .A2(new_n319), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n309), .A2(new_n310), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(new_n312), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n328), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  AND3_X1   g604(.A1(new_n314), .A2(KEYINPUT92), .A3(new_n322), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n322), .B1(new_n314), .B2(KEYINPUT92), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n806), .A2(new_n807), .A3(new_n320), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n805), .B1(new_n808), .B2(new_n332), .ZN(new_n809));
  OAI211_X1 g608(.A(new_n809), .B(new_n278), .C1(new_n275), .C2(new_n272), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(KEYINPUT116), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT116), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n276), .A2(new_n812), .A3(new_n278), .A4(new_n809), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n269), .B1(new_n274), .B2(KEYINPUT54), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n251), .A2(new_n260), .A3(new_n262), .ZN(new_n817));
  INV_X1    g616(.A(new_n273), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n819), .A2(KEYINPUT54), .A3(new_n263), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n816), .A2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT55), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n816), .A2(KEYINPUT55), .A3(new_n820), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n825), .A2(new_n334), .A3(new_n271), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(KEYINPUT117), .B1(new_n814), .B2(new_n827), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n825), .A2(new_n334), .A3(new_n271), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(new_n823), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT117), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n830), .A2(new_n831), .A3(new_n813), .A4(new_n811), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n828), .A2(new_n656), .A3(new_n832), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n825), .A2(new_n271), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n684), .A2(new_n834), .A3(new_n809), .A4(new_n823), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n633), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n730), .A2(new_n280), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(KEYINPUT115), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT115), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n839), .B1(new_n730), .B2(new_n280), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  OR2_X1    g640(.A1(new_n836), .A2(new_n841), .ZN(new_n842));
  AND3_X1   g641(.A1(new_n842), .A2(new_n578), .A3(new_n468), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n607), .A2(new_n610), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n845), .A2(new_n335), .ZN(new_n846));
  XOR2_X1   g645(.A(new_n846), .B(G113gat), .Z(G1340gat));
  NOR2_X1   g646(.A1(new_n845), .A2(new_n279), .ZN(new_n848));
  XNOR2_X1  g647(.A(new_n848), .B(new_n383), .ZN(G1341gat));
  NOR2_X1   g648(.A1(new_n845), .A2(new_n687), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n850), .B(new_n392), .ZN(G1342gat));
  AND2_X1   g650(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n845), .A2(new_n656), .A3(new_n852), .ZN(new_n853));
  NOR2_X1   g652(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n853), .B(new_n854), .ZN(G1343gat));
  INV_X1    g654(.A(new_n835), .ZN(new_n856));
  AND3_X1   g655(.A1(new_n819), .A2(KEYINPUT54), .A3(new_n263), .ZN(new_n857));
  OAI21_X1  g656(.A(KEYINPUT118), .B1(new_n857), .B2(new_n815), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT118), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n816), .A2(new_n859), .A3(new_n820), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n858), .A2(new_n822), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n829), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n684), .B1(new_n862), .B2(new_n810), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n856), .B1(new_n863), .B2(KEYINPUT119), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT119), .ZN(new_n865));
  INV_X1    g664(.A(new_n810), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n866), .B1(new_n829), .B2(new_n861), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n865), .B1(new_n867), .B2(new_n684), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n633), .B1(new_n864), .B2(new_n868), .ZN(new_n869));
  OAI211_X1 g668(.A(KEYINPUT57), .B(new_n610), .C1(new_n869), .C2(new_n841), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT120), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(KEYINPUT55), .B1(new_n821), .B2(KEYINPUT118), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n826), .B1(new_n873), .B2(new_n860), .ZN(new_n874));
  OAI211_X1 g673(.A(KEYINPUT119), .B(new_n656), .C1(new_n874), .C2(new_n866), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n868), .A2(new_n835), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n687), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n838), .A2(new_n840), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n879), .A2(KEYINPUT120), .A3(KEYINPUT57), .A4(new_n610), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n610), .B1(new_n836), .B2(new_n841), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT57), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n872), .A2(new_n880), .A3(new_n883), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n678), .A2(new_n686), .A3(new_n590), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n884), .A2(new_n334), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(G141gat), .ZN(new_n887));
  INV_X1    g686(.A(new_n881), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n888), .A2(new_n481), .A3(new_n334), .A4(new_n885), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(KEYINPUT58), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT58), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n887), .A2(new_n889), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n891), .A2(new_n893), .ZN(G1344gat));
  NOR2_X1   g693(.A1(new_n495), .A2(new_n496), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n678), .A2(new_n895), .A3(new_n744), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n843), .A2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT59), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n881), .A2(KEYINPUT57), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n834), .A2(new_n823), .ZN(new_n900));
  OR3_X1    g699(.A1(new_n900), .A2(new_n656), .A3(KEYINPUT121), .ZN(new_n901));
  OAI21_X1  g700(.A(KEYINPUT121), .B1(new_n900), .B2(new_n656), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n901), .A2(new_n809), .A3(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(new_n863), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n633), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  OAI211_X1 g704(.A(new_n882), .B(new_n610), .C1(new_n905), .C2(new_n837), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n899), .A2(new_n280), .A3(new_n885), .A4(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT122), .ZN(new_n908));
  OR2_X1    g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n483), .B1(new_n907), .B2(new_n908), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n898), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n884), .A2(new_n280), .A3(new_n885), .ZN(new_n912));
  AND3_X1   g711(.A1(new_n912), .A2(new_n898), .A3(new_n895), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n897), .B1(new_n911), .B2(new_n913), .ZN(G1345gat));
  NAND3_X1  g713(.A1(new_n884), .A2(new_n633), .A3(new_n885), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(G155gat), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n687), .A2(G155gat), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n888), .A2(new_n885), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT123), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n916), .A2(new_n918), .A3(KEYINPUT123), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(G1346gat));
  NAND3_X1  g722(.A1(new_n888), .A2(new_n684), .A3(new_n885), .ZN(new_n924));
  INV_X1    g723(.A(G162gat), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n884), .A2(new_n885), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n684), .A2(G162gat), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT124), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n929), .B(new_n930), .ZN(G1347gat));
  NAND2_X1  g730(.A1(new_n844), .A2(new_n590), .ZN(new_n932));
  INV_X1    g731(.A(new_n932), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n842), .B(new_n686), .C1(KEYINPUT125), .C2(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT125), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n932), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n937), .A2(new_n337), .A3(new_n334), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n842), .A2(new_n686), .A3(new_n933), .ZN(new_n939));
  OAI21_X1  g738(.A(G169gat), .B1(new_n939), .B2(new_n335), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n938), .A2(new_n940), .ZN(G1348gat));
  NOR3_X1   g740(.A1(new_n939), .A2(new_n266), .A3(new_n279), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n937), .A2(new_n280), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n942), .B1(new_n943), .B2(new_n266), .ZN(G1349gat));
  XNOR2_X1  g743(.A(KEYINPUT27), .B(G183gat), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n937), .A2(new_n633), .A3(new_n945), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n375), .B1(new_n939), .B2(new_n687), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(KEYINPUT60), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT60), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n946), .A2(new_n950), .A3(new_n947), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n949), .A2(new_n951), .ZN(G1350gat));
  OAI21_X1  g751(.A(G190gat), .B1(new_n939), .B2(new_n656), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n953), .A2(KEYINPUT126), .ZN(new_n954));
  OAI21_X1  g753(.A(KEYINPUT61), .B1(new_n953), .B2(KEYINPUT126), .ZN(new_n955));
  OR2_X1    g754(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n937), .A2(new_n346), .A3(new_n684), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n954), .A2(new_n955), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(G1351gat));
  NOR2_X1   g758(.A1(new_n678), .A2(new_n468), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(new_n686), .ZN(new_n961));
  NOR4_X1   g760(.A1(new_n881), .A2(G197gat), .A3(new_n335), .A4(new_n961), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n899), .A2(new_n906), .ZN(new_n963));
  INV_X1    g762(.A(new_n961), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n963), .A2(new_n334), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n962), .B1(new_n965), .B2(G197gat), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT127), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  AOI211_X1 g767(.A(KEYINPUT127), .B(new_n962), .C1(new_n965), .C2(G197gat), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n968), .A2(new_n969), .ZN(G1352gat));
  NOR3_X1   g769(.A1(new_n678), .A2(G204gat), .A3(new_n468), .ZN(new_n971));
  NAND4_X1  g770(.A1(new_n842), .A2(new_n686), .A3(new_n745), .A4(new_n971), .ZN(new_n972));
  XOR2_X1   g771(.A(new_n972), .B(KEYINPUT62), .Z(new_n973));
  AND3_X1   g772(.A1(new_n963), .A2(new_n280), .A3(new_n964), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n973), .B1(new_n974), .B2(new_n268), .ZN(G1353gat));
  NAND3_X1  g774(.A1(new_n963), .A2(new_n633), .A3(new_n964), .ZN(new_n976));
  AND3_X1   g775(.A1(new_n976), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n977));
  AOI21_X1  g776(.A(KEYINPUT63), .B1(new_n976), .B2(G211gat), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n888), .A2(new_n964), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n633), .A2(new_n439), .ZN(new_n980));
  OAI22_X1  g779(.A1(new_n977), .A2(new_n978), .B1(new_n979), .B2(new_n980), .ZN(G1354gat));
  NAND4_X1  g780(.A1(new_n963), .A2(G218gat), .A3(new_n684), .A4(new_n964), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n440), .B1(new_n979), .B2(new_n656), .ZN(new_n983));
  AND2_X1   g782(.A1(new_n982), .A2(new_n983), .ZN(G1355gat));
endmodule


