//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 1 1 0 0 0 1 0 1 0 1 0 1 1 1 0 0 0 1 0 0 1 1 1 1 0 0 1 0 0 1 1 1 0 1 1 0 0 0 0 1 0 1 1 0 1 1 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:22 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998;
  INV_X1    g000(.A(G119), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT67), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT67), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G119), .ZN(new_n190));
  AND3_X1   g004(.A1(new_n188), .A2(new_n190), .A3(G116), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT85), .B(KEYINPUT5), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n188), .A2(new_n190), .A3(G116), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n187), .A2(G116), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n195), .A2(new_n197), .A3(new_n192), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n194), .A2(new_n198), .A3(G113), .ZN(new_n199));
  XNOR2_X1  g013(.A(KEYINPUT67), .B(G119), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n196), .B1(new_n200), .B2(G116), .ZN(new_n201));
  INV_X1    g015(.A(G113), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT2), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT2), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G113), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  AOI21_X1  g020(.A(KEYINPUT68), .B1(new_n201), .B2(new_n206), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n195), .A2(new_n206), .A3(KEYINPUT68), .A4(new_n197), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n199), .B1(new_n207), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G104), .ZN(new_n211));
  NOR3_X1   g025(.A1(new_n211), .A2(KEYINPUT3), .A3(G107), .ZN(new_n212));
  AND2_X1   g026(.A1(KEYINPUT82), .A2(G104), .ZN(new_n213));
  NOR2_X1   g027(.A1(KEYINPUT82), .A2(G104), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n212), .B1(new_n215), .B2(G107), .ZN(new_n216));
  INV_X1    g030(.A(G107), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n217), .B1(new_n213), .B2(new_n214), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(KEYINPUT3), .ZN(new_n219));
  INV_X1    g033(.A(G101), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n216), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n218), .B1(G104), .B2(new_n217), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G101), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT86), .B1(new_n210), .B2(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n195), .A2(new_n197), .A3(new_n206), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n202), .B1(new_n191), .B2(new_n193), .ZN(new_n229));
  AOI22_X1  g043(.A1(new_n228), .A2(new_n208), .B1(new_n229), .B2(new_n198), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT86), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n230), .A2(new_n231), .A3(new_n221), .A4(new_n223), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n225), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT84), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n228), .A2(new_n208), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n195), .A2(new_n197), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n236), .A2(new_n203), .A3(new_n205), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n220), .B1(new_n216), .B2(new_n219), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT4), .ZN(new_n239));
  AOI22_X1  g053(.A1(new_n235), .A2(new_n237), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT3), .ZN(new_n241));
  OR2_X1    g055(.A1(KEYINPUT82), .A2(G104), .ZN(new_n242));
  NAND2_X1  g056(.A1(KEYINPUT82), .A2(G104), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n241), .B1(new_n244), .B2(new_n217), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n242), .A2(G107), .A3(new_n243), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n241), .A2(new_n217), .A3(G104), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(G101), .B1(new_n245), .B2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n249), .A2(KEYINPUT4), .A3(new_n221), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n234), .B1(new_n240), .B2(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n237), .B1(new_n207), .B2(new_n209), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n238), .A2(new_n239), .ZN(new_n253));
  AND4_X1   g067(.A1(new_n234), .A2(new_n252), .A3(new_n250), .A4(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n233), .B1(new_n251), .B2(new_n254), .ZN(new_n255));
  XNOR2_X1  g069(.A(G110), .B(G122), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  OAI211_X1 g072(.A(new_n233), .B(new_n256), .C1(new_n251), .C2(new_n254), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n258), .A2(KEYINPUT6), .A3(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT6), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n255), .A2(new_n261), .A3(new_n257), .ZN(new_n262));
  INV_X1    g076(.A(G128), .ZN(new_n263));
  INV_X1    g077(.A(G146), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G143), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n263), .B1(new_n265), .B2(KEYINPUT1), .ZN(new_n266));
  XNOR2_X1  g080(.A(G143), .B(G146), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n266), .B(new_n267), .ZN(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT0), .B(G128), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT64), .ZN(new_n271));
  INV_X1    g085(.A(G143), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G146), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n265), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n270), .A2(new_n271), .A3(new_n274), .ZN(new_n275));
  OAI21_X1  g089(.A(KEYINPUT64), .B1(new_n267), .B2(new_n269), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT65), .ZN(new_n277));
  NAND2_X1  g091(.A1(KEYINPUT0), .A2(G128), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n277), .B1(new_n274), .B2(new_n278), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n267), .A2(KEYINPUT65), .A3(KEYINPUT0), .A4(G128), .ZN(new_n280));
  AOI22_X1  g094(.A1(new_n275), .A2(new_n276), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  MUX2_X1   g095(.A(new_n268), .B(new_n281), .S(G125), .Z(new_n282));
  INV_X1    g096(.A(G953), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(G224), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n282), .B(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n260), .A2(new_n262), .A3(new_n285), .ZN(new_n286));
  AND2_X1   g100(.A1(new_n284), .A2(KEYINPUT7), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n282), .B(new_n287), .ZN(new_n288));
  XOR2_X1   g102(.A(new_n256), .B(KEYINPUT8), .Z(new_n289));
  INV_X1    g103(.A(KEYINPUT5), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n229), .B1(new_n290), .B2(new_n236), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n224), .B1(new_n235), .B2(new_n291), .ZN(new_n292));
  AOI211_X1 g106(.A(new_n289), .B(new_n292), .C1(new_n224), .C2(new_n230), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n288), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(G902), .B1(new_n294), .B2(new_n259), .ZN(new_n295));
  OAI21_X1  g109(.A(G210), .B1(G237), .B2(G902), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n286), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT87), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n286), .A2(new_n295), .ZN(new_n299));
  INV_X1    g113(.A(new_n296), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT87), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n286), .A2(new_n302), .A3(new_n295), .A4(new_n296), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n298), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  AND2_X1   g118(.A1(new_n283), .A2(G952), .ZN(new_n305));
  NAND2_X1  g119(.A1(G234), .A2(G237), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  AND3_X1   g122(.A1(new_n306), .A2(G902), .A3(G953), .ZN(new_n309));
  XNOR2_X1  g123(.A(KEYINPUT21), .B(G898), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n308), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(G214), .B1(G237), .B2(G902), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  AND2_X1   g128(.A1(new_n304), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G469), .ZN(new_n316));
  INV_X1    g130(.A(G902), .ZN(new_n317));
  XNOR2_X1  g131(.A(G110), .B(G140), .ZN(new_n318));
  INV_X1    g132(.A(G227), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n319), .A2(G953), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n318), .B(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n250), .A2(new_n281), .A3(new_n253), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n268), .A2(new_n221), .A3(new_n223), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT10), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n268), .A2(new_n221), .A3(new_n223), .A4(KEYINPUT10), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n323), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(KEYINPUT83), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT69), .ZN(new_n330));
  INV_X1    g144(.A(G131), .ZN(new_n331));
  INV_X1    g145(.A(G134), .ZN(new_n332));
  OAI21_X1  g146(.A(KEYINPUT11), .B1(new_n332), .B2(G137), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT11), .ZN(new_n334));
  INV_X1    g148(.A(G137), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n334), .A2(new_n335), .A3(G134), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(KEYINPUT66), .B1(new_n335), .B2(G134), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT66), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n339), .A2(new_n332), .A3(G137), .ZN(new_n340));
  AND4_X1   g154(.A1(new_n331), .A2(new_n337), .A3(new_n338), .A4(new_n340), .ZN(new_n341));
  AND2_X1   g155(.A1(new_n338), .A2(new_n340), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n331), .B1(new_n342), .B2(new_n337), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n330), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n337), .A2(new_n338), .A3(new_n340), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(G131), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n342), .A2(new_n331), .A3(new_n337), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n346), .A2(KEYINPUT69), .A3(new_n347), .ZN(new_n348));
  AND2_X1   g162(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT83), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n323), .A2(new_n350), .A3(new_n326), .A4(new_n327), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n329), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n344), .A2(new_n348), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n323), .A2(new_n353), .A3(new_n326), .A4(new_n327), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n322), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n268), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n224), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n324), .ZN(new_n358));
  AOI21_X1  g172(.A(KEYINPUT12), .B1(new_n358), .B2(new_n349), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n346), .A2(new_n347), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(KEYINPUT12), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n361), .B1(new_n357), .B2(new_n324), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n354), .A2(new_n322), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n316), .B(new_n317), .C1(new_n355), .C2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n364), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n352), .A2(new_n367), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n354), .B1(new_n359), .B2(new_n362), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n321), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n368), .A2(new_n370), .A3(G469), .ZN(new_n371));
  NAND2_X1  g185(.A1(G469), .A2(G902), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n366), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(KEYINPUT9), .B(G234), .ZN(new_n374));
  OAI21_X1  g188(.A(G221), .B1(new_n374), .B2(G902), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(G140), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(G125), .ZN(new_n378));
  INV_X1    g192(.A(G125), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G140), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n378), .A2(new_n380), .A3(KEYINPUT74), .ZN(new_n381));
  OR3_X1    g195(.A1(new_n379), .A2(KEYINPUT74), .A3(G140), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n381), .A2(new_n382), .A3(KEYINPUT16), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT16), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n378), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G146), .ZN(new_n387));
  NOR2_X1   g201(.A1(G237), .A2(G953), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n388), .A2(G143), .A3(G214), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(G143), .B1(new_n388), .B2(G214), .ZN(new_n391));
  OAI21_X1  g205(.A(G131), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n391), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(new_n331), .A3(new_n389), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT17), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n392), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n383), .A2(new_n264), .A3(new_n385), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n393), .A2(new_n389), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n398), .A2(KEYINPUT17), .A3(G131), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n387), .A2(new_n396), .A3(new_n397), .A4(new_n399), .ZN(new_n400));
  XOR2_X1   g214(.A(KEYINPUT89), .B(G104), .Z(new_n401));
  XNOR2_X1  g215(.A(G113), .B(G122), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n401), .B(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n381), .A2(new_n382), .A3(G146), .ZN(new_n405));
  AND2_X1   g219(.A1(new_n378), .A2(new_n380), .ZN(new_n406));
  AOI21_X1  g220(.A(KEYINPUT76), .B1(new_n406), .B2(new_n264), .ZN(new_n407));
  AND4_X1   g221(.A1(KEYINPUT76), .A2(new_n378), .A3(new_n380), .A4(new_n264), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n405), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(KEYINPUT18), .A2(G131), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n393), .A2(new_n389), .A3(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n398), .A2(KEYINPUT18), .A3(G131), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n409), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n400), .A2(new_n404), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(KEYINPUT90), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT90), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n400), .A2(new_n413), .A3(new_n416), .A4(new_n404), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT19), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n419), .B1(new_n381), .B2(new_n382), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n406), .A2(KEYINPUT19), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n264), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n392), .A2(new_n394), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n387), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n413), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(KEYINPUT88), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT88), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n424), .A2(new_n413), .A3(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n426), .A2(new_n403), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n418), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(KEYINPUT91), .ZN(new_n431));
  NOR2_X1   g245(.A1(G475), .A2(G902), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT91), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n418), .A2(new_n429), .A3(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n431), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  AND2_X1   g249(.A1(new_n432), .A2(KEYINPUT92), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n432), .A2(KEYINPUT92), .ZN(new_n437));
  NOR3_X1   g251(.A1(new_n436), .A2(new_n437), .A3(KEYINPUT20), .ZN(new_n438));
  AOI22_X1  g252(.A1(new_n435), .A2(KEYINPUT20), .B1(new_n430), .B2(new_n438), .ZN(new_n439));
  AND2_X1   g253(.A1(new_n400), .A2(new_n413), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n418), .B1(new_n404), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n317), .ZN(new_n442));
  AND2_X1   g256(.A1(new_n442), .A2(G475), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n439), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT13), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n446), .B1(new_n263), .B2(G143), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n272), .A2(KEYINPUT13), .A3(G128), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n263), .A2(G143), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n447), .A2(new_n448), .A3(KEYINPUT94), .A4(new_n449), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n450), .B(G134), .C1(KEYINPUT94), .C2(new_n448), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n263), .A2(G143), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n272), .A2(G128), .ZN(new_n453));
  OR3_X1    g267(.A1(new_n452), .A2(new_n453), .A3(G134), .ZN(new_n454));
  INV_X1    g268(.A(G122), .ZN(new_n455));
  OAI21_X1  g269(.A(KEYINPUT93), .B1(new_n455), .B2(G116), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT93), .ZN(new_n457));
  INV_X1    g271(.A(G116), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n457), .A2(new_n458), .A3(G122), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n455), .A2(G116), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n460), .A2(new_n217), .A3(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n217), .B1(new_n460), .B2(new_n461), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n451), .B(new_n454), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  OR2_X1    g279(.A1(new_n460), .A2(KEYINPUT14), .ZN(new_n466));
  AOI22_X1  g280(.A1(new_n460), .A2(KEYINPUT14), .B1(G116), .B2(new_n455), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n217), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(G134), .B1(new_n452), .B2(new_n453), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n454), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(new_n462), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n465), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(KEYINPUT95), .ZN(new_n473));
  INV_X1    g287(.A(G217), .ZN(new_n474));
  NOR3_X1   g288(.A1(new_n374), .A2(new_n474), .A3(G953), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT95), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n465), .B(new_n477), .C1(new_n468), .C2(new_n471), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n473), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n472), .A2(KEYINPUT95), .A3(new_n475), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n479), .A2(new_n317), .A3(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT96), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n479), .A2(KEYINPUT96), .A3(new_n317), .A4(new_n480), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT15), .ZN(new_n485));
  AOI22_X1  g299(.A1(new_n483), .A2(new_n484), .B1(new_n485), .B2(G478), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n484), .A2(new_n485), .A3(G478), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n445), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n315), .A2(new_n376), .A3(new_n490), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n332), .A2(G137), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n335), .A2(G134), .ZN(new_n493));
  OAI21_X1  g307(.A(G131), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AND2_X1   g308(.A1(new_n347), .A2(new_n494), .ZN(new_n495));
  AOI22_X1  g309(.A1(new_n281), .A2(new_n360), .B1(new_n495), .B2(new_n268), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n252), .B1(new_n496), .B2(KEYINPUT30), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n344), .A2(new_n281), .A3(new_n348), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n495), .A2(new_n268), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(KEYINPUT30), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(KEYINPUT70), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT70), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n498), .A2(new_n502), .A3(KEYINPUT30), .A4(new_n499), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n497), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n252), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n498), .A2(new_n505), .A3(new_n499), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n388), .A2(G210), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n509), .B(KEYINPUT27), .ZN(new_n510));
  XNOR2_X1  g324(.A(KEYINPUT26), .B(G101), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n510), .B(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n508), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n507), .A2(KEYINPUT28), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT28), .ZN(new_n516));
  OAI22_X1  g330(.A1(new_n506), .A2(new_n516), .B1(new_n505), .B2(new_n496), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n512), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(KEYINPUT29), .B1(new_n514), .B2(new_n518), .ZN(new_n519));
  OR3_X1    g333(.A1(new_n507), .A2(KEYINPUT72), .A3(KEYINPUT28), .ZN(new_n520));
  OAI21_X1  g334(.A(KEYINPUT72), .B1(new_n507), .B2(KEYINPUT28), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n505), .B1(new_n498), .B2(new_n499), .ZN(new_n522));
  OAI21_X1  g336(.A(KEYINPUT28), .B1(new_n507), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n520), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT29), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n513), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n317), .B1(new_n524), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(G472), .B1(new_n519), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g343(.A1(G472), .A2(G902), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n501), .A2(new_n503), .ZN(new_n532));
  INV_X1    g346(.A(new_n497), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT31), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n506), .A2(new_n512), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n534), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n513), .B1(new_n515), .B2(new_n517), .ZN(new_n539));
  OAI21_X1  g353(.A(KEYINPUT31), .B1(new_n504), .B2(new_n536), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT71), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n538), .A2(new_n540), .A3(KEYINPUT71), .A4(new_n539), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n531), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n529), .B1(new_n545), .B2(KEYINPUT32), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n543), .A2(new_n544), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT32), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n531), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(KEYINPUT73), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT73), .ZN(new_n551));
  INV_X1    g365(.A(new_n549), .ZN(new_n552));
  AOI211_X1 g366(.A(new_n551), .B(new_n552), .C1(new_n543), .C2(new_n544), .ZN(new_n553));
  NOR3_X1   g367(.A1(new_n546), .A2(new_n550), .A3(new_n553), .ZN(new_n554));
  OR2_X1    g368(.A1(new_n407), .A2(new_n408), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n387), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n187), .A2(new_n263), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n557), .B1(new_n200), .B2(new_n263), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(KEYINPUT24), .B(G110), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(G110), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT23), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n563), .B1(new_n200), .B2(G128), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n562), .B(new_n564), .C1(new_n558), .C2(new_n563), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT75), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n561), .A2(new_n565), .A3(KEYINPUT75), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n556), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n564), .B1(new_n558), .B2(new_n563), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(G110), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n573), .B1(new_n560), .B2(new_n559), .ZN(new_n574));
  AND2_X1   g388(.A1(new_n387), .A2(new_n397), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(KEYINPUT22), .B(G137), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n283), .A2(G221), .A3(G234), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n578), .B(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n571), .A2(new_n577), .A3(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n580), .B(KEYINPUT77), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n582), .B1(new_n570), .B2(new_n576), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT78), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT25), .ZN(new_n585));
  AOI21_X1  g399(.A(G902), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n581), .A2(new_n583), .A3(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n584), .A2(new_n585), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n588), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n581), .A2(new_n583), .A3(new_n590), .A4(new_n586), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n474), .B1(G234), .B2(new_n317), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n589), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(KEYINPUT79), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT79), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n589), .A2(new_n595), .A3(new_n591), .A4(new_n592), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n592), .A2(G902), .ZN(new_n597));
  XOR2_X1   g411(.A(new_n597), .B(KEYINPUT80), .Z(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n581), .A2(new_n583), .A3(new_n599), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n594), .A2(new_n596), .A3(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g416(.A(KEYINPUT81), .B1(new_n554), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n550), .A2(new_n553), .ZN(new_n604));
  INV_X1    g418(.A(G472), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n514), .A2(new_n518), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(new_n525), .ZN(new_n607));
  INV_X1    g421(.A(new_n528), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n605), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n547), .A2(new_n530), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n609), .B1(new_n610), .B2(new_n548), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n604), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT81), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n612), .A2(new_n613), .A3(new_n601), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n491), .B1(new_n603), .B2(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(new_n220), .ZN(G3));
  AOI21_X1  g430(.A(G902), .B1(new_n543), .B2(new_n544), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n545), .B1(new_n618), .B2(G472), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n619), .A2(KEYINPUT97), .A3(new_n601), .A4(new_n376), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT97), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n610), .B1(new_n605), .B2(new_n617), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n376), .A2(new_n601), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(KEYINPUT33), .B1(new_n479), .B2(new_n480), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT98), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n472), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(new_n475), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n627), .B1(KEYINPUT33), .B2(new_n630), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n317), .A2(G478), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n481), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n635), .A2(G478), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n443), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n430), .A2(new_n438), .ZN(new_n639));
  INV_X1    g453(.A(new_n434), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n433), .B1(new_n418), .B2(new_n429), .ZN(new_n641));
  INV_X1    g455(.A(new_n432), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT20), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n639), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n637), .B1(new_n638), .B2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n301), .A2(new_n297), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n312), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n647), .A2(new_n649), .A3(new_n311), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n626), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT99), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT34), .B(G104), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G6));
  XNOR2_X1  g468(.A(new_n435), .B(KEYINPUT20), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n655), .A2(new_n638), .A3(new_n489), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n649), .A2(new_n656), .A3(new_n311), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n626), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT35), .B(G107), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G9));
  NAND2_X1  g474(.A1(new_n571), .A2(new_n577), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n582), .A2(KEYINPUT36), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n599), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n594), .A2(new_n596), .A3(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n622), .A2(new_n666), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n667), .A2(new_n315), .A3(new_n376), .A4(new_n490), .ZN(new_n668));
  XOR2_X1   g482(.A(KEYINPUT37), .B(G110), .Z(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G12));
  NAND3_X1  g484(.A1(new_n665), .A2(new_n375), .A3(new_n373), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n649), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n283), .A2(G900), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n673), .A2(G902), .A3(new_n306), .ZN(new_n674));
  OR2_X1    g488(.A1(new_n674), .A2(KEYINPUT100), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(KEYINPUT100), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n675), .A2(new_n307), .A3(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n656), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n547), .A2(new_n549), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n551), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n547), .A2(KEYINPUT73), .A3(new_n549), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  OAI211_X1 g497(.A(new_n672), .B(new_n679), .C1(new_n683), .C2(new_n546), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G128), .ZN(G30));
  XOR2_X1   g499(.A(KEYINPUT101), .B(KEYINPUT39), .Z(new_n686));
  XNOR2_X1  g500(.A(new_n677), .B(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n376), .A2(new_n687), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n688), .A2(KEYINPUT40), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n688), .A2(KEYINPUT40), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n312), .B1(new_n486), .B2(new_n487), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n691), .B1(new_n645), .B2(new_n638), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n689), .A2(new_n690), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n304), .B(KEYINPUT38), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n610), .A2(new_n548), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n508), .A2(new_n513), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n507), .A2(new_n522), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n317), .B1(new_n699), .B2(new_n512), .ZN(new_n700));
  OAI21_X1  g514(.A(G472), .B1(new_n697), .B2(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n604), .A2(new_n696), .A3(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n694), .A2(new_n666), .A3(new_n695), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G143), .ZN(G45));
  NAND2_X1  g518(.A1(new_n646), .A2(new_n677), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  OAI211_X1 g520(.A(new_n672), .B(new_n706), .C1(new_n683), .C2(new_n546), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G146), .ZN(G48));
  AOI21_X1  g522(.A(new_n602), .B1(new_n604), .B2(new_n611), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n317), .B1(new_n355), .B2(new_n365), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(G469), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n711), .A2(new_n375), .A3(new_n366), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n709), .A2(new_n650), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(KEYINPUT41), .B(G113), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(KEYINPUT102), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n714), .B(new_n716), .ZN(G15));
  NAND4_X1  g531(.A1(new_n612), .A2(new_n601), .A3(new_n657), .A4(new_n713), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G116), .ZN(G18));
  INV_X1    g533(.A(new_n311), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n665), .A2(new_n444), .A3(new_n720), .A4(new_n488), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n721), .A2(new_n649), .A3(new_n712), .ZN(new_n722));
  AND2_X1   g536(.A1(new_n612), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(new_n187), .ZN(G21));
  AND2_X1   g538(.A1(new_n524), .A2(new_n513), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n538), .A2(new_n540), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n530), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  OAI211_X1 g541(.A(new_n601), .B(new_n727), .C1(new_n617), .C2(new_n605), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  AND4_X1   g543(.A1(new_n720), .A2(new_n692), .A3(new_n713), .A4(new_n648), .ZN(new_n730));
  AND2_X1   g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(new_n455), .ZN(G24));
  OAI211_X1 g546(.A(new_n727), .B(new_n665), .C1(new_n617), .C2(new_n605), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n733), .A2(new_n705), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n649), .A2(new_n712), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G125), .ZN(G27));
  NAND2_X1  g551(.A1(new_n696), .A2(new_n680), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(KEYINPUT106), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT106), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n696), .A2(new_n740), .A3(new_n680), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n739), .A2(new_n529), .A3(new_n741), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n298), .A2(new_n303), .ZN(new_n743));
  INV_X1    g557(.A(new_n375), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n366), .A2(new_n372), .ZN(new_n745));
  AOI22_X1  g559(.A1(new_n367), .A2(new_n352), .B1(new_n369), .B2(new_n321), .ZN(new_n746));
  AOI21_X1  g560(.A(KEYINPUT103), .B1(new_n746), .B2(G469), .ZN(new_n747));
  AND4_X1   g561(.A1(KEYINPUT103), .A2(new_n368), .A3(G469), .A4(new_n370), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n744), .B1(new_n745), .B2(new_n749), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n313), .B1(new_n299), .B2(new_n300), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n743), .A2(KEYINPUT104), .A3(new_n750), .A4(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT104), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n298), .A2(new_n301), .A3(new_n303), .A4(new_n312), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT103), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n371), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n746), .A2(KEYINPUT103), .A3(G469), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n756), .A2(new_n366), .A3(new_n757), .A4(new_n372), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n375), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n753), .B1(new_n754), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n752), .A2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT42), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n705), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n742), .A2(new_n601), .A3(new_n761), .A4(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n761), .A2(new_n612), .A3(new_n601), .A4(new_n706), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n765), .A2(KEYINPUT105), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT105), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n709), .A2(new_n761), .A3(new_n767), .A4(new_n706), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n762), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n764), .B1(new_n766), .B2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G131), .ZN(G33));
  NAND3_X1  g585(.A1(new_n709), .A2(new_n679), .A3(new_n761), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G134), .ZN(G36));
  INV_X1    g587(.A(new_n637), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n444), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(KEYINPUT43), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT107), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n622), .A2(new_n665), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(KEYINPUT108), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT44), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n778), .A2(KEYINPUT44), .A3(new_n780), .ZN(new_n784));
  INV_X1    g598(.A(new_n366), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n746), .A2(KEYINPUT45), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n746), .A2(KEYINPUT45), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n786), .A2(G469), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(new_n372), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT46), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n785), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n791), .B1(new_n790), .B2(new_n789), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(new_n375), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n751), .A2(new_n298), .A3(new_n303), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n794), .A2(new_n687), .A3(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n783), .A2(new_n784), .A3(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G137), .ZN(G39));
  XNOR2_X1  g612(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n793), .B(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n554), .A2(new_n602), .A3(new_n706), .A4(new_n795), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(new_n377), .ZN(G42));
  NOR2_X1   g618(.A1(new_n702), .A2(new_n602), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n754), .A2(new_n307), .A3(new_n712), .ZN(new_n806));
  AND4_X1   g620(.A1(new_n444), .A2(new_n805), .A3(new_n637), .A4(new_n806), .ZN(new_n807));
  XOR2_X1   g621(.A(new_n807), .B(KEYINPUT115), .Z(new_n808));
  NOR3_X1   g622(.A1(new_n776), .A2(new_n307), .A3(new_n728), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n695), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT114), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT50), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n811), .A2(new_n313), .A3(new_n713), .A4(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n810), .A2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n812), .A2(new_n813), .ZN(new_n818));
  INV_X1    g632(.A(new_n733), .ZN(new_n819));
  INV_X1    g633(.A(new_n776), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n820), .A2(new_n806), .ZN(new_n821));
  AOI22_X1  g635(.A1(new_n817), .A2(new_n818), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n711), .A2(new_n366), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n801), .B1(new_n375), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n810), .A2(new_n754), .ZN(new_n825));
  INV_X1    g639(.A(new_n818), .ZN(new_n826));
  AOI22_X1  g640(.A1(new_n824), .A2(new_n825), .B1(new_n816), .B2(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n808), .A2(new_n822), .A3(new_n827), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(KEYINPUT51), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n742), .A2(new_n601), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(new_n821), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(KEYINPUT48), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n805), .A2(new_n646), .A3(new_n806), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n809), .A2(new_n735), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n832), .A2(new_n305), .A3(new_n833), .A4(new_n834), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n835), .B(KEYINPUT116), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n829), .A2(new_n836), .ZN(new_n837));
  AOI22_X1  g651(.A1(new_n612), .A2(new_n722), .B1(new_n729), .B2(new_n730), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n714), .A2(new_n838), .A3(new_n668), .A4(new_n718), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n304), .A2(new_n646), .A3(new_n314), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n840), .A2(KEYINPUT111), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n304), .A2(new_n314), .A3(new_n444), .A4(new_n489), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n842), .B1(new_n840), .B2(KEYINPUT111), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n844), .A2(new_n625), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n839), .A2(new_n615), .A3(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT112), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n709), .A2(new_n679), .A3(new_n761), .ZN(new_n848));
  AOI21_X1  g662(.A(KEYINPUT104), .B1(new_n795), .B2(new_n750), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n754), .A2(new_n753), .A3(new_n759), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n734), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n655), .A2(new_n638), .A3(new_n488), .A4(new_n677), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n671), .A2(new_n852), .A3(new_n754), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n612), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n847), .B1(new_n848), .B2(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n772), .A2(KEYINPUT112), .A3(new_n851), .A4(new_n854), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n846), .A2(new_n858), .A3(new_n770), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n692), .A2(new_n648), .A3(new_n677), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n861), .A2(new_n759), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n696), .A2(new_n701), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n862), .B(new_n666), .C1(new_n683), .C2(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n864), .A2(new_n684), .A3(new_n707), .A4(new_n736), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT52), .ZN(new_n866));
  AOI21_X1  g680(.A(KEYINPUT113), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n612), .B(new_n672), .C1(new_n679), .C2(new_n706), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n868), .A2(KEYINPUT52), .A3(new_n736), .A4(new_n864), .ZN(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n867), .B(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n860), .A2(new_n871), .A3(KEYINPUT53), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT54), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n865), .A2(new_n866), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(new_n869), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n846), .A2(new_n858), .A3(new_n770), .A4(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT53), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n872), .A2(new_n873), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT53), .B1(new_n860), .B2(new_n871), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n876), .A2(new_n877), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n879), .B1(new_n882), .B2(new_n873), .ZN(new_n883));
  OAI22_X1  g697(.A1(new_n837), .A2(new_n883), .B1(G952), .B2(G953), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n823), .A2(KEYINPUT49), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(KEYINPUT110), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n444), .A2(new_n774), .A3(new_n312), .A4(new_n375), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n887), .B1(KEYINPUT49), .B2(new_n823), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n805), .A2(new_n811), .A3(new_n886), .A4(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n884), .A2(new_n889), .ZN(G75));
  NOR2_X1   g704(.A1(new_n283), .A2(G952), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n317), .B1(new_n872), .B2(new_n878), .ZN(new_n893));
  AOI21_X1  g707(.A(KEYINPUT56), .B1(new_n893), .B2(G210), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n285), .B(KEYINPUT118), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n895), .B(KEYINPUT55), .Z(new_n896));
  NAND2_X1  g710(.A1(new_n260), .A2(new_n262), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT117), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n896), .B(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n892), .B1(new_n894), .B2(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n901), .B1(new_n894), .B2(new_n900), .ZN(G51));
  XOR2_X1   g716(.A(new_n372), .B(KEYINPUT57), .Z(new_n903));
  NAND2_X1  g717(.A1(new_n872), .A2(new_n878), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n904), .A2(KEYINPUT54), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n873), .B1(new_n872), .B2(new_n878), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n903), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OR2_X1    g721(.A1(new_n355), .A2(new_n365), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n893), .A2(G469), .A3(new_n787), .A4(new_n786), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n891), .B1(new_n909), .B2(new_n910), .ZN(G54));
  NAND3_X1  g725(.A1(new_n893), .A2(KEYINPUT58), .A3(G475), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n640), .A2(new_n641), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n912), .A2(new_n914), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n915), .A2(new_n916), .A3(new_n891), .ZN(G60));
  NOR2_X1   g731(.A1(new_n905), .A2(new_n906), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n631), .B(KEYINPUT119), .ZN(new_n919));
  NAND2_X1  g733(.A1(G478), .A2(G902), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT59), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n892), .B1(new_n918), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n919), .B1(new_n883), .B2(new_n921), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n923), .A2(new_n924), .ZN(G63));
  NAND2_X1  g739(.A1(G217), .A2(G902), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT60), .Z(new_n927));
  NOR2_X1   g741(.A1(new_n867), .A2(new_n870), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n865), .A2(KEYINPUT113), .A3(new_n866), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n930), .A2(new_n859), .A3(new_n877), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n876), .A2(new_n877), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n927), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n581), .A2(new_n583), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n891), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT121), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n904), .A2(new_n936), .A3(new_n663), .A4(new_n927), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n663), .B(new_n927), .C1(new_n931), .C2(new_n932), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(KEYINPUT121), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n935), .A2(new_n937), .A3(new_n939), .ZN(new_n940));
  XNOR2_X1  g754(.A(KEYINPUT120), .B(KEYINPUT61), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n935), .A2(KEYINPUT61), .A3(new_n938), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(G66));
  INV_X1    g758(.A(new_n310), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n283), .B1(new_n945), .B2(G224), .ZN(new_n946));
  INV_X1    g760(.A(new_n846), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n946), .B1(new_n947), .B2(new_n283), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n898), .B1(G898), .B2(new_n283), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT122), .Z(new_n950));
  XNOR2_X1  g764(.A(new_n948), .B(new_n950), .ZN(G69));
  OAI21_X1  g765(.A(new_n532), .B1(KEYINPUT30), .B2(new_n496), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n420), .A2(new_n421), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n952), .B(new_n953), .Z(new_n954));
  NAND2_X1  g768(.A1(new_n603), .A2(new_n614), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n646), .B1(new_n444), .B2(new_n489), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n956), .A2(new_n688), .A3(new_n754), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n803), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n868), .A2(new_n736), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n703), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(KEYINPUT62), .ZN(new_n961));
  AND3_X1   g775(.A1(new_n958), .A2(new_n797), .A3(new_n961), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n960), .A2(KEYINPUT62), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n963), .B(KEYINPUT124), .ZN(new_n964));
  AOI21_X1  g778(.A(G953), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT123), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n954), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n962), .A2(new_n964), .ZN(new_n968));
  AOI21_X1  g782(.A(KEYINPUT123), .B1(new_n968), .B2(new_n283), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n692), .A2(new_n648), .ZN(new_n970));
  AND3_X1   g784(.A1(new_n794), .A2(new_n687), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n830), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT125), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n971), .A2(new_n830), .A3(KEYINPUT125), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n803), .A2(new_n848), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n976), .A2(new_n797), .A3(new_n959), .A4(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n770), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n283), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n954), .A2(new_n673), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n967), .B1(new_n969), .B2(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n673), .B1(new_n319), .B2(G953), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(new_n984), .ZN(new_n986));
  OAI211_X1 g800(.A(new_n967), .B(new_n986), .C1(new_n969), .C2(new_n982), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n985), .A2(new_n987), .ZN(G72));
  NOR2_X1   g802(.A1(new_n968), .A2(new_n947), .ZN(new_n989));
  NAND2_X1  g803(.A1(G472), .A2(G902), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT63), .Z(new_n991));
  XNOR2_X1  g805(.A(new_n991), .B(KEYINPUT126), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n697), .B1(new_n989), .B2(new_n992), .ZN(new_n993));
  NOR3_X1   g807(.A1(new_n978), .A2(new_n979), .A3(new_n947), .ZN(new_n994));
  OAI211_X1 g808(.A(new_n513), .B(new_n508), .C1(new_n994), .C2(new_n992), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n993), .A2(new_n892), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n514), .A2(new_n991), .ZN(new_n997));
  NOR3_X1   g811(.A1(new_n882), .A2(new_n697), .A3(new_n997), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n996), .A2(new_n998), .ZN(G57));
endmodule


