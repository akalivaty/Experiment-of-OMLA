

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781;

  AND2_X1 U379 ( .A1(n395), .A2(n394), .ZN(n393) );
  NAND2_X1 U380 ( .A1(n422), .A2(n416), .ZN(n396) );
  XNOR2_X1 U381 ( .A(n357), .B(n462), .ZN(n761) );
  XNOR2_X1 U382 ( .A(n460), .B(n511), .ZN(n357) );
  XNOR2_X2 U383 ( .A(n577), .B(n404), .ZN(n603) );
  NAND2_X2 U384 ( .A1(n549), .A2(n528), .ZN(n529) );
  XNOR2_X2 U385 ( .A(n591), .B(n457), .ZN(n576) );
  XNOR2_X2 U386 ( .A(G902), .B(KEYINPUT15), .ZN(n634) );
  XNOR2_X2 U387 ( .A(n405), .B(n360), .ZN(n539) );
  AND2_X2 U388 ( .A1(n374), .A2(n373), .ZN(n372) );
  AND2_X2 U389 ( .A1(n530), .A2(n668), .ZN(n379) );
  NOR2_X1 U390 ( .A1(n703), .A2(n702), .ZN(n444) );
  XNOR2_X1 U391 ( .A(n551), .B(n550), .ZN(n660) );
  XNOR2_X1 U392 ( .A(n427), .B(G125), .ZN(n464) );
  XNOR2_X1 U393 ( .A(n387), .B(G137), .ZN(n402) );
  XNOR2_X2 U394 ( .A(n765), .B(G146), .ZN(n453) );
  BUF_X1 U395 ( .A(n453), .Z(n358) );
  OR2_X2 U396 ( .A1(n746), .A2(G902), .ZN(n405) );
  XNOR2_X1 U397 ( .A(n464), .B(n428), .ZN(n491) );
  NAND2_X1 U398 ( .A1(n420), .A2(n634), .ZN(n419) );
  INV_X1 U399 ( .A(n477), .ZN(n420) );
  NOR2_X1 U400 ( .A1(G953), .A2(G237), .ZN(n492) );
  XNOR2_X1 U401 ( .A(n383), .B(KEYINPUT66), .ZN(n563) );
  INV_X1 U402 ( .A(G237), .ZN(n473) );
  INV_X1 U403 ( .A(G902), .ZN(n474) );
  XNOR2_X1 U404 ( .A(G119), .B(G137), .ZN(n431) );
  XNOR2_X1 U405 ( .A(n398), .B(n397), .ZN(n508) );
  INV_X1 U406 ( .A(KEYINPUT8), .ZN(n397) );
  XOR2_X1 U407 ( .A(n491), .B(n490), .Z(n767) );
  INV_X1 U408 ( .A(G146), .ZN(n427) );
  NOR2_X1 U409 ( .A1(n541), .A2(n368), .ZN(n370) );
  NAND2_X1 U410 ( .A1(n390), .A2(n389), .ZN(n391) );
  XNOR2_X1 U411 ( .A(n539), .B(KEYINPUT1), .ZN(n703) );
  XNOR2_X1 U412 ( .A(n438), .B(n437), .ZN(n527) );
  NOR2_X1 U413 ( .A1(n642), .A2(G902), .ZN(n438) );
  XNOR2_X1 U414 ( .A(n411), .B(G104), .ZN(n461) );
  INV_X1 U415 ( .A(G110), .ZN(n411) );
  NAND2_X1 U416 ( .A1(n472), .A2(KEYINPUT2), .ZN(n635) );
  OR2_X2 U417 ( .A1(n700), .A2(n359), .ZN(n403) );
  XNOR2_X1 U418 ( .A(n621), .B(n380), .ZN(n579) );
  INV_X1 U419 ( .A(KEYINPUT107), .ZN(n380) );
  OR2_X1 U420 ( .A1(n722), .A2(n705), .ZN(n424) );
  BUF_X1 U421 ( .A(n527), .Z(n706) );
  INV_X2 U422 ( .A(G953), .ZN(n776) );
  AND2_X1 U423 ( .A1(n378), .A2(n403), .ZN(n751) );
  XNOR2_X1 U424 ( .A(n453), .B(n399), .ZN(n746) );
  XNOR2_X1 U425 ( .A(n401), .B(n400), .ZN(n399) );
  XNOR2_X1 U426 ( .A(n365), .B(n410), .ZN(n400) );
  XNOR2_X1 U427 ( .A(n490), .B(n461), .ZN(n401) );
  NOR2_X1 U428 ( .A1(n553), .A2(n660), .ZN(n552) );
  NAND2_X1 U429 ( .A1(n385), .A2(n384), .ZN(n383) );
  NAND2_X1 U430 ( .A1(G234), .A2(G237), .ZN(n479) );
  NOR2_X1 U431 ( .A1(n417), .A2(n423), .ZN(n416) );
  INV_X1 U432 ( .A(n718), .ZN(n423) );
  AND2_X1 U433 ( .A1(n418), .A2(n392), .ZN(n389) );
  INV_X1 U434 ( .A(KEYINPUT83), .ZN(n392) );
  XNOR2_X1 U435 ( .A(G116), .B(G131), .ZN(n449) );
  XOR2_X1 U436 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n494) );
  XNOR2_X1 U437 ( .A(G113), .B(G143), .ZN(n496) );
  XOR2_X1 U438 ( .A(KEYINPUT95), .B(KEYINPUT97), .Z(n497) );
  XNOR2_X1 U439 ( .A(G122), .B(G104), .ZN(n498) );
  INV_X1 U440 ( .A(KEYINPUT73), .ZN(n631) );
  XNOR2_X1 U441 ( .A(n387), .B(n463), .ZN(n465) );
  XNOR2_X1 U442 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n463) );
  XNOR2_X1 U443 ( .A(n566), .B(KEYINPUT64), .ZN(n567) );
  INV_X1 U444 ( .A(KEYINPUT48), .ZN(n619) );
  XNOR2_X1 U445 ( .A(n444), .B(n443), .ZN(n536) );
  NAND2_X1 U446 ( .A1(n477), .A2(n472), .ZN(n421) );
  XNOR2_X1 U447 ( .A(n435), .B(n434), .ZN(n642) );
  XNOR2_X1 U448 ( .A(n429), .B(n491), .ZN(n435) );
  XOR2_X1 U449 ( .A(G131), .B(G140), .Z(n490) );
  NAND2_X1 U450 ( .A1(n776), .A2(G227), .ZN(n410) );
  XNOR2_X1 U451 ( .A(n598), .B(n597), .ZN(n628) );
  INV_X1 U452 ( .A(KEYINPUT39), .ZN(n597) );
  NAND2_X1 U453 ( .A1(n376), .A2(n518), .ZN(n375) );
  NAND2_X1 U454 ( .A1(n372), .A2(n371), .ZN(n376) );
  INV_X1 U455 ( .A(KEYINPUT19), .ZN(n404) );
  XNOR2_X1 U456 ( .A(n503), .B(n382), .ZN(n543) );
  XNOR2_X1 U457 ( .A(n504), .B(n505), .ZN(n382) );
  AND2_X1 U458 ( .A1(n403), .A2(G472), .ZN(n409) );
  XNOR2_X1 U459 ( .A(n671), .B(n670), .ZN(n672) );
  AND2_X1 U460 ( .A1(n403), .A2(G217), .ZN(n406) );
  XNOR2_X1 U461 ( .A(n642), .B(KEYINPUT121), .ZN(n643) );
  XNOR2_X1 U462 ( .A(n661), .B(KEYINPUT59), .ZN(n662) );
  AND2_X1 U463 ( .A1(n403), .A2(G475), .ZN(n407) );
  AND2_X1 U464 ( .A1(n403), .A2(G210), .ZN(n408) );
  XOR2_X1 U465 ( .A(KEYINPUT86), .B(n645), .Z(n749) );
  XNOR2_X1 U466 ( .A(n580), .B(n381), .ZN(n581) );
  XNOR2_X1 U467 ( .A(KEYINPUT108), .B(KEYINPUT36), .ZN(n381) );
  AND2_X1 U468 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U469 ( .A(n754), .B(n753), .ZN(n386) );
  XNOR2_X1 U470 ( .A(n748), .B(n747), .ZN(n750) );
  OR2_X1 U471 ( .A1(n641), .A2(n640), .ZN(n359) );
  XOR2_X1 U472 ( .A(n426), .B(n425), .Z(n360) );
  AND2_X1 U473 ( .A1(G217), .A2(n439), .ZN(n361) );
  XOR2_X1 U474 ( .A(G140), .B(KEYINPUT91), .Z(n362) );
  XOR2_X1 U475 ( .A(G110), .B(G128), .Z(n363) );
  XOR2_X1 U476 ( .A(n486), .B(n485), .Z(n364) );
  NAND2_X2 U477 ( .A1(n393), .A2(n391), .ZN(n577) );
  XOR2_X1 U478 ( .A(G101), .B(G107), .Z(n365) );
  AND2_X1 U479 ( .A1(n418), .A2(n421), .ZN(n366) );
  AND2_X1 U480 ( .A1(n403), .A2(KEYINPUT2), .ZN(n367) );
  XNOR2_X1 U481 ( .A(KEYINPUT75), .B(KEYINPUT34), .ZN(n368) );
  NAND2_X1 U482 ( .A1(n370), .A2(n369), .ZN(n371) );
  INV_X1 U483 ( .A(n717), .ZN(n369) );
  NAND2_X1 U484 ( .A1(n541), .A2(n368), .ZN(n373) );
  NAND2_X1 U485 ( .A1(n717), .A2(n368), .ZN(n374) );
  XNOR2_X2 U486 ( .A(n375), .B(KEYINPUT35), .ZN(n560) );
  XNOR2_X1 U487 ( .A(n620), .B(n619), .ZN(n641) );
  INV_X1 U488 ( .A(n418), .ZN(n388) );
  XNOR2_X1 U489 ( .A(n651), .B(n650), .ZN(n652) );
  OR2_X1 U490 ( .A1(n649), .A2(n419), .ZN(n418) );
  XNOR2_X1 U491 ( .A(n761), .B(n471), .ZN(n649) );
  INV_X1 U492 ( .A(n622), .ZN(n377) );
  NAND2_X1 U493 ( .A1(n633), .A2(n632), .ZN(n636) );
  NAND2_X2 U494 ( .A1(n636), .A2(n635), .ZN(n378) );
  NAND2_X1 U495 ( .A1(n406), .A2(n378), .ZN(n644) );
  NAND2_X1 U496 ( .A1(n407), .A2(n378), .ZN(n663) );
  NAND2_X1 U497 ( .A1(n408), .A2(n378), .ZN(n653) );
  NAND2_X1 U498 ( .A1(n409), .A2(n378), .ZN(n673) );
  XNOR2_X2 U499 ( .A(n459), .B(n458), .ZN(n717) );
  NAND2_X1 U500 ( .A1(n379), .A2(n552), .ZN(n558) );
  NAND2_X1 U501 ( .A1(n575), .A2(n576), .ZN(n621) );
  INV_X1 U502 ( .A(KEYINPUT44), .ZN(n384) );
  INV_X1 U503 ( .A(n669), .ZN(n385) );
  NOR2_X1 U504 ( .A1(n386), .A2(n755), .ZN(G63) );
  XNOR2_X2 U505 ( .A(KEYINPUT68), .B(KEYINPUT4), .ZN(n387) );
  NAND2_X1 U506 ( .A1(n388), .A2(KEYINPUT83), .ZN(n394) );
  INV_X1 U507 ( .A(n396), .ZN(n390) );
  NAND2_X1 U508 ( .A1(n396), .A2(KEYINPUT83), .ZN(n395) );
  NAND2_X1 U509 ( .A1(n776), .A2(G234), .ZN(n398) );
  XNOR2_X2 U510 ( .A(n512), .B(n402), .ZN(n765) );
  XNOR2_X2 U511 ( .A(n467), .B(G134), .ZN(n512) );
  OR2_X1 U512 ( .A1(n700), .A2(G953), .ZN(n759) );
  NAND2_X1 U513 ( .A1(n603), .A2(n364), .ZN(n489) );
  NAND2_X1 U514 ( .A1(n751), .A2(G478), .ZN(n754) );
  XNOR2_X2 U515 ( .A(n415), .B(n414), .ZN(n460) );
  XNOR2_X2 U516 ( .A(n413), .B(G107), .ZN(n511) );
  XNOR2_X2 U517 ( .A(G122), .B(G116), .ZN(n413) );
  XNOR2_X2 U518 ( .A(KEYINPUT3), .B(G119), .ZN(n414) );
  XNOR2_X2 U519 ( .A(G113), .B(G101), .ZN(n415) );
  NAND2_X1 U520 ( .A1(n366), .A2(n422), .ZN(n582) );
  INV_X1 U521 ( .A(n421), .ZN(n417) );
  NAND2_X1 U522 ( .A1(n649), .A2(n477), .ZN(n422) );
  BUF_X1 U523 ( .A(n560), .Z(n669) );
  NAND2_X1 U524 ( .A1(n556), .A2(n555), .ZN(n557) );
  INV_X1 U525 ( .A(KEYINPUT72), .ZN(n445) );
  XNOR2_X1 U526 ( .A(n446), .B(n445), .ZN(n448) );
  INV_X1 U527 ( .A(KEYINPUT10), .ZN(n428) );
  INV_X1 U528 ( .A(KEYINPUT71), .ZN(n443) );
  XNOR2_X1 U529 ( .A(n448), .B(n447), .ZN(n451) );
  NOR2_X1 U530 ( .A1(n618), .A2(n617), .ZN(n620) );
  BUF_X1 U531 ( .A(n717), .Z(n735) );
  XNOR2_X1 U532 ( .A(n433), .B(n432), .ZN(n434) );
  BUF_X1 U533 ( .A(n649), .Z(n651) );
  XNOR2_X1 U534 ( .A(n752), .B(KEYINPUT120), .ZN(n753) );
  XNOR2_X1 U535 ( .A(n746), .B(n745), .ZN(n747) );
  AND2_X1 U536 ( .A1(n628), .A2(n687), .ZN(n599) );
  XNOR2_X2 U537 ( .A(G143), .B(G128), .ZN(n467) );
  XNOR2_X1 U538 ( .A(KEYINPUT70), .B(KEYINPUT69), .ZN(n426) );
  INV_X1 U539 ( .A(G469), .ZN(n425) );
  NAND2_X1 U540 ( .A1(G221), .A2(n508), .ZN(n429) );
  XOR2_X1 U541 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n430) );
  XNOR2_X1 U542 ( .A(n430), .B(n362), .ZN(n433) );
  XNOR2_X1 U543 ( .A(n363), .B(n431), .ZN(n432) );
  NAND2_X1 U544 ( .A1(n634), .A2(G234), .ZN(n436) );
  XNOR2_X1 U545 ( .A(n436), .B(KEYINPUT20), .ZN(n439) );
  XNOR2_X1 U546 ( .A(KEYINPUT25), .B(n361), .ZN(n437) );
  AND2_X1 U547 ( .A1(n439), .A2(G221), .ZN(n441) );
  INV_X1 U548 ( .A(KEYINPUT21), .ZN(n440) );
  XNOR2_X1 U549 ( .A(n441), .B(n440), .ZN(n705) );
  NOR2_X1 U550 ( .A1(n527), .A2(n705), .ZN(n442) );
  XNOR2_X1 U551 ( .A(n442), .B(KEYINPUT67), .ZN(n702) );
  NAND2_X1 U552 ( .A1(n492), .A2(G210), .ZN(n446) );
  XOR2_X1 U553 ( .A(KEYINPUT92), .B(KEYINPUT5), .Z(n447) );
  XNOR2_X1 U554 ( .A(n460), .B(n449), .ZN(n450) );
  XNOR2_X1 U555 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U556 ( .A(n358), .B(n452), .ZN(n671) );
  OR2_X1 U557 ( .A1(n671), .A2(G902), .ZN(n456) );
  INV_X1 U558 ( .A(KEYINPUT93), .ZN(n454) );
  XNOR2_X1 U559 ( .A(n454), .B(G472), .ZN(n455) );
  XNOR2_X2 U560 ( .A(n456), .B(n455), .ZN(n591) );
  INV_X1 U561 ( .A(KEYINPUT6), .ZN(n457) );
  NAND2_X1 U562 ( .A1(n536), .A2(n576), .ZN(n459) );
  INV_X1 U563 ( .A(KEYINPUT33), .ZN(n458) );
  XNOR2_X1 U564 ( .A(n461), .B(KEYINPUT16), .ZN(n462) );
  XNOR2_X1 U565 ( .A(n465), .B(n464), .ZN(n470) );
  NAND2_X1 U566 ( .A1(n776), .A2(G224), .ZN(n466) );
  XNOR2_X1 U567 ( .A(n466), .B(KEYINPUT74), .ZN(n468) );
  XNOR2_X1 U568 ( .A(n467), .B(n468), .ZN(n469) );
  XNOR2_X1 U569 ( .A(n470), .B(n469), .ZN(n471) );
  INV_X1 U570 ( .A(n634), .ZN(n472) );
  NAND2_X1 U571 ( .A1(n474), .A2(n473), .ZN(n478) );
  NAND2_X1 U572 ( .A1(n478), .A2(G210), .ZN(n476) );
  INV_X1 U573 ( .A(KEYINPUT87), .ZN(n475) );
  XNOR2_X1 U574 ( .A(n476), .B(n475), .ZN(n477) );
  NAND2_X1 U575 ( .A1(n478), .A2(G214), .ZN(n718) );
  XNOR2_X1 U576 ( .A(n479), .B(KEYINPUT14), .ZN(n481) );
  NAND2_X1 U577 ( .A1(n481), .A2(G952), .ZN(n480) );
  XNOR2_X1 U578 ( .A(n480), .B(KEYINPUT88), .ZN(n734) );
  NOR2_X1 U579 ( .A1(G953), .A2(n734), .ZN(n573) );
  NAND2_X1 U580 ( .A1(G902), .A2(n481), .ZN(n482) );
  XNOR2_X1 U581 ( .A(KEYINPUT89), .B(n482), .ZN(n483) );
  NAND2_X1 U582 ( .A1(n483), .A2(G953), .ZN(n570) );
  NOR2_X1 U583 ( .A1(G898), .A2(n570), .ZN(n484) );
  OR2_X1 U584 ( .A1(n573), .A2(n484), .ZN(n486) );
  INV_X1 U585 ( .A(KEYINPUT90), .ZN(n485) );
  INV_X1 U586 ( .A(KEYINPUT85), .ZN(n487) );
  XNOR2_X1 U587 ( .A(n487), .B(KEYINPUT0), .ZN(n488) );
  XNOR2_X1 U588 ( .A(n489), .B(n488), .ZN(n524) );
  BUF_X2 U589 ( .A(n524), .Z(n541) );
  XNOR2_X1 U590 ( .A(KEYINPUT98), .B(KEYINPUT13), .ZN(n504) );
  NAND2_X1 U591 ( .A1(G214), .A2(n492), .ZN(n493) );
  XNOR2_X1 U592 ( .A(n494), .B(n493), .ZN(n495) );
  XOR2_X1 U593 ( .A(n495), .B(KEYINPUT96), .Z(n501) );
  XNOR2_X1 U594 ( .A(n497), .B(n496), .ZN(n499) );
  XNOR2_X1 U595 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U596 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U597 ( .A(n502), .B(n767), .ZN(n661) );
  NOR2_X1 U598 ( .A1(G902), .A2(n661), .ZN(n503) );
  INV_X1 U599 ( .A(G475), .ZN(n505) );
  INV_X1 U600 ( .A(n543), .ZN(n517) );
  XOR2_X1 U601 ( .A(KEYINPUT100), .B(KEYINPUT9), .Z(n507) );
  XNOR2_X1 U602 ( .A(KEYINPUT7), .B(KEYINPUT99), .ZN(n506) );
  XNOR2_X1 U603 ( .A(n507), .B(n506), .ZN(n510) );
  NAND2_X1 U604 ( .A1(G217), .A2(n508), .ZN(n509) );
  XNOR2_X1 U605 ( .A(n510), .B(n509), .ZN(n514) );
  XNOR2_X1 U606 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U607 ( .A(n514), .B(n513), .ZN(n752) );
  OR2_X1 U608 ( .A1(n752), .A2(G902), .ZN(n516) );
  INV_X1 U609 ( .A(G478), .ZN(n515) );
  XNOR2_X1 U610 ( .A(n516), .B(n515), .ZN(n523) );
  INV_X1 U611 ( .A(n523), .ZN(n542) );
  NAND2_X1 U612 ( .A1(n517), .A2(n542), .ZN(n608) );
  INV_X1 U613 ( .A(n608), .ZN(n518) );
  INV_X1 U614 ( .A(n560), .ZN(n519) );
  NAND2_X1 U615 ( .A1(n519), .A2(KEYINPUT82), .ZN(n522) );
  NOR2_X1 U616 ( .A1(n384), .A2(KEYINPUT82), .ZN(n520) );
  NAND2_X1 U617 ( .A1(n560), .A2(n520), .ZN(n521) );
  NAND2_X1 U618 ( .A1(n522), .A2(n521), .ZN(n530) );
  NAND2_X1 U619 ( .A1(n543), .A2(n523), .ZN(n722) );
  OR2_X2 U620 ( .A1(n524), .A2(n424), .ZN(n526) );
  INV_X1 U621 ( .A(KEYINPUT22), .ZN(n525) );
  XNOR2_X2 U622 ( .A(n526), .B(n525), .ZN(n532) );
  AND2_X2 U623 ( .A1(n532), .A2(n706), .ZN(n549) );
  INV_X1 U624 ( .A(n703), .ZN(n622) );
  NOR2_X1 U625 ( .A1(n622), .A2(n591), .ZN(n528) );
  XOR2_X2 U626 ( .A(KEYINPUT103), .B(n529), .Z(n668) );
  INV_X1 U627 ( .A(n576), .ZN(n531) );
  XNOR2_X1 U628 ( .A(n533), .B(KEYINPUT80), .ZN(n535) );
  NOR2_X1 U629 ( .A1(n622), .A2(n706), .ZN(n534) );
  NAND2_X1 U630 ( .A1(n535), .A2(n534), .ZN(n658) );
  NAND2_X1 U631 ( .A1(n536), .A2(n591), .ZN(n713) );
  NOR2_X1 U632 ( .A1(n713), .A2(n541), .ZN(n538) );
  XNOR2_X1 U633 ( .A(KEYINPUT31), .B(KEYINPUT94), .ZN(n537) );
  XNOR2_X1 U634 ( .A(n538), .B(n537), .ZN(n694) );
  BUF_X1 U635 ( .A(n539), .Z(n587) );
  NOR2_X1 U636 ( .A1(n702), .A2(n587), .ZN(n594) );
  INV_X1 U637 ( .A(n591), .ZN(n708) );
  NAND2_X1 U638 ( .A1(n594), .A2(n708), .ZN(n540) );
  OR2_X1 U639 ( .A1(n541), .A2(n540), .ZN(n679) );
  NAND2_X1 U640 ( .A1(n694), .A2(n679), .ZN(n546) );
  NAND2_X1 U641 ( .A1(n543), .A2(n542), .ZN(n693) );
  XNOR2_X1 U642 ( .A(KEYINPUT101), .B(n693), .ZN(n629) );
  NOR2_X1 U643 ( .A1(n543), .A2(n542), .ZN(n687) );
  NOR2_X1 U644 ( .A1(n629), .A2(n687), .ZN(n544) );
  XNOR2_X1 U645 ( .A(n544), .B(KEYINPUT102), .ZN(n724) );
  XNOR2_X1 U646 ( .A(n724), .B(KEYINPUT77), .ZN(n545) );
  NAND2_X1 U647 ( .A1(n546), .A2(n545), .ZN(n547) );
  NAND2_X1 U648 ( .A1(n658), .A2(n547), .ZN(n553) );
  NOR2_X1 U649 ( .A1(n377), .A2(n576), .ZN(n548) );
  NAND2_X1 U650 ( .A1(n549), .A2(n548), .ZN(n551) );
  INV_X1 U651 ( .A(KEYINPUT32), .ZN(n550) );
  INV_X1 U652 ( .A(n553), .ZN(n556) );
  INV_X1 U653 ( .A(KEYINPUT82), .ZN(n554) );
  NOR2_X1 U654 ( .A1(n554), .A2(KEYINPUT44), .ZN(n555) );
  NAND2_X1 U655 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U656 ( .A(n559), .B(KEYINPUT81), .ZN(n565) );
  INV_X1 U657 ( .A(n660), .ZN(n561) );
  NAND2_X1 U658 ( .A1(n668), .A2(n561), .ZN(n562) );
  NOR2_X1 U659 ( .A1(n563), .A2(n562), .ZN(n564) );
  NOR2_X1 U660 ( .A1(n565), .A2(n564), .ZN(n568) );
  XOR2_X1 U661 ( .A(KEYINPUT79), .B(KEYINPUT45), .Z(n566) );
  XNOR2_X1 U662 ( .A(n568), .B(n567), .ZN(n637) );
  NOR2_X1 U663 ( .A1(n637), .A2(n634), .ZN(n569) );
  XNOR2_X1 U664 ( .A(n569), .B(KEYINPUT78), .ZN(n633) );
  INV_X1 U665 ( .A(n687), .ZN(n690) );
  XNOR2_X1 U666 ( .A(KEYINPUT104), .B(n570), .ZN(n571) );
  NOR2_X1 U667 ( .A1(G900), .A2(n571), .ZN(n572) );
  NOR2_X1 U668 ( .A1(n573), .A2(n572), .ZN(n596) );
  NOR2_X1 U669 ( .A1(n705), .A2(n596), .ZN(n574) );
  NAND2_X1 U670 ( .A1(n706), .A2(n574), .ZN(n585) );
  NOR2_X1 U671 ( .A1(n690), .A2(n585), .ZN(n575) );
  INV_X1 U672 ( .A(n577), .ZN(n578) );
  NOR2_X1 U673 ( .A1(n579), .A2(n578), .ZN(n580) );
  NAND2_X1 U674 ( .A1(n581), .A2(n622), .ZN(n697) );
  XNOR2_X1 U675 ( .A(n582), .B(KEYINPUT38), .ZN(n719) );
  NAND2_X1 U676 ( .A1(n719), .A2(n718), .ZN(n725) );
  NOR2_X1 U677 ( .A1(n722), .A2(n725), .ZN(n584) );
  XNOR2_X1 U678 ( .A(KEYINPUT41), .B(KEYINPUT106), .ZN(n583) );
  XNOR2_X1 U679 ( .A(n584), .B(n583), .ZN(n736) );
  NOR2_X1 U680 ( .A1(n708), .A2(n585), .ZN(n586) );
  XNOR2_X1 U681 ( .A(n586), .B(KEYINPUT28), .ZN(n589) );
  INV_X1 U682 ( .A(n587), .ZN(n588) );
  NAND2_X1 U683 ( .A1(n589), .A2(n588), .ZN(n602) );
  NOR2_X1 U684 ( .A1(n736), .A2(n602), .ZN(n590) );
  XNOR2_X1 U685 ( .A(KEYINPUT42), .B(n590), .ZN(n781) );
  NAND2_X1 U686 ( .A1(n591), .A2(n718), .ZN(n592) );
  XOR2_X1 U687 ( .A(KEYINPUT30), .B(n592), .Z(n593) );
  NAND2_X1 U688 ( .A1(n594), .A2(n593), .ZN(n595) );
  NOR2_X1 U689 ( .A1(n596), .A2(n595), .ZN(n610) );
  AND2_X1 U690 ( .A1(n610), .A2(n719), .ZN(n598) );
  XNOR2_X1 U691 ( .A(n599), .B(KEYINPUT40), .ZN(n780) );
  NOR2_X1 U692 ( .A1(n781), .A2(n780), .ZN(n600) );
  XNOR2_X1 U693 ( .A(n600), .B(KEYINPUT46), .ZN(n601) );
  NAND2_X1 U694 ( .A1(n697), .A2(n601), .ZN(n618) );
  INV_X1 U695 ( .A(n602), .ZN(n604) );
  NAND2_X1 U696 ( .A1(n604), .A2(n603), .ZN(n686) );
  INV_X1 U697 ( .A(KEYINPUT77), .ZN(n606) );
  INV_X1 U698 ( .A(n724), .ZN(n605) );
  OR2_X1 U699 ( .A1(n606), .A2(n605), .ZN(n607) );
  NOR2_X1 U700 ( .A1(n686), .A2(n607), .ZN(n611) );
  NOR2_X1 U701 ( .A1(n608), .A2(n582), .ZN(n609) );
  AND2_X1 U702 ( .A1(n610), .A2(n609), .ZN(n657) );
  NOR2_X1 U703 ( .A1(n611), .A2(n657), .ZN(n616) );
  NOR2_X1 U704 ( .A1(n724), .A2(n686), .ZN(n612) );
  XOR2_X1 U705 ( .A(n612), .B(KEYINPUT47), .Z(n614) );
  NAND2_X1 U706 ( .A1(n612), .A2(KEYINPUT77), .ZN(n613) );
  NAND2_X1 U707 ( .A1(n614), .A2(n613), .ZN(n615) );
  NAND2_X1 U708 ( .A1(n616), .A2(n615), .ZN(n617) );
  NOR2_X1 U709 ( .A1(n622), .A2(n621), .ZN(n623) );
  NAND2_X1 U710 ( .A1(n718), .A2(n623), .ZN(n624) );
  XOR2_X1 U711 ( .A(KEYINPUT105), .B(n624), .Z(n625) );
  XOR2_X1 U712 ( .A(KEYINPUT43), .B(n625), .Z(n627) );
  INV_X1 U713 ( .A(n582), .ZN(n626) );
  OR2_X1 U714 ( .A1(n627), .A2(n626), .ZN(n659) );
  NAND2_X1 U715 ( .A1(n629), .A2(n628), .ZN(n698) );
  NAND2_X1 U716 ( .A1(n659), .A2(n698), .ZN(n630) );
  NOR2_X1 U717 ( .A1(n641), .A2(n630), .ZN(n768) );
  XNOR2_X1 U718 ( .A(n768), .B(n631), .ZN(n632) );
  BUF_X1 U719 ( .A(n637), .Z(n700) );
  NAND2_X1 U720 ( .A1(KEYINPUT2), .A2(n698), .ZN(n638) );
  XOR2_X1 U721 ( .A(KEYINPUT76), .B(n638), .Z(n639) );
  NAND2_X1 U722 ( .A1(n639), .A2(n659), .ZN(n640) );
  XNOR2_X1 U723 ( .A(n644), .B(n643), .ZN(n646) );
  NOR2_X1 U724 ( .A1(n776), .A2(G952), .ZN(n645) );
  NAND2_X1 U725 ( .A1(n646), .A2(n749), .ZN(n648) );
  INV_X1 U726 ( .A(KEYINPUT122), .ZN(n647) );
  XNOR2_X1 U727 ( .A(n648), .B(n647), .ZN(G66) );
  XNOR2_X1 U728 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n650) );
  XNOR2_X1 U729 ( .A(n653), .B(n652), .ZN(n654) );
  NAND2_X1 U730 ( .A1(n654), .A2(n749), .ZN(n656) );
  INV_X1 U731 ( .A(KEYINPUT56), .ZN(n655) );
  XNOR2_X1 U732 ( .A(n656), .B(n655), .ZN(G51) );
  XOR2_X1 U733 ( .A(G143), .B(n657), .Z(G45) );
  XNOR2_X1 U734 ( .A(n658), .B(G101), .ZN(G3) );
  XNOR2_X1 U735 ( .A(n659), .B(G140), .ZN(G42) );
  XOR2_X1 U736 ( .A(G119), .B(n660), .Z(G21) );
  XNOR2_X1 U737 ( .A(n663), .B(n662), .ZN(n664) );
  NAND2_X1 U738 ( .A1(n664), .A2(n749), .ZN(n667) );
  XOR2_X1 U739 ( .A(KEYINPUT119), .B(KEYINPUT60), .Z(n665) );
  XNOR2_X1 U740 ( .A(n665), .B(KEYINPUT65), .ZN(n666) );
  XNOR2_X1 U741 ( .A(n667), .B(n666), .ZN(G60) );
  XNOR2_X1 U742 ( .A(n668), .B(G110), .ZN(G12) );
  XOR2_X1 U743 ( .A(G122), .B(n669), .Z(G24) );
  XNOR2_X1 U744 ( .A(KEYINPUT109), .B(KEYINPUT62), .ZN(n670) );
  XNOR2_X1 U745 ( .A(n673), .B(n672), .ZN(n674) );
  NAND2_X1 U746 ( .A1(n674), .A2(n749), .ZN(n676) );
  XNOR2_X1 U747 ( .A(KEYINPUT84), .B(KEYINPUT63), .ZN(n675) );
  XNOR2_X1 U748 ( .A(n676), .B(n675), .ZN(G57) );
  NOR2_X1 U749 ( .A1(n679), .A2(n690), .ZN(n677) );
  XOR2_X1 U750 ( .A(KEYINPUT110), .B(n677), .Z(n678) );
  XNOR2_X1 U751 ( .A(G104), .B(n678), .ZN(G6) );
  NOR2_X1 U752 ( .A1(n693), .A2(n679), .ZN(n683) );
  XOR2_X1 U753 ( .A(KEYINPUT26), .B(KEYINPUT111), .Z(n681) );
  XNOR2_X1 U754 ( .A(G107), .B(KEYINPUT27), .ZN(n680) );
  XNOR2_X1 U755 ( .A(n681), .B(n680), .ZN(n682) );
  XNOR2_X1 U756 ( .A(n683), .B(n682), .ZN(G9) );
  NOR2_X1 U757 ( .A1(n686), .A2(n693), .ZN(n685) );
  XNOR2_X1 U758 ( .A(G128), .B(KEYINPUT29), .ZN(n684) );
  XNOR2_X1 U759 ( .A(n685), .B(n684), .ZN(G30) );
  INV_X1 U760 ( .A(n686), .ZN(n688) );
  NAND2_X1 U761 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U762 ( .A(n689), .B(G146), .ZN(G48) );
  NOR2_X1 U763 ( .A1(n694), .A2(n690), .ZN(n691) );
  XOR2_X1 U764 ( .A(KEYINPUT112), .B(n691), .Z(n692) );
  XNOR2_X1 U765 ( .A(G113), .B(n692), .ZN(G15) );
  NOR2_X1 U766 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U767 ( .A(G116), .B(n695), .Z(G18) );
  XOR2_X1 U768 ( .A(G125), .B(KEYINPUT37), .Z(n696) );
  XNOR2_X1 U769 ( .A(n697), .B(n696), .ZN(G27) );
  XNOR2_X1 U770 ( .A(G134), .B(n698), .ZN(G36) );
  XOR2_X1 U771 ( .A(KEYINPUT53), .B(KEYINPUT118), .Z(n744) );
  NAND2_X1 U772 ( .A1(n359), .A2(n768), .ZN(n699) );
  NOR2_X1 U773 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U774 ( .A1(n701), .A2(G953), .ZN(n742) );
  XOR2_X1 U775 ( .A(KEYINPUT52), .B(KEYINPUT116), .Z(n732) );
  NAND2_X1 U776 ( .A1(n377), .A2(n702), .ZN(n704) );
  XNOR2_X1 U777 ( .A(n704), .B(KEYINPUT50), .ZN(n712) );
  NAND2_X1 U778 ( .A1(n706), .A2(n705), .ZN(n707) );
  XOR2_X1 U779 ( .A(KEYINPUT49), .B(n707), .Z(n709) );
  NAND2_X1 U780 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U781 ( .A(KEYINPUT113), .B(n710), .ZN(n711) );
  NAND2_X1 U782 ( .A1(n712), .A2(n711), .ZN(n714) );
  NAND2_X1 U783 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U784 ( .A(KEYINPUT51), .B(n715), .ZN(n716) );
  NOR2_X1 U785 ( .A1(n736), .A2(n716), .ZN(n730) );
  NOR2_X1 U786 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U787 ( .A(n720), .B(KEYINPUT114), .ZN(n721) );
  NOR2_X1 U788 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U789 ( .A(KEYINPUT115), .B(n723), .Z(n727) );
  NOR2_X1 U790 ( .A1(n725), .A2(n724), .ZN(n726) );
  NOR2_X1 U791 ( .A1(n727), .A2(n726), .ZN(n728) );
  NOR2_X1 U792 ( .A1(n735), .A2(n728), .ZN(n729) );
  NOR2_X1 U793 ( .A1(n730), .A2(n729), .ZN(n731) );
  XOR2_X1 U794 ( .A(n732), .B(n731), .Z(n733) );
  NOR2_X1 U795 ( .A1(n734), .A2(n733), .ZN(n738) );
  NOR2_X1 U796 ( .A1(n736), .A2(n735), .ZN(n737) );
  NOR2_X1 U797 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U798 ( .A(n739), .B(KEYINPUT117), .ZN(n740) );
  NOR2_X1 U799 ( .A1(n740), .A2(n367), .ZN(n741) );
  NAND2_X1 U800 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U801 ( .A(n744), .B(n743), .ZN(G75) );
  NAND2_X1 U802 ( .A1(n751), .A2(G469), .ZN(n748) );
  XOR2_X1 U803 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n745) );
  INV_X1 U804 ( .A(n749), .ZN(n755) );
  NOR2_X1 U805 ( .A1(n750), .A2(n755), .ZN(G54) );
  NAND2_X1 U806 ( .A1(G953), .A2(G224), .ZN(n756) );
  XNOR2_X1 U807 ( .A(KEYINPUT61), .B(n756), .ZN(n757) );
  NAND2_X1 U808 ( .A1(n757), .A2(G898), .ZN(n758) );
  NAND2_X1 U809 ( .A1(n759), .A2(n758), .ZN(n764) );
  OR2_X1 U810 ( .A1(G898), .A2(n776), .ZN(n760) );
  NAND2_X1 U811 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U812 ( .A(n762), .B(KEYINPUT123), .ZN(n763) );
  XNOR2_X1 U813 ( .A(n764), .B(n763), .ZN(G69) );
  BUF_X1 U814 ( .A(n765), .Z(n766) );
  XNOR2_X1 U815 ( .A(n767), .B(n766), .ZN(n771) );
  XOR2_X1 U816 ( .A(n768), .B(n771), .Z(n769) );
  NOR2_X1 U817 ( .A1(G953), .A2(n769), .ZN(n770) );
  XOR2_X1 U818 ( .A(KEYINPUT124), .B(n770), .Z(n779) );
  XNOR2_X1 U819 ( .A(n771), .B(G227), .ZN(n772) );
  XNOR2_X1 U820 ( .A(n772), .B(KEYINPUT125), .ZN(n773) );
  NAND2_X1 U821 ( .A1(n773), .A2(G900), .ZN(n774) );
  XOR2_X1 U822 ( .A(KEYINPUT126), .B(n774), .Z(n775) );
  NOR2_X1 U823 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U824 ( .A(KEYINPUT127), .B(n777), .ZN(n778) );
  NAND2_X1 U825 ( .A1(n779), .A2(n778), .ZN(G72) );
  XOR2_X1 U826 ( .A(G131), .B(n780), .Z(G33) );
  XOR2_X1 U827 ( .A(G137), .B(n781), .Z(G39) );
endmodule

