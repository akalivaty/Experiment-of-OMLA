//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 0 0 0 0 1 1 0 0 0 1 1 1 1 0 0 1 0 0 1 1 1 1 0 1 1 1 1 0 0 1 0 0 0 0 0 0 0 0 0 1 1 1 1 1 1 1 0 1 1 1 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:13 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n551,
    new_n552, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n612, new_n613, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n841, new_n842, new_n843,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT64), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT65), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n453), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G125), .ZN(new_n462));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n461), .A2(G137), .A3(new_n460), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n460), .A2(G101), .A3(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n464), .A2(new_n467), .ZN(G160));
  NAND2_X1  g043(.A1(new_n461), .A2(new_n460), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G136), .ZN(new_n471));
  XOR2_X1   g046(.A(new_n471), .B(KEYINPUT66), .Z(new_n472));
  OAI21_X1  g047(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n473));
  INV_X1    g048(.A(G112), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n473), .B1(new_n474), .B2(G2105), .ZN(new_n475));
  XNOR2_X1  g050(.A(new_n475), .B(KEYINPUT67), .ZN(new_n476));
  OR2_X1    g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n460), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n476), .B1(G124), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n472), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT68), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n481), .B(new_n482), .ZN(G162));
  OAI21_X1  g058(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n485), .B1(G114), .B2(new_n460), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n461), .A2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G126), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  AND2_X1   g064(.A1(new_n460), .A2(G138), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n461), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n461), .A2(new_n493), .A3(new_n490), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n489), .B1(new_n492), .B2(new_n494), .ZN(G164));
  INV_X1    g070(.A(G543), .ZN(new_n496));
  OR2_X1    g071(.A1(KEYINPUT6), .A2(G651), .ZN(new_n497));
  NAND2_X1  g072(.A1(KEYINPUT6), .A2(G651), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G50), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT69), .ZN(new_n501));
  XNOR2_X1  g076(.A(new_n500), .B(new_n501), .ZN(new_n502));
  XNOR2_X1  g077(.A(KEYINPUT5), .B(G543), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n503), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n497), .A2(new_n498), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(new_n503), .ZN(new_n507));
  INV_X1    g082(.A(G88), .ZN(new_n508));
  OAI22_X1  g083(.A1(new_n504), .A2(new_n505), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n502), .A2(new_n509), .ZN(G166));
  XNOR2_X1  g085(.A(KEYINPUT72), .B(KEYINPUT7), .ZN(new_n511));
  AND3_X1   g086(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OR2_X1    g088(.A1(new_n511), .A2(new_n512), .ZN(new_n514));
  AND2_X1   g089(.A1(new_n506), .A2(new_n503), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n513), .A2(new_n514), .B1(new_n515), .B2(G89), .ZN(new_n516));
  AND2_X1   g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NOR2_X1   g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  OAI21_X1  g093(.A(KEYINPUT70), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT5), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(new_n496), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT70), .ZN(new_n522));
  NAND2_X1  g097(.A1(KEYINPUT5), .A2(G543), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  AND2_X1   g099(.A1(G63), .A2(G651), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n519), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n499), .A2(G51), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT71), .ZN(new_n528));
  AND3_X1   g103(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n528), .B1(new_n526), .B2(new_n527), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n516), .B1(new_n529), .B2(new_n530), .ZN(G286));
  INV_X1    g106(.A(G286), .ZN(G168));
  NAND3_X1  g107(.A1(new_n519), .A2(new_n524), .A3(G64), .ZN(new_n533));
  NAND2_X1  g108(.A1(G77), .A2(G543), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n505), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n499), .A2(G52), .ZN(new_n536));
  INV_X1    g111(.A(G90), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n536), .B1(new_n537), .B2(new_n507), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n535), .A2(new_n538), .ZN(G171));
  XNOR2_X1  g114(.A(KEYINPUT74), .B(G81), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n515), .A2(new_n540), .B1(G43), .B2(new_n499), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n519), .A2(new_n524), .A3(G56), .ZN(new_n542));
  NAND2_X1  g117(.A1(G68), .A2(G543), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n505), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT73), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n541), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AOI211_X1 g121(.A(KEYINPUT73), .B(new_n505), .C1(new_n542), .C2(new_n543), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(G188));
  NAND2_X1  g128(.A1(G78), .A2(G543), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n517), .A2(new_n518), .ZN(new_n555));
  INV_X1    g130(.A(G65), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  AOI22_X1  g132(.A1(G91), .A2(new_n515), .B1(new_n557), .B2(G651), .ZN(new_n558));
  INV_X1    g133(.A(new_n498), .ZN(new_n559));
  NOR2_X1   g134(.A1(KEYINPUT6), .A2(G651), .ZN(new_n560));
  OAI211_X1 g135(.A(G53), .B(G543), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT9), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n558), .A2(new_n562), .ZN(G299));
  INV_X1    g138(.A(G171), .ZN(G301));
  OR2_X1    g139(.A1(new_n502), .A2(new_n509), .ZN(G303));
  NAND2_X1  g140(.A1(new_n499), .A2(G49), .ZN(new_n566));
  XOR2_X1   g141(.A(new_n566), .B(KEYINPUT75), .Z(new_n567));
  AND2_X1   g142(.A1(new_n519), .A2(new_n524), .ZN(new_n568));
  OAI21_X1  g143(.A(G651), .B1(new_n568), .B2(G74), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n515), .A2(G87), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(G288));
  INV_X1    g148(.A(G73), .ZN(new_n574));
  OR3_X1    g149(.A1(new_n574), .A2(new_n496), .A3(KEYINPUT76), .ZN(new_n575));
  OAI21_X1  g150(.A(KEYINPUT76), .B1(new_n574), .B2(new_n496), .ZN(new_n576));
  INV_X1    g151(.A(G61), .ZN(new_n577));
  OAI211_X1 g152(.A(new_n575), .B(new_n576), .C1(new_n577), .C2(new_n555), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n578), .A2(G651), .B1(new_n515), .B2(G86), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT77), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n506), .A2(G543), .ZN(new_n581));
  INV_X1    g156(.A(G48), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n499), .A2(KEYINPUT77), .A3(G48), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n579), .A2(new_n585), .ZN(G305));
  NAND2_X1  g161(.A1(new_n568), .A2(G60), .ZN(new_n587));
  NAND2_X1  g162(.A1(G72), .A2(G543), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n505), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n499), .A2(G47), .ZN(new_n590));
  INV_X1    g165(.A(G85), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n591), .B2(new_n507), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(G290));
  INV_X1    g169(.A(KEYINPUT10), .ZN(new_n595));
  INV_X1    g170(.A(G92), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n507), .B2(new_n596), .ZN(new_n597));
  NAND4_X1  g172(.A1(new_n506), .A2(new_n503), .A3(KEYINPUT10), .A4(G92), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(G79), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G66), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n555), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n602), .A2(G651), .B1(G54), .B2(new_n499), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(new_n605), .B2(G171), .ZN(G284));
  OAI21_X1  g182(.A(new_n606), .B1(new_n605), .B2(G171), .ZN(G321));
  NAND2_X1  g183(.A1(G299), .A2(new_n605), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G168), .B2(new_n605), .ZN(G297));
  OAI21_X1  g185(.A(new_n609), .B1(G168), .B2(new_n605), .ZN(G280));
  INV_X1    g186(.A(new_n604), .ZN(new_n612));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(G860), .ZN(G148));
  NAND2_X1  g189(.A1(new_n612), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(G868), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(G868), .B2(new_n548), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g193(.A1(new_n479), .A2(G123), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n460), .A2(G111), .ZN(new_n620));
  OAI21_X1  g195(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n621));
  INV_X1    g196(.A(G135), .ZN(new_n622));
  OAI221_X1 g197(.A(new_n619), .B1(new_n620), .B2(new_n621), .C1(new_n622), .C2(new_n469), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(G2096), .Z(new_n624));
  NAND3_X1  g199(.A1(new_n460), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT12), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT13), .ZN(new_n627));
  INV_X1    g202(.A(G2100), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n627), .A2(new_n628), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n624), .A2(new_n629), .A3(new_n630), .ZN(G156));
  INV_X1    g206(.A(KEYINPUT14), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2427), .B(G2438), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2430), .ZN(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT15), .B(G2435), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n632), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n636), .B1(new_n635), .B2(new_n634), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2451), .B(G2454), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT16), .ZN(new_n639));
  XNOR2_X1  g214(.A(G1341), .B(G1348), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n637), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2443), .B(G2446), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  AND3_X1   g220(.A1(new_n644), .A2(G14), .A3(new_n645), .ZN(G401));
  XOR2_X1   g221(.A(KEYINPUT78), .B(KEYINPUT18), .Z(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2084), .B(G2090), .Z(new_n649));
  XNOR2_X1  g224(.A(G2067), .B(G2678), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(KEYINPUT17), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n649), .A2(new_n650), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n648), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2072), .B(G2078), .Z(new_n655));
  AOI21_X1  g230(.A(new_n655), .B1(new_n651), .B2(new_n647), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n654), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2096), .B(G2100), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(G227));
  XNOR2_X1  g234(.A(G1981), .B(G1986), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1961), .B(G1966), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT79), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1956), .B(G2474), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1971), .B(G1976), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT19), .ZN(new_n667));
  OR3_X1    g242(.A1(new_n665), .A2(KEYINPUT81), .A3(new_n667), .ZN(new_n668));
  OAI21_X1  g243(.A(KEYINPUT81), .B1(new_n665), .B2(new_n667), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n663), .A2(new_n664), .ZN(new_n670));
  INV_X1    g245(.A(new_n667), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n671), .B1(new_n663), .B2(new_n664), .ZN(new_n672));
  AOI22_X1  g247(.A1(new_n668), .A2(new_n669), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  OAI21_X1  g248(.A(KEYINPUT80), .B1(new_n670), .B2(new_n667), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n663), .A2(new_n664), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT80), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n675), .A2(new_n676), .A3(new_n671), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n678), .A2(KEYINPUT20), .ZN(new_n679));
  INV_X1    g254(.A(KEYINPUT20), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(new_n674), .B2(new_n677), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n673), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1991), .B(G1996), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT82), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  OAI211_X1 g263(.A(new_n673), .B(new_n683), .C1(new_n679), .C2(new_n681), .ZN(new_n689));
  AND3_X1   g264(.A1(new_n685), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n688), .B1(new_n685), .B2(new_n689), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n661), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n685), .A2(new_n689), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(new_n687), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n685), .A2(new_n688), .A3(new_n689), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n694), .A2(new_n660), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n692), .A2(new_n696), .ZN(G229));
  NOR2_X1   g272(.A1(G29), .A2(G35), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(G162), .B2(G29), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT29), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(G2090), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n479), .A2(G128), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n460), .A2(G116), .ZN(new_n703));
  OAI21_X1  g278(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n704));
  INV_X1    g279(.A(G140), .ZN(new_n705));
  OAI221_X1 g280(.A(new_n702), .B1(new_n703), .B2(new_n704), .C1(new_n705), .C2(new_n469), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G29), .ZN(new_n707));
  INV_X1    g282(.A(G29), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G26), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT88), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT28), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n707), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(G2067), .ZN(new_n713));
  INV_X1    g288(.A(G16), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G20), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT23), .ZN(new_n716));
  INV_X1    g291(.A(G299), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n716), .B1(new_n717), .B2(new_n714), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(G1956), .ZN(new_n719));
  NOR2_X1   g294(.A1(G16), .A2(G19), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(new_n548), .B2(G16), .ZN(new_n721));
  AOI211_X1 g296(.A(new_n713), .B(new_n719), .C1(G1341), .C2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n714), .A2(G4), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(new_n612), .B2(new_n714), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT87), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(G1348), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n722), .B(new_n726), .C1(G1341), .C2(new_n721), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n701), .A2(new_n727), .ZN(new_n728));
  AND2_X1   g303(.A1(new_n708), .A2(G33), .ZN(new_n729));
  AND2_X1   g304(.A1(new_n461), .A2(G127), .ZN(new_n730));
  AND2_X1   g305(.A1(G115), .A2(G2104), .ZN(new_n731));
  OAI21_X1  g306(.A(G2105), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT89), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n732), .A2(new_n733), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT25), .ZN(new_n736));
  NAND2_X1  g311(.A1(G103), .A2(G2104), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n736), .B1(new_n737), .B2(G2105), .ZN(new_n738));
  NAND4_X1  g313(.A1(new_n460), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n739));
  AOI22_X1  g314(.A1(new_n470), .A2(G139), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n734), .A2(new_n735), .A3(new_n740), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT90), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n729), .B1(new_n742), .B2(G29), .ZN(new_n743));
  INV_X1    g318(.A(G2072), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n743), .A2(new_n744), .ZN(new_n746));
  INV_X1    g321(.A(G34), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n747), .A2(KEYINPUT24), .ZN(new_n748));
  AOI21_X1  g323(.A(G29), .B1(new_n747), .B2(KEYINPUT24), .ZN(new_n749));
  AOI22_X1  g324(.A1(G160), .A2(G29), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(G2084), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT91), .Z(new_n752));
  NAND3_X1  g327(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT26), .Z(new_n754));
  INV_X1    g329(.A(G129), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n754), .B1(new_n487), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n460), .A2(G105), .A3(G2104), .ZN(new_n757));
  INV_X1    g332(.A(G141), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n757), .B1(new_n469), .B2(new_n758), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n761), .A2(new_n708), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n708), .B2(G32), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT27), .B(G1996), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n752), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n745), .A2(new_n746), .A3(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT92), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n766), .A2(new_n767), .ZN(new_n769));
  NAND2_X1  g344(.A1(G168), .A2(G16), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n770), .B(KEYINPUT93), .C1(G16), .C2(G21), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(KEYINPUT93), .B2(new_n770), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n772), .A2(G1966), .ZN(new_n773));
  OAI22_X1  g348(.A1(new_n763), .A2(new_n764), .B1(G2084), .B2(new_n750), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT31), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n775), .A2(G11), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(G11), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT30), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n778), .A2(G28), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n708), .B1(new_n778), .B2(G28), .ZN(new_n780));
  OAI211_X1 g355(.A(new_n776), .B(new_n777), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n623), .A2(new_n708), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT94), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n783), .B2(new_n782), .ZN(new_n785));
  NOR2_X1   g360(.A1(G27), .A2(G29), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G164), .B2(G29), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G2078), .ZN(new_n788));
  NOR3_X1   g363(.A1(new_n774), .A2(new_n785), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n772), .A2(G1966), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n714), .A2(G5), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G171), .B2(new_n714), .ZN(new_n792));
  INV_X1    g367(.A(G1961), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  AND4_X1   g369(.A1(new_n773), .A2(new_n789), .A3(new_n790), .A4(new_n794), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n768), .A2(new_n769), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n796), .A2(KEYINPUT95), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT95), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n768), .A2(new_n798), .A3(new_n769), .A4(new_n795), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n728), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n714), .A2(G24), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(new_n593), .B2(new_n714), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G1986), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n708), .A2(G25), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n470), .A2(G131), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n479), .A2(G119), .ZN(new_n806));
  OR2_X1    g381(.A1(G95), .A2(G2105), .ZN(new_n807));
  OAI211_X1 g382(.A(new_n807), .B(G2104), .C1(G107), .C2(new_n460), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n805), .A2(new_n806), .A3(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n804), .B1(new_n810), .B2(new_n708), .ZN(new_n811));
  XOR2_X1   g386(.A(KEYINPUT35), .B(G1991), .Z(new_n812));
  XOR2_X1   g387(.A(new_n811), .B(new_n812), .Z(new_n813));
  NOR2_X1   g388(.A1(new_n803), .A2(new_n813), .ZN(new_n814));
  MUX2_X1   g389(.A(G6), .B(G305), .S(G16), .Z(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT84), .ZN(new_n816));
  XNOR2_X1  g391(.A(KEYINPUT32), .B(G1981), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  AND2_X1   g393(.A1(new_n714), .A2(G23), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(G288), .B2(G16), .ZN(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT33), .B(G1976), .ZN(new_n821));
  AND2_X1   g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n714), .A2(G22), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(G166), .B2(new_n714), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(G1971), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n820), .A2(new_n821), .ZN(new_n826));
  NOR3_X1   g401(.A1(new_n822), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n818), .A2(new_n827), .ZN(new_n828));
  XOR2_X1   g403(.A(KEYINPUT83), .B(KEYINPUT34), .Z(new_n829));
  OAI21_X1  g404(.A(new_n814), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT85), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n828), .A2(new_n829), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT36), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n835), .A2(KEYINPUT86), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n836), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n832), .A2(new_n833), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n800), .B1(new_n837), .B2(new_n839), .ZN(G311));
  INV_X1    g415(.A(new_n800), .ZN(new_n841));
  AND3_X1   g416(.A1(new_n832), .A2(new_n833), .A3(new_n838), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n838), .B1(new_n832), .B2(new_n833), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n841), .B1(new_n842), .B2(new_n843), .ZN(G150));
  NAND2_X1  g419(.A1(new_n612), .A2(G559), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT38), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n519), .A2(new_n524), .A3(G67), .ZN(new_n847));
  NAND2_X1  g422(.A1(G80), .A2(G543), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n505), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n506), .A2(new_n503), .A3(G93), .ZN(new_n850));
  OAI211_X1 g425(.A(G55), .B(G543), .C1(new_n559), .C2(new_n560), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT96), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n850), .A2(KEYINPUT96), .A3(new_n851), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n849), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  AND2_X1   g431(.A1(new_n542), .A2(new_n543), .ZN(new_n857));
  OAI21_X1  g432(.A(KEYINPUT73), .B1(new_n857), .B2(new_n505), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n544), .A2(new_n545), .ZN(new_n859));
  NAND4_X1  g434(.A1(new_n856), .A2(new_n858), .A3(new_n859), .A4(new_n541), .ZN(new_n860));
  AND3_X1   g435(.A1(new_n850), .A2(KEYINPUT96), .A3(new_n851), .ZN(new_n861));
  AOI21_X1  g436(.A(KEYINPUT96), .B1(new_n850), .B2(new_n851), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OAI22_X1  g438(.A1(new_n546), .A2(new_n547), .B1(new_n863), .B2(new_n849), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n860), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n846), .B(new_n866), .ZN(new_n867));
  OR2_X1    g442(.A1(new_n867), .A2(KEYINPUT39), .ZN(new_n868));
  INV_X1    g443(.A(G860), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(KEYINPUT39), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n856), .A2(new_n869), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT37), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(new_n873), .ZN(G145));
  XNOR2_X1  g449(.A(new_n623), .B(G160), .ZN(new_n875));
  XNOR2_X1  g450(.A(G162), .B(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n479), .A2(G130), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n460), .A2(G118), .ZN(new_n878));
  OAI21_X1  g453(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n880), .B1(G142), .B2(new_n470), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(new_n626), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(new_n809), .ZN(new_n883));
  INV_X1    g458(.A(new_n742), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n492), .A2(new_n494), .ZN(new_n885));
  INV_X1    g460(.A(G114), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n484), .B1(new_n886), .B2(G2105), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n887), .B1(G126), .B2(new_n479), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(new_n706), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(new_n761), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n884), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n890), .B(new_n760), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(new_n741), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n883), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT97), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n892), .A2(new_n894), .A3(new_n883), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AOI211_X1 g473(.A(KEYINPUT97), .B(new_n883), .C1(new_n892), .C2(new_n894), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n876), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n876), .A2(new_n895), .ZN(new_n901));
  AOI21_X1  g476(.A(G37), .B1(new_n901), .B2(new_n897), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g479(.A(KEYINPUT99), .B1(new_n856), .B2(G868), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n572), .A2(new_n593), .ZN(new_n906));
  OAI22_X1  g481(.A1(new_n567), .A2(new_n571), .B1(new_n589), .B2(new_n592), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(KEYINPUT98), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT98), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n906), .A2(new_n910), .A3(new_n907), .ZN(new_n911));
  XNOR2_X1  g486(.A(G166), .B(G305), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n909), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n912), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n914), .A2(new_n910), .A3(new_n907), .A4(new_n906), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n916), .B(KEYINPUT42), .ZN(new_n917));
  XOR2_X1   g492(.A(new_n865), .B(new_n615), .Z(new_n918));
  NAND2_X1  g493(.A1(new_n604), .A2(G299), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n599), .A2(new_n558), .A3(new_n562), .A4(new_n603), .ZN(new_n920));
  AOI21_X1  g495(.A(KEYINPUT41), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n919), .A2(KEYINPUT41), .A3(new_n920), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n918), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n919), .A2(new_n920), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n923), .B1(new_n925), .B2(new_n918), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n605), .B1(new_n917), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n927), .B1(new_n926), .B2(new_n917), .ZN(new_n928));
  MUX2_X1   g503(.A(KEYINPUT99), .B(new_n905), .S(new_n928), .Z(G295));
  MUX2_X1   g504(.A(KEYINPUT99), .B(new_n905), .S(new_n928), .Z(G331));
  NOR2_X1   g505(.A1(new_n922), .A2(new_n921), .ZN(new_n931));
  OAI221_X1 g506(.A(new_n516), .B1(new_n535), .B2(new_n538), .C1(new_n529), .C2(new_n530), .ZN(new_n932));
  NAND2_X1  g507(.A1(G286), .A2(G171), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n865), .A2(new_n934), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n860), .A2(new_n864), .A3(new_n933), .A4(new_n932), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n931), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT102), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT102), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n931), .A2(new_n935), .A3(new_n939), .A4(new_n936), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n935), .A2(new_n936), .ZN(new_n941));
  AOI21_X1  g516(.A(KEYINPUT103), .B1(new_n941), .B2(new_n925), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT103), .ZN(new_n943));
  AOI211_X1 g518(.A(new_n943), .B(new_n924), .C1(new_n935), .C2(new_n936), .ZN(new_n944));
  OAI211_X1 g519(.A(new_n938), .B(new_n940), .C1(new_n942), .C2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n916), .ZN(new_n946));
  INV_X1    g521(.A(G37), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT104), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n949), .B1(new_n945), .B2(new_n916), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n938), .A2(new_n940), .ZN(new_n951));
  INV_X1    g526(.A(new_n936), .ZN(new_n952));
  AOI22_X1  g527(.A1(new_n860), .A2(new_n864), .B1(new_n932), .B2(new_n933), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n925), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(new_n943), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n941), .A2(KEYINPUT103), .A3(new_n925), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n916), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n951), .A2(new_n957), .A3(KEYINPUT104), .A4(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n948), .B1(new_n950), .B2(new_n959), .ZN(new_n960));
  XNOR2_X1  g535(.A(KEYINPUT101), .B(KEYINPUT43), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT105), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT43), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n950), .A2(new_n959), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n954), .A2(new_n937), .ZN(new_n966));
  AOI21_X1  g541(.A(G37), .B1(new_n916), .B2(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n964), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  OAI211_X1 g543(.A(new_n962), .B(KEYINPUT44), .C1(new_n963), .C2(new_n968), .ZN(new_n969));
  AND2_X1   g544(.A1(new_n968), .A2(new_n963), .ZN(new_n970));
  XOR2_X1   g545(.A(KEYINPUT100), .B(KEYINPUT44), .Z(new_n971));
  AOI21_X1  g546(.A(G37), .B1(new_n945), .B2(new_n916), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n961), .B1(new_n965), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n961), .ZN(new_n974));
  INV_X1    g549(.A(new_n967), .ZN(new_n975));
  AOI211_X1 g550(.A(new_n974), .B(new_n975), .C1(new_n950), .C2(new_n959), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  OAI22_X1  g552(.A1(new_n969), .A2(new_n970), .B1(new_n971), .B2(new_n977), .ZN(G397));
  INV_X1    g553(.A(G1384), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n889), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT45), .ZN(new_n981));
  INV_X1    g556(.A(G40), .ZN(new_n982));
  NOR3_X1   g557(.A1(new_n464), .A2(new_n467), .A3(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n980), .A2(new_n981), .A3(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(G1996), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n760), .B(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G2067), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n706), .B(new_n988), .ZN(new_n989));
  OR2_X1    g564(.A1(new_n810), .A2(new_n812), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n810), .A2(new_n812), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n987), .A2(new_n989), .A3(new_n990), .A4(new_n991), .ZN(new_n992));
  XOR2_X1   g567(.A(new_n593), .B(G1986), .Z(new_n993));
  OAI21_X1  g568(.A(new_n985), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(G1384), .B1(new_n885), .B2(new_n888), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n995), .A2(new_n983), .A3(new_n988), .ZN(new_n996));
  OR2_X1    g571(.A1(new_n996), .A2(KEYINPUT116), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(KEYINPUT116), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT50), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n983), .B1(new_n995), .B2(new_n999), .ZN(new_n1000));
  NOR3_X1   g575(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n997), .B(new_n998), .C1(new_n1002), .C2(G1348), .ZN(new_n1003));
  NOR3_X1   g578(.A1(new_n1003), .A2(KEYINPUT60), .A3(new_n604), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n1003), .B(new_n612), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1004), .B1(new_n1005), .B2(KEYINPUT60), .ZN(new_n1006));
  XNOR2_X1  g581(.A(KEYINPUT114), .B(G1956), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1008), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT57), .ZN(new_n1010));
  OR2_X1    g585(.A1(new_n1010), .A2(KEYINPUT115), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(KEYINPUT115), .ZN(new_n1012));
  NAND3_X1  g587(.A1(G299), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n558), .A2(new_n562), .A3(KEYINPUT115), .A4(new_n1010), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n981), .B1(G164), .B2(G1384), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n995), .A2(KEYINPUT45), .ZN(new_n1017));
  XNOR2_X1  g592(.A(KEYINPUT56), .B(G2072), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1016), .A2(new_n1017), .A3(new_n983), .A4(new_n1018), .ZN(new_n1019));
  AND3_X1   g594(.A1(new_n1009), .A2(new_n1015), .A3(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1015), .B1(new_n1009), .B2(new_n1019), .ZN(new_n1021));
  OAI211_X1 g596(.A(KEYINPUT119), .B(KEYINPUT61), .C1(new_n1020), .C2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1023));
  NAND2_X1  g598(.A1(G160), .A2(G40), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1024), .B1(new_n980), .B2(KEYINPUT50), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n995), .A2(new_n999), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1007), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  AND4_X1   g602(.A1(new_n1016), .A2(new_n983), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1028));
  OAI211_X1 g603(.A(KEYINPUT119), .B(new_n1023), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT61), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1009), .A2(new_n1015), .A3(new_n1019), .A4(KEYINPUT119), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1022), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(KEYINPUT117), .A2(KEYINPUT59), .ZN(new_n1034));
  XNOR2_X1  g609(.A(new_n1034), .B(KEYINPUT118), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1016), .A2(new_n1017), .A3(new_n986), .A4(new_n983), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n995), .A2(new_n983), .ZN(new_n1037));
  XOR2_X1   g612(.A(KEYINPUT58), .B(G1341), .Z(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1036), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(new_n548), .ZN(new_n1041));
  NOR2_X1   g616(.A1(KEYINPUT117), .A2(KEYINPUT59), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1035), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1035), .ZN(new_n1045));
  AOI211_X1 g620(.A(new_n1042), .B(new_n1045), .C1(new_n1040), .C2(new_n548), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  AND3_X1   g622(.A1(new_n1033), .A2(KEYINPUT120), .A3(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(KEYINPUT120), .B1(new_n1033), .B2(new_n1047), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1006), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  AND2_X1   g625(.A1(new_n1003), .A2(new_n612), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1020), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1021), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1050), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(G303), .A2(G8), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT55), .ZN(new_n1056));
  XNOR2_X1  g631(.A(new_n1055), .B(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1017), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n983), .B1(new_n995), .B2(KEYINPUT45), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  OAI22_X1  g636(.A1(G2090), .A2(new_n1058), .B1(new_n1061), .B2(G1971), .ZN(new_n1062));
  AND3_X1   g637(.A1(new_n1057), .A2(new_n1062), .A3(G8), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1057), .B1(new_n1062), .B2(G8), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n572), .A2(G1976), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT106), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1067), .B1(new_n1037), .B2(G8), .ZN(new_n1068));
  INV_X1    g643(.A(G8), .ZN(new_n1069));
  AOI211_X1 g644(.A(KEYINPUT106), .B(new_n1069), .C1(new_n995), .C2(new_n983), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1066), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(KEYINPUT107), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT107), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1066), .B(new_n1073), .C1(new_n1068), .C2(new_n1070), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1072), .A2(new_n1074), .A3(KEYINPUT52), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1037), .A2(G8), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(KEYINPUT106), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1037), .A2(new_n1067), .A3(G8), .ZN(new_n1078));
  AOI22_X1  g653(.A1(new_n1077), .A2(new_n1078), .B1(G1976), .B2(new_n572), .ZN(new_n1079));
  INV_X1    g654(.A(G1976), .ZN(new_n1080));
  AOI21_X1  g655(.A(KEYINPUT52), .B1(G288), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1082));
  INV_X1    g657(.A(G1981), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n579), .A2(new_n585), .A3(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1083), .B1(new_n579), .B2(new_n585), .ZN(new_n1086));
  OAI21_X1  g661(.A(KEYINPUT49), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1086), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT49), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1088), .A2(new_n1089), .A3(new_n1084), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1087), .A2(new_n1090), .ZN(new_n1091));
  AOI22_X1  g666(.A1(new_n1079), .A2(new_n1081), .B1(new_n1082), .B2(new_n1091), .ZN(new_n1092));
  AND3_X1   g667(.A1(new_n1075), .A2(new_n1092), .A3(KEYINPUT110), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT110), .B1(new_n1075), .B2(new_n1092), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1065), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT121), .ZN(new_n1097));
  XOR2_X1   g672(.A(KEYINPUT111), .B(G2084), .Z(new_n1098));
  AND3_X1   g673(.A1(new_n1025), .A2(new_n1026), .A3(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1024), .B1(new_n980), .B2(new_n981), .ZN(new_n1100));
  AOI21_X1  g675(.A(G1966), .B1(new_n1100), .B2(new_n1017), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1097), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1025), .A2(new_n1026), .A3(new_n1098), .ZN(new_n1103));
  INV_X1    g678(.A(G1966), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1104), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1103), .A2(new_n1105), .A3(KEYINPUT121), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1102), .A2(G168), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT122), .ZN(new_n1108));
  OAI21_X1  g683(.A(G8), .B1(new_n1108), .B2(KEYINPUT51), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1109), .B1(new_n1108), .B2(KEYINPUT51), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1107), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(G8), .ZN(new_n1113));
  AOI21_X1  g688(.A(KEYINPUT51), .B1(G286), .B2(G8), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1111), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(G286), .A2(G8), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1117), .B1(new_n1102), .B2(new_n1106), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(G2078), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1016), .A2(new_n1017), .A3(new_n1120), .A4(new_n983), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  AOI22_X1  g697(.A1(new_n1122), .A2(KEYINPUT53), .B1(new_n1058), .B2(new_n793), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT53), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1121), .A2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(G301), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT123), .ZN(new_n1127));
  OAI21_X1  g702(.A(KEYINPUT54), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1058), .A2(new_n793), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1100), .A2(KEYINPUT53), .A3(new_n1120), .A4(new_n1017), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1129), .A2(new_n1125), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(G171), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1129), .A2(new_n1125), .A3(G301), .A4(new_n1130), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  AOI22_X1  g709(.A1(new_n1116), .A2(new_n1119), .B1(new_n1128), .B2(new_n1134), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1132), .A2(new_n1127), .A3(KEYINPUT54), .A4(new_n1133), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1096), .A2(new_n1135), .A3(KEYINPUT124), .A4(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT124), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT54), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1127), .B1(new_n1131), .B2(G171), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1134), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  AOI22_X1  g716(.A1(new_n1107), .A2(new_n1110), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1141), .B(new_n1136), .C1(new_n1118), .C2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1138), .B1(new_n1143), .B2(new_n1095), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n1054), .A2(new_n1137), .A3(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1112), .A2(G8), .A3(G168), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT112), .ZN(new_n1147));
  XNOR2_X1  g722(.A(new_n1146), .B(new_n1147), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n1148), .B(new_n1065), .C1(new_n1093), .C2(new_n1094), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT63), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1075), .A2(new_n1092), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1152), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1065), .A2(new_n1148), .A3(new_n1153), .A4(KEYINPUT63), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT113), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NOR3_X1   g731(.A1(new_n1063), .A2(new_n1064), .A3(new_n1150), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1157), .A2(KEYINPUT113), .A3(new_n1153), .A4(new_n1148), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1151), .A2(new_n1156), .A3(new_n1158), .ZN(new_n1159));
  OAI211_X1 g734(.A(new_n1065), .B(new_n1126), .C1(new_n1093), .C2(new_n1094), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1118), .B1(new_n1111), .B2(new_n1115), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT62), .ZN(new_n1163));
  OAI21_X1  g738(.A(KEYINPUT125), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT125), .ZN(new_n1166));
  OAI211_X1 g741(.A(new_n1166), .B(KEYINPUT62), .C1(new_n1142), .C2(new_n1118), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1161), .A2(new_n1164), .A3(new_n1165), .A4(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1153), .A2(new_n1063), .ZN(new_n1169));
  XOR2_X1   g744(.A(new_n1082), .B(KEYINPUT108), .Z(new_n1170));
  AND2_X1   g745(.A1(new_n1082), .A2(new_n1091), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n572), .A2(new_n1080), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1084), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1170), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1169), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT109), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1169), .A2(KEYINPUT109), .A3(new_n1174), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1159), .A2(new_n1168), .A3(new_n1179), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n994), .B1(new_n1145), .B2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n984), .B1(new_n989), .B2(new_n761), .ZN(new_n1182));
  OR3_X1    g757(.A1(new_n984), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1183));
  OAI21_X1  g758(.A(KEYINPUT46), .B1(new_n984), .B2(G1996), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1182), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  XNOR2_X1  g760(.A(new_n1185), .B(KEYINPUT47), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n992), .A2(new_n985), .ZN(new_n1187));
  NOR3_X1   g762(.A1(G290), .A2(new_n984), .A3(G1986), .ZN(new_n1188));
  XNOR2_X1  g763(.A(new_n1188), .B(KEYINPUT126), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1187), .B1(new_n1189), .B2(KEYINPUT48), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1190), .B1(KEYINPUT48), .B2(new_n1189), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n987), .A2(new_n989), .ZN(new_n1192));
  OAI22_X1  g767(.A1(new_n1192), .A2(new_n991), .B1(G2067), .B2(new_n706), .ZN(new_n1193));
  AOI211_X1 g768(.A(new_n1186), .B(new_n1191), .C1(new_n985), .C2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1181), .A2(new_n1194), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g770(.A1(new_n965), .A2(new_n961), .A3(new_n967), .ZN(new_n1197));
  OAI21_X1  g771(.A(new_n1197), .B1(new_n960), .B2(new_n961), .ZN(new_n1198));
  INV_X1    g772(.A(G319), .ZN(new_n1199));
  NOR3_X1   g773(.A1(G401), .A2(new_n1199), .A3(G227), .ZN(new_n1200));
  NAND3_X1  g774(.A1(new_n692), .A2(new_n696), .A3(new_n1200), .ZN(new_n1201));
  AOI21_X1  g775(.A(new_n1201), .B1(new_n900), .B2(new_n902), .ZN(new_n1202));
  AOI21_X1  g776(.A(KEYINPUT127), .B1(new_n1198), .B2(new_n1202), .ZN(new_n1203));
  OAI211_X1 g777(.A(KEYINPUT127), .B(new_n1202), .C1(new_n973), .C2(new_n976), .ZN(new_n1204));
  INV_X1    g778(.A(new_n1204), .ZN(new_n1205));
  NOR2_X1   g779(.A1(new_n1203), .A2(new_n1205), .ZN(G308));
  NAND2_X1  g780(.A1(new_n1198), .A2(new_n1202), .ZN(G225));
endmodule


