//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 1 1 0 0 1 0 0 1 0 1 0 0 0 0 1 1 1 0 0 0 1 0 1 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 1 1 1 1 1 1 0 0 1 0 1 1 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:09 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1213,
    new_n1214, new_n1215, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1263,
    new_n1264, new_n1265;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  INV_X1    g0009(.A(G68), .ZN(new_n210));
  INV_X1    g0010(.A(G238), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(G87), .ZN(new_n213));
  INV_X1    g0013(.A(G250), .ZN(new_n214));
  INV_X1    g0014(.A(G97), .ZN(new_n215));
  INV_X1    g0015(.A(G257), .ZN(new_n216));
  OAI22_X1  g0016(.A1(new_n213), .A2(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  AOI211_X1 g0017(.A(new_n212), .B(new_n217), .C1(G107), .C2(G264), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G116), .A2(G270), .ZN(new_n219));
  AND2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G50), .ZN(new_n221));
  INV_X1    g0021(.A(G226), .ZN(new_n222));
  INV_X1    g0022(.A(G77), .ZN(new_n223));
  INV_X1    g0023(.A(G244), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(G58), .ZN(new_n226));
  INV_X1    g0026(.A(G232), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n206), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT1), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n204), .A2(KEYINPUT64), .ZN(new_n231));
  INV_X1    g0031(.A(KEYINPUT64), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(G20), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g0034(.A1(G1), .A2(G13), .ZN(new_n235));
  NOR2_X1   g0035(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT65), .ZN(new_n237));
  OAI21_X1  g0037(.A(G50), .B1(G58), .B2(G68), .ZN(new_n238));
  INV_X1    g0038(.A(new_n238), .ZN(new_n239));
  AOI211_X1 g0039(.A(new_n209), .B(new_n230), .C1(new_n237), .C2(new_n239), .ZN(G361));
  XOR2_X1   g0040(.A(G238), .B(G244), .Z(new_n241));
  XNOR2_X1  g0041(.A(G226), .B(G232), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  XNOR2_X1  g0045(.A(G250), .B(G257), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(G264), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n247), .B(G270), .Z(new_n248));
  XOR2_X1   g0048(.A(new_n245), .B(new_n248), .Z(G358));
  XNOR2_X1  g0049(.A(G87), .B(G97), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(KEYINPUT67), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G107), .B(G116), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g0053(.A(G68), .B(G77), .Z(new_n254));
  XNOR2_X1  g0054(.A(G50), .B(G58), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n253), .B(new_n256), .ZN(G351));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  INV_X1    g0058(.A(G41), .ZN(new_n259));
  OAI211_X1 g0059(.A(G1), .B(G13), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT3), .B(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G1698), .ZN(new_n263));
  XNOR2_X1  g0063(.A(new_n263), .B(KEYINPUT70), .ZN(new_n264));
  XOR2_X1   g0064(.A(KEYINPUT71), .B(G223), .Z(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n258), .A2(KEYINPUT3), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT3), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n270), .A2(G1698), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G222), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n272), .B1(new_n223), .B2(new_n262), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n261), .B1(new_n266), .B2(new_n273), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n260), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  OR2_X1    g0077(.A1(KEYINPUT69), .A2(G226), .ZN(new_n278));
  NAND2_X1  g0078(.A1(KEYINPUT69), .A2(G226), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n203), .B(G274), .C1(G41), .C2(G45), .ZN(new_n281));
  XNOR2_X1  g0081(.A(new_n281), .B(KEYINPUT68), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n274), .A2(new_n280), .A3(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G190), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(new_n235), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n203), .A2(G20), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n288), .A2(G50), .A3(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n291));
  NOR2_X1   g0091(.A1(G58), .A2(G68), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n221), .ZN(new_n293));
  NOR2_X1   g0093(.A1(G20), .A2(G33), .ZN(new_n294));
  AOI22_X1  g0094(.A1(new_n293), .A2(G20), .B1(G150), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n234), .A2(G33), .ZN(new_n296));
  XNOR2_X1  g0096(.A(KEYINPUT8), .B(G58), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n295), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(new_n287), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT72), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(KEYINPUT72), .B1(new_n298), .B2(new_n287), .ZN(new_n302));
  OAI221_X1 g0102(.A(new_n290), .B1(G50), .B2(new_n291), .C1(new_n301), .C2(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n303), .A2(KEYINPUT9), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(KEYINPUT9), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n285), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n283), .A2(G200), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT76), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(KEYINPUT10), .ZN(new_n311));
  OR2_X1    g0111(.A1(new_n310), .A2(KEYINPUT10), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n309), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G169), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n283), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(new_n303), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT73), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n315), .A2(KEYINPUT73), .A3(new_n303), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n318), .B(new_n319), .C1(G179), .C2(new_n283), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n307), .A2(new_n310), .A3(KEYINPUT10), .A4(new_n308), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n313), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT75), .ZN(new_n324));
  XNOR2_X1  g0124(.A(new_n291), .B(new_n324), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n325), .A2(G77), .ZN(new_n326));
  INV_X1    g0126(.A(new_n294), .ZN(new_n327));
  OAI22_X1  g0127(.A1(new_n234), .A2(new_n223), .B1(new_n297), .B2(new_n327), .ZN(new_n328));
  XOR2_X1   g0128(.A(new_n328), .B(KEYINPUT74), .Z(new_n329));
  XOR2_X1   g0129(.A(KEYINPUT15), .B(G87), .Z(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n329), .B1(new_n296), .B2(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n326), .B1(new_n332), .B2(new_n287), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n325), .A2(new_n288), .A3(new_n289), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n334), .A2(new_n223), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n271), .A2(G232), .ZN(new_n338));
  INV_X1    g0138(.A(G107), .ZN(new_n339));
  OAI221_X1 g0139(.A(new_n338), .B1(new_n339), .B2(new_n262), .C1(new_n264), .C2(new_n211), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n261), .ZN(new_n341));
  INV_X1    g0141(.A(G179), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n277), .A2(G244), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n341), .A2(new_n342), .A3(new_n282), .A4(new_n343), .ZN(new_n344));
  AND3_X1   g0144(.A1(new_n341), .A2(new_n282), .A3(new_n343), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n337), .B(new_n344), .C1(new_n345), .C2(G169), .ZN(new_n346));
  AOI211_X1 g0146(.A(new_n326), .B(new_n335), .C1(new_n332), .C2(new_n287), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n341), .A2(G190), .A3(new_n282), .A4(new_n343), .ZN(new_n348));
  INV_X1    g0148(.A(G200), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n347), .B(new_n348), .C1(new_n345), .C2(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n323), .A2(new_n346), .A3(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(G1698), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n267), .B(new_n269), .C1(G226), .C2(new_n352), .ZN(new_n353));
  NOR2_X1   g0153(.A1(G223), .A2(G1698), .ZN(new_n354));
  OAI22_X1  g0154(.A1(new_n353), .A2(new_n354), .B1(new_n258), .B2(new_n213), .ZN(new_n355));
  OR2_X1    g0155(.A1(new_n281), .A2(KEYINPUT68), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n281), .A2(KEYINPUT68), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n355), .A2(new_n261), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(KEYINPUT79), .B1(new_n276), .B2(new_n227), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT79), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n260), .A2(new_n360), .A3(G232), .A4(new_n275), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  OAI21_X1  g0163(.A(KEYINPUT81), .B1(new_n363), .B2(G190), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n349), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT81), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n358), .A2(new_n366), .A3(new_n284), .A4(new_n362), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n364), .A2(new_n365), .A3(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n268), .A2(KEYINPUT77), .A3(G33), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n267), .ZN(new_n370));
  AOI21_X1  g0170(.A(KEYINPUT77), .B1(new_n268), .B2(G33), .ZN(new_n371));
  OAI211_X1 g0171(.A(KEYINPUT7), .B(new_n234), .C1(new_n370), .C2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT7), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n373), .B1(new_n262), .B2(G20), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(G68), .ZN(new_n376));
  XNOR2_X1  g0176(.A(G58), .B(G68), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n377), .A2(G20), .B1(G159), .B2(new_n294), .ZN(new_n378));
  AOI21_X1  g0178(.A(KEYINPUT16), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(KEYINPUT7), .B1(new_n262), .B2(G20), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n234), .A2(new_n270), .A3(new_n373), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n380), .A2(new_n381), .A3(G68), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n382), .A2(new_n378), .A3(KEYINPUT16), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n287), .ZN(new_n384));
  OAI21_X1  g0184(.A(KEYINPUT78), .B1(new_n379), .B2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n297), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(new_n289), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n291), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n389), .A2(new_n287), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n388), .A2(new_n390), .B1(new_n389), .B2(new_n297), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT16), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n210), .B1(new_n372), .B2(new_n374), .ZN(new_n393));
  INV_X1    g0193(.A(new_n378), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n392), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT78), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n395), .A2(new_n396), .A3(new_n287), .A4(new_n383), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n368), .A2(new_n385), .A3(new_n391), .A4(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT17), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AND2_X1   g0200(.A1(new_n385), .A2(new_n397), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n401), .A2(KEYINPUT17), .A3(new_n391), .A4(new_n368), .ZN(new_n402));
  AND3_X1   g0202(.A1(new_n358), .A2(new_n342), .A3(new_n362), .ZN(new_n403));
  AOI21_X1  g0203(.A(G169), .B1(new_n358), .B2(new_n362), .ZN(new_n404));
  OAI21_X1  g0204(.A(KEYINPUT80), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n363), .A2(new_n314), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT80), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n358), .A2(new_n342), .A3(new_n362), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n385), .A2(new_n391), .A3(new_n397), .ZN(new_n411));
  AND3_X1   g0211(.A1(new_n410), .A2(new_n411), .A3(KEYINPUT18), .ZN(new_n412));
  AOI21_X1  g0212(.A(KEYINPUT18), .B1(new_n410), .B2(new_n411), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n400), .B(new_n402), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  AND2_X1   g0215(.A1(G33), .A2(G97), .ZN(new_n416));
  NOR2_X1   g0216(.A1(G226), .A2(G1698), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n417), .B1(new_n227), .B2(G1698), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n416), .B1(new_n418), .B2(new_n262), .ZN(new_n419));
  OAI221_X1 g0219(.A(new_n282), .B1(new_n211), .B2(new_n276), .C1(new_n419), .C2(new_n260), .ZN(new_n420));
  XNOR2_X1  g0220(.A(new_n420), .B(KEYINPUT13), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(KEYINPUT14), .B1(new_n422), .B2(new_n314), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(G179), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT14), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n421), .A2(new_n425), .A3(G169), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n423), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  XNOR2_X1  g0227(.A(new_n291), .B(KEYINPUT75), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n428), .A2(KEYINPUT12), .A3(new_n210), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n389), .A2(KEYINPUT12), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n334), .A2(KEYINPUT12), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n430), .B1(new_n431), .B2(G68), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n294), .A2(G50), .ZN(new_n433));
  OAI221_X1 g0233(.A(new_n433), .B1(new_n204), .B2(G68), .C1(new_n296), .C2(new_n223), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n287), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n435), .A2(KEYINPUT11), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n435), .A2(KEYINPUT11), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n429), .B(new_n432), .C1(new_n436), .C2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n427), .A2(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n421), .A2(new_n284), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n440), .A2(new_n438), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n441), .B1(new_n349), .B2(new_n422), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n415), .A2(new_n439), .A3(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n351), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n262), .A2(G244), .A3(new_n352), .ZN(new_n446));
  NOR2_X1   g0246(.A1(KEYINPUT83), .A2(KEYINPUT4), .ZN(new_n447));
  OR2_X1    g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n270), .A2(new_n352), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n449), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n450));
  NAND2_X1  g0250(.A1(KEYINPUT83), .A2(KEYINPUT4), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n446), .A2(new_n447), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n448), .A2(new_n450), .A3(new_n451), .A4(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n261), .ZN(new_n454));
  INV_X1    g0254(.A(G45), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n455), .A2(G1), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n456), .B(KEYINPUT84), .C1(KEYINPUT5), .C2(new_n259), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n203), .B(G45), .C1(new_n259), .C2(KEYINPUT5), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT84), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  OR2_X1    g0261(.A1(KEYINPUT85), .A2(KEYINPUT5), .ZN(new_n462));
  NAND2_X1  g0262(.A1(KEYINPUT85), .A2(KEYINPUT5), .ZN(new_n463));
  AOI21_X1  g0263(.A(G41), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(G274), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n461), .A2(new_n466), .A3(new_n260), .ZN(new_n467));
  OAI211_X1 g0267(.A(G257), .B(new_n260), .C1(new_n464), .C2(new_n458), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n454), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n470), .A2(new_n349), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n291), .A2(G97), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n203), .A2(G33), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n390), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n475), .A2(new_n215), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  OR2_X1    g0277(.A1(new_n215), .A2(KEYINPUT6), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT82), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n215), .A2(new_n339), .A3(KEYINPUT6), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n479), .B1(new_n478), .B2(new_n480), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n339), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(new_n483), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n485), .A2(G107), .A3(new_n481), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n234), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n339), .B1(new_n372), .B2(new_n374), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n327), .A2(new_n223), .ZN(new_n489));
  NOR3_X1   g0289(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n473), .B(new_n477), .C1(new_n490), .C2(new_n288), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n469), .A2(new_n284), .ZN(new_n492));
  NOR3_X1   g0292(.A1(new_n471), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n470), .A2(new_n342), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n469), .A2(new_n314), .ZN(new_n495));
  AND3_X1   g0295(.A1(new_n494), .A2(new_n491), .A3(new_n495), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n325), .A2(new_n330), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n231), .A2(new_n233), .B1(new_n416), .B2(KEYINPUT19), .ZN(new_n499));
  NOR3_X1   g0299(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n500));
  OAI21_X1  g0300(.A(KEYINPUT87), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n232), .A2(G20), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n204), .A2(KEYINPUT64), .ZN(new_n503));
  OAI211_X1 g0303(.A(G33), .B(G97), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT19), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n234), .A2(new_n262), .A3(G68), .ZN(new_n507));
  INV_X1    g0307(.A(new_n500), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT87), .ZN(new_n509));
  XNOR2_X1  g0309(.A(KEYINPUT64), .B(G20), .ZN(new_n510));
  AND3_X1   g0310(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n508), .B(new_n509), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n501), .A2(new_n506), .A3(new_n507), .A4(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n498), .B1(new_n513), .B2(new_n287), .ZN(new_n514));
  INV_X1    g0314(.A(new_n475), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n330), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n224), .A2(G1698), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n262), .B(new_n517), .C1(G238), .C2(G1698), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G33), .A2(G116), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n260), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n465), .B1(new_n214), .B2(KEYINPUT86), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n456), .ZN(new_n522));
  OAI211_X1 g0322(.A(KEYINPUT86), .B(G250), .C1(new_n455), .C2(G1), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n261), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n520), .A2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n514), .A2(new_n516), .B1(new_n526), .B2(new_n314), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n342), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n526), .A2(G200), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n515), .A2(G87), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n525), .A2(G190), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n530), .A2(new_n514), .A3(new_n531), .A4(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n214), .A2(new_n352), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n216), .A2(G1698), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n267), .A2(new_n535), .A3(new_n269), .A4(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(G294), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n537), .B1(new_n258), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n261), .ZN(new_n540));
  OAI211_X1 g0340(.A(G264), .B(new_n260), .C1(new_n464), .C2(new_n458), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n467), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n314), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n467), .A2(new_n540), .A3(new_n342), .A4(new_n541), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n234), .A2(new_n262), .A3(G87), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT22), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n547), .A2(KEYINPUT88), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(new_n548), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n234), .A2(new_n262), .A3(new_n550), .A4(G87), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(KEYINPUT23), .A2(G107), .ZN(new_n553));
  AOI21_X1  g0353(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n553), .B1(new_n554), .B2(G20), .ZN(new_n555));
  NOR2_X1   g0355(.A1(KEYINPUT23), .A2(G107), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n555), .B1(new_n510), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n552), .A2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT24), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n552), .A2(KEYINPUT24), .A3(new_n557), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n560), .A2(new_n287), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n515), .A2(G107), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n389), .A2(new_n339), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT89), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n564), .A2(new_n565), .A3(KEYINPUT25), .ZN(new_n566));
  XOR2_X1   g0366(.A(KEYINPUT89), .B(KEYINPUT25), .Z(new_n567));
  NOR2_X1   g0367(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(new_n568), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n563), .A2(KEYINPUT90), .A3(new_n566), .A4(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT90), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n566), .B1(new_n475), .B2(new_n339), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n571), .B1(new_n572), .B2(new_n568), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n545), .B1(new_n562), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n534), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n325), .A2(G116), .A3(new_n288), .A4(new_n474), .ZN(new_n577));
  INV_X1    g0377(.A(G116), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n428), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(G33), .A2(G283), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n258), .A2(G97), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n234), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n286), .A2(new_n235), .B1(G20), .B2(new_n578), .ZN(new_n583));
  AND3_X1   g0383(.A1(new_n582), .A2(KEYINPUT20), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(KEYINPUT20), .B1(new_n582), .B2(new_n583), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n577), .B(new_n579), .C1(new_n584), .C2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(G264), .A2(G1698), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n262), .B(new_n587), .C1(new_n216), .C2(G1698), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n588), .B(new_n261), .C1(G303), .C2(new_n262), .ZN(new_n589));
  OAI211_X1 g0389(.A(G270), .B(new_n260), .C1(new_n464), .C2(new_n458), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n589), .A2(new_n467), .A3(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n591), .A2(new_n284), .ZN(new_n592));
  AOI211_X1 g0392(.A(new_n586), .B(new_n592), .C1(G200), .C2(new_n591), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n586), .A2(G169), .A3(new_n591), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT21), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n591), .A2(new_n342), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n586), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n586), .A2(new_n591), .A3(KEYINPUT21), .A4(G169), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n596), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n593), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n542), .A2(G200), .ZN(new_n602));
  AND2_X1   g0402(.A1(new_n540), .A2(new_n541), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n603), .A2(G190), .A3(new_n467), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n562), .A2(new_n574), .A3(new_n602), .A4(new_n604), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n497), .A2(new_n576), .A3(new_n601), .A4(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n445), .A2(new_n606), .ZN(G372));
  INV_X1    g0407(.A(new_n442), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n439), .B1(new_n608), .B2(new_n346), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n400), .A2(new_n402), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT95), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n611), .B1(new_n412), .B2(new_n413), .ZN(new_n612));
  INV_X1    g0412(.A(new_n413), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n410), .A2(new_n411), .A3(KEYINPUT18), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n613), .A2(KEYINPUT95), .A3(new_n614), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n609), .A2(new_n610), .B1(new_n612), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n313), .A2(new_n321), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n320), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  XNOR2_X1  g0419(.A(KEYINPUT94), .B(KEYINPUT26), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n496), .A2(new_n533), .A3(new_n620), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n605), .B1(new_n600), .B2(new_n575), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n494), .A2(new_n491), .A3(new_n495), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n491), .A2(new_n492), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n625), .B1(new_n349), .B2(new_n470), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT92), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT91), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n513), .A2(new_n287), .ZN(new_n630));
  INV_X1    g0430(.A(new_n498), .ZN(new_n631));
  AND4_X1   g0431(.A1(new_n629), .A2(new_n630), .A3(new_n631), .A4(new_n531), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n629), .B1(new_n514), .B2(new_n531), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n628), .B(new_n530), .C1(new_n632), .C2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n532), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n630), .A2(new_n631), .A3(new_n531), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(KEYINPUT91), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n514), .A2(new_n629), .A3(new_n531), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n628), .B1(new_n639), .B2(new_n530), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n529), .B1(new_n635), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(KEYINPUT93), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT93), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n643), .B(new_n529), .C1(new_n635), .C2(new_n640), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n627), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n621), .B1(new_n645), .B2(KEYINPUT26), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(new_n529), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n619), .B1(new_n445), .B2(new_n648), .ZN(G369));
  INV_X1    g0449(.A(G13), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n510), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n203), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(KEYINPUT27), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT27), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n651), .A2(new_n654), .A3(new_n203), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n653), .A2(G213), .A3(G343), .A4(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT96), .ZN(new_n657));
  XNOR2_X1  g0457(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n586), .ZN(new_n659));
  MUX2_X1   g0459(.A(new_n600), .B(new_n601), .S(new_n659), .Z(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(G330), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n562), .A2(new_n574), .ZN(new_n662));
  INV_X1    g0462(.A(new_n658), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n605), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n575), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n575), .A2(new_n663), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n661), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n600), .A2(new_n663), .ZN(new_n671));
  XOR2_X1   g0471(.A(new_n671), .B(KEYINPUT97), .Z(new_n672));
  INV_X1    g0472(.A(new_n668), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(new_n667), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n670), .A2(new_n676), .ZN(G399));
  INV_X1    g0477(.A(new_n207), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(G41), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(G1), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n500), .A2(new_n578), .ZN(new_n682));
  OAI22_X1  g0482(.A1(new_n681), .A2(new_n682), .B1(new_n238), .B2(new_n680), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n683), .B(KEYINPUT28), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n658), .B1(new_n646), .B2(new_n529), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT29), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n493), .B1(new_n623), .B2(new_n622), .ZN(new_n688));
  INV_X1    g0488(.A(new_n644), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n530), .B1(new_n632), .B2(new_n633), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(KEYINPUT92), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n691), .A2(new_n532), .A3(new_n634), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n643), .B1(new_n692), .B2(new_n529), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n688), .B1(new_n689), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(KEYINPUT99), .B1(new_n694), .B2(new_n496), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT99), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n645), .A2(new_n696), .A3(new_n623), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT26), .ZN(new_n699));
  AOI211_X1 g0499(.A(new_n699), .B(new_n623), .C1(new_n642), .C2(new_n644), .ZN(new_n700));
  INV_X1    g0500(.A(new_n534), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n620), .B1(new_n496), .B2(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n529), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n658), .B1(new_n698), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n687), .B1(new_n705), .B2(new_n686), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n454), .A2(new_n525), .A3(new_n467), .A4(new_n468), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n597), .A2(new_n603), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT30), .ZN(new_n709));
  OR3_X1    g0509(.A1(new_n707), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n709), .B1(new_n707), .B2(new_n708), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n591), .A2(new_n342), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n469), .A2(new_n526), .A3(new_n542), .A4(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n710), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(new_n658), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT31), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT98), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n717), .B(new_n718), .ZN(new_n719));
  OAI22_X1  g0519(.A1(new_n606), .A2(new_n658), .B1(new_n716), .B2(new_n715), .ZN(new_n720));
  OAI21_X1  g0520(.A(G330), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n706), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n684), .B1(new_n723), .B2(G1), .ZN(G364));
  NOR2_X1   g0524(.A1(G13), .A2(G33), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  OR3_X1    g0526(.A1(new_n660), .A2(G20), .A3(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n678), .A2(new_n262), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n239), .A2(new_n455), .ZN(new_n729));
  OAI211_X1 g0529(.A(new_n728), .B(new_n729), .C1(new_n256), .C2(new_n455), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n207), .A2(G355), .A3(new_n262), .ZN(new_n731));
  OAI211_X1 g0531(.A(new_n730), .B(new_n731), .C1(G116), .C2(new_n207), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n726), .A2(G20), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n235), .B1(G20), .B2(new_n314), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n681), .B1(G45), .B2(new_n651), .ZN(new_n737));
  NOR4_X1   g0537(.A1(new_n234), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  XOR2_X1   g0539(.A(KEYINPUT101), .B(G159), .Z(new_n740));
  NOR3_X1   g0540(.A1(new_n739), .A2(KEYINPUT32), .A3(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n349), .A2(G179), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n742), .A2(G20), .A3(G190), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n234), .A2(new_n342), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G190), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(G200), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  OAI221_X1 g0547(.A(new_n262), .B1(new_n213), .B2(new_n743), .C1(new_n747), .C2(new_n226), .ZN(new_n748));
  NOR3_X1   g0548(.A1(new_n284), .A2(G179), .A3(G200), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n234), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  AOI211_X1 g0551(.A(new_n741), .B(new_n748), .C1(G97), .C2(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(KEYINPUT32), .B1(new_n739), .B2(new_n740), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n510), .A2(new_n284), .A3(new_n742), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G107), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n744), .A2(new_n284), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(new_n349), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n756), .B1(new_n759), .B2(new_n210), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n744), .A2(new_n284), .A3(new_n349), .ZN(new_n761));
  AND2_X1   g0561(.A1(new_n761), .A2(KEYINPUT100), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n761), .A2(KEYINPUT100), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n760), .B1(new_n765), .B2(G77), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n752), .A2(new_n753), .A3(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n745), .A2(new_n349), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n767), .B1(G50), .B2(new_n768), .ZN(new_n769));
  XOR2_X1   g0569(.A(KEYINPUT33), .B(G317), .Z(new_n770));
  NOR2_X1   g0570(.A1(new_n759), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(G322), .ZN(new_n772));
  INV_X1    g0572(.A(G303), .ZN(new_n773));
  OAI22_X1  g0573(.A1(new_n747), .A2(new_n772), .B1(new_n773), .B2(new_n743), .ZN(new_n774));
  AOI211_X1 g0574(.A(new_n771), .B(new_n774), .C1(G283), .C2(new_n755), .ZN(new_n775));
  AND2_X1   g0575(.A1(new_n738), .A2(G329), .ZN(new_n776));
  AOI211_X1 g0576(.A(new_n262), .B(new_n776), .C1(G326), .C2(new_n768), .ZN(new_n777));
  OAI211_X1 g0577(.A(new_n775), .B(new_n777), .C1(new_n538), .C2(new_n750), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n778), .B1(G311), .B2(new_n765), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n734), .B1(new_n769), .B2(new_n779), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n727), .A2(new_n736), .A3(new_n737), .A4(new_n780), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n660), .B(G330), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n781), .B1(new_n737), .B2(new_n782), .ZN(G396));
  NAND2_X1  g0583(.A1(new_n337), .A2(new_n658), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n346), .A2(new_n350), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(KEYINPUT103), .ZN(new_n786));
  INV_X1    g0586(.A(KEYINPUT103), .ZN(new_n787));
  NAND4_X1  g0587(.A1(new_n346), .A2(new_n350), .A3(new_n787), .A4(new_n784), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n621), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n791), .B1(new_n694), .B2(new_n699), .ZN(new_n792));
  INV_X1    g0592(.A(new_n529), .ZN(new_n793));
  OAI211_X1 g0593(.A(new_n663), .B(new_n790), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(KEYINPUT104), .ZN(new_n795));
  INV_X1    g0595(.A(KEYINPUT104), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n796), .B1(new_n685), .B2(new_n790), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n346), .A2(new_n663), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n798), .B1(new_n786), .B2(new_n788), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n795), .A2(new_n797), .B1(new_n685), .B2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n721), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(KEYINPUT105), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n737), .B1(new_n801), .B2(new_n721), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n764), .A2(new_n578), .B1(new_n215), .B2(new_n750), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n746), .A2(G294), .B1(G311), .B2(new_n738), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(new_n213), .B2(new_n754), .ZN(new_n808));
  INV_X1    g0608(.A(G283), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n759), .A2(new_n809), .ZN(new_n810));
  NOR4_X1   g0610(.A1(new_n806), .A2(new_n808), .A3(new_n262), .A4(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n768), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n811), .B1(new_n339), .B2(new_n743), .C1(new_n773), .C2(new_n812), .ZN(new_n813));
  XOR2_X1   g0613(.A(KEYINPUT102), .B(G143), .Z(new_n814));
  NAND2_X1  g0614(.A1(new_n746), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(G150), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n815), .B1(new_n759), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n764), .A2(new_n740), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n817), .B(new_n818), .C1(G137), .C2(new_n768), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(KEYINPUT34), .Z(new_n820));
  NOR2_X1   g0620(.A1(new_n754), .A2(new_n210), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n270), .B(new_n821), .C1(G58), .C2(new_n751), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n820), .B(new_n822), .C1(new_n221), .C2(new_n743), .ZN(new_n823));
  INV_X1    g0623(.A(G132), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n739), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n813), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(new_n734), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n734), .A2(new_n725), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n223), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n799), .A2(new_n725), .ZN(new_n830));
  NAND4_X1  g0630(.A1(new_n827), .A2(new_n737), .A3(new_n829), .A4(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n805), .A2(new_n831), .ZN(G384));
  AOI21_X1  g0632(.A(KEYINPUT16), .B1(new_n382), .B2(new_n378), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n391), .B1(new_n384), .B2(new_n833), .ZN(new_n834));
  XOR2_X1   g0634(.A(new_n834), .B(KEYINPUT107), .Z(new_n835));
  NAND3_X1  g0635(.A1(new_n653), .A2(G213), .A3(new_n655), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n414), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(KEYINPUT108), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT108), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n414), .A2(new_n840), .A3(new_n837), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n836), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n411), .B1(new_n410), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n398), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT37), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n410), .A2(new_n843), .ZN(new_n848));
  OAI211_X1 g0648(.A(KEYINPUT37), .B(new_n398), .C1(new_n835), .C2(new_n848), .ZN(new_n849));
  NAND4_X1  g0649(.A1(new_n842), .A2(KEYINPUT38), .A3(new_n847), .A4(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT39), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT38), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT109), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n846), .B1(new_n844), .B2(new_n853), .ZN(new_n854));
  XOR2_X1   g0654(.A(new_n854), .B(new_n845), .Z(new_n855));
  NAND2_X1  g0655(.A1(new_n411), .A2(new_n843), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n615), .A2(new_n612), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n856), .B1(new_n857), .B2(new_n610), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n852), .B1(new_n855), .B2(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n850), .A2(new_n851), .A3(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  AND3_X1   g0661(.A1(new_n414), .A2(new_n840), .A3(new_n837), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n840), .B1(new_n414), .B2(new_n837), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n847), .B(new_n849), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n852), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n851), .B1(new_n865), .B2(new_n850), .ZN(new_n866));
  OAI21_X1  g0666(.A(KEYINPUT110), .B1(new_n861), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n865), .A2(new_n850), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(KEYINPUT39), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT110), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n869), .A2(new_n870), .A3(new_n860), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n867), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n439), .A2(new_n658), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n346), .A2(new_n658), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n876), .B1(new_n795), .B2(new_n797), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n438), .A2(new_n658), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT106), .ZN(new_n879));
  XNOR2_X1  g0679(.A(new_n878), .B(new_n879), .ZN(new_n880));
  AND3_X1   g0680(.A1(new_n439), .A2(new_n442), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n880), .B1(new_n439), .B2(new_n442), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n877), .A2(new_n868), .A3(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n615), .A2(new_n612), .A3(new_n836), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n874), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n618), .B1(new_n706), .B2(new_n444), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n887), .B(new_n888), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n717), .B(KEYINPUT111), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n715), .A2(new_n716), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n626), .A2(new_n601), .A3(new_n623), .A4(new_n605), .ZN(new_n892));
  INV_X1    g0692(.A(new_n576), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n891), .B1(new_n894), .B2(new_n663), .ZN(new_n895));
  AOI211_X1 g0695(.A(new_n799), .B(new_n883), .C1(new_n890), .C2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n868), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT40), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n850), .A2(new_n859), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n896), .A2(new_n900), .A3(KEYINPUT40), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT111), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n717), .B(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n444), .B1(new_n720), .B2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n902), .B(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(G330), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n889), .B(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n203), .B2(new_n651), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n484), .A2(new_n486), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n578), .B1(new_n912), .B2(KEYINPUT35), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n913), .B(new_n237), .C1(KEYINPUT35), .C2(new_n912), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n914), .B(KEYINPUT36), .ZN(new_n915));
  OAI21_X1  g0715(.A(G77), .B1(new_n226), .B2(new_n210), .ZN(new_n916));
  OAI22_X1  g0716(.A1(new_n916), .A2(new_n238), .B1(G50), .B2(new_n210), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n917), .A2(G1), .A3(new_n650), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n910), .A2(new_n915), .A3(new_n918), .ZN(G367));
  INV_X1    g0719(.A(new_n674), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n491), .A2(new_n658), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n497), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n496), .A2(new_n658), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n920), .A2(new_n924), .ZN(new_n925));
  XOR2_X1   g0725(.A(KEYINPUT112), .B(KEYINPUT42), .Z(new_n926));
  XNOR2_X1  g0726(.A(new_n925), .B(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n623), .B1(new_n922), .B2(new_n665), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n663), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n689), .A2(new_n693), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n639), .A2(new_n663), .ZN(new_n932));
  MUX2_X1   g0732(.A(new_n931), .B(new_n529), .S(new_n932), .Z(new_n933));
  INV_X1    g0733(.A(KEYINPUT43), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n930), .A2(new_n935), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n936), .B(KEYINPUT113), .Z(new_n937));
  NOR2_X1   g0737(.A1(new_n933), .A2(new_n934), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n930), .A2(new_n935), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n924), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n670), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n940), .B(new_n942), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n679), .B(KEYINPUT41), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n675), .A2(new_n941), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT45), .ZN(new_n947));
  OAI21_X1  g0747(.A(KEYINPUT44), .B1(new_n676), .B2(new_n924), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT44), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n675), .A2(new_n941), .A3(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n947), .A2(new_n948), .A3(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n951), .A2(new_n669), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n952), .B(KEYINPUT116), .Z(new_n953));
  NAND2_X1  g0753(.A1(new_n951), .A2(new_n669), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(KEYINPUT114), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT115), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n672), .B2(new_n673), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(new_n661), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(new_n920), .ZN(new_n959));
  AND2_X1   g0759(.A1(new_n723), .A2(new_n959), .ZN(new_n960));
  OR2_X1    g0760(.A1(new_n954), .A2(KEYINPUT114), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n953), .A2(new_n955), .A3(new_n960), .A4(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n945), .B1(new_n962), .B2(new_n723), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n203), .B1(new_n651), .B2(G45), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n943), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n933), .A2(new_n733), .ZN(new_n967));
  INV_X1    g0767(.A(G137), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n739), .A2(new_n968), .B1(new_n210), .B2(new_n750), .ZN(new_n969));
  OAI221_X1 g0769(.A(new_n262), .B1(new_n223), .B2(new_n754), .C1(new_n759), .C2(new_n740), .ZN(new_n970));
  AOI211_X1 g0770(.A(new_n969), .B(new_n970), .C1(G150), .C2(new_n746), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n765), .A2(G50), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n768), .A2(new_n814), .ZN(new_n973));
  INV_X1    g0773(.A(new_n743), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(G58), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n971), .A2(new_n972), .A3(new_n973), .A4(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n747), .A2(new_n773), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n768), .A2(G311), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n738), .A2(G317), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n755), .A2(G97), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  AOI211_X1 g0781(.A(new_n977), .B(new_n981), .C1(G294), .C2(new_n758), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n751), .A2(G107), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n765), .A2(G283), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n974), .A2(G116), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT46), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n262), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n982), .A2(new_n983), .A3(new_n984), .A4(new_n987), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n985), .A2(new_n986), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n976), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT47), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n734), .ZN(new_n992));
  INV_X1    g0792(.A(new_n728), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n735), .B1(new_n207), .B2(new_n331), .C1(new_n248), .C2(new_n993), .ZN(new_n994));
  NAND4_X1  g0794(.A1(new_n967), .A2(new_n737), .A3(new_n992), .A4(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n966), .A2(new_n995), .ZN(G387));
  NOR2_X1   g0796(.A1(new_n750), .A2(new_n331), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n739), .A2(new_n816), .ZN(new_n998));
  AOI211_X1 g0798(.A(new_n997), .B(new_n998), .C1(new_n386), .C2(new_n758), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n768), .A2(G159), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n999), .B(new_n1000), .C1(new_n221), .C2(new_n747), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(new_n765), .B2(G68), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n974), .A2(G77), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n1002), .A2(new_n262), .A3(new_n980), .A4(new_n1003), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(G311), .A2(new_n758), .B1(new_n746), .B2(G317), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n1005), .B1(new_n772), .B2(new_n812), .C1(new_n764), .C2(new_n773), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT48), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n1007), .B1(new_n809), .B2(new_n750), .C1(new_n538), .C2(new_n743), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT49), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n755), .A2(G116), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n738), .A2(G326), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1010), .A2(new_n270), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  AND2_X1   g0813(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1004), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(new_n734), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n386), .A2(new_n221), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT50), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n210), .A2(new_n223), .ZN(new_n1019));
  NOR4_X1   g0819(.A1(new_n1018), .A2(G45), .A3(new_n1019), .A4(new_n682), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n245), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n728), .B1(new_n1021), .B2(new_n455), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n207), .A2(new_n262), .A3(new_n682), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1020), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n207), .A2(G107), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n735), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1016), .A2(new_n737), .A3(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(new_n668), .B2(new_n733), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(new_n959), .B2(new_n965), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n679), .B1(new_n723), .B2(new_n959), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1029), .B1(new_n960), .B2(new_n1030), .ZN(G393));
  AND2_X1   g0831(.A1(new_n953), .A2(new_n954), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n679), .B(new_n962), .C1(new_n1032), .C2(new_n960), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n941), .A2(new_n733), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n758), .A2(G303), .B1(G322), .B2(new_n738), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n756), .B(new_n1035), .C1(new_n764), .C2(new_n538), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(G311), .A2(new_n746), .B1(new_n768), .B2(G317), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT52), .Z(new_n1038));
  OAI211_X1 g0838(.A(new_n1038), .B(new_n270), .C1(new_n809), .C2(new_n743), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n1036), .B(new_n1039), .C1(G116), .C2(new_n751), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n765), .A2(new_n386), .B1(G50), .B2(new_n758), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n738), .A2(new_n814), .B1(new_n755), .B2(G87), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n751), .A2(G77), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(G150), .A2(new_n768), .B1(new_n746), .B2(G159), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n1045), .A2(KEYINPUT51), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n743), .A2(new_n210), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n262), .B1(new_n1045), .B2(KEYINPUT51), .ZN(new_n1048));
  NOR4_X1   g0848(.A1(new_n1044), .A2(new_n1046), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n734), .B1(new_n1040), .B2(new_n1049), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n735), .B1(new_n215), .B2(new_n207), .C1(new_n253), .C2(new_n993), .ZN(new_n1051));
  AND4_X1   g0851(.A1(new_n737), .A2(new_n1034), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(new_n1032), .B2(new_n965), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1033), .A2(new_n1053), .ZN(G390));
  AND2_X1   g0854(.A1(new_n867), .A2(new_n871), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(new_n725), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n828), .A2(new_n297), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n339), .A2(new_n759), .B1(new_n747), .B2(new_n578), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n821), .B(new_n1058), .C1(G283), .C2(new_n768), .ZN(new_n1059));
  AND2_X1   g0859(.A1(new_n1059), .A2(new_n1043), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n1060), .B1(new_n215), .B2(new_n764), .C1(new_n538), .C2(new_n739), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n262), .B(new_n1061), .C1(G87), .C2(new_n974), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n738), .A2(G125), .B1(new_n751), .B2(G159), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n1063), .B1(new_n221), .B2(new_n754), .C1(new_n759), .C2(new_n968), .ZN(new_n1064));
  XOR2_X1   g0864(.A(KEYINPUT54), .B(G143), .Z(new_n1065));
  INV_X1    g0865(.A(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n764), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n768), .A2(G128), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1068), .B(new_n262), .C1(new_n747), .C2(new_n824), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n974), .A2(G150), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT53), .ZN(new_n1071));
  NOR4_X1   g0871(.A1(new_n1064), .A2(new_n1067), .A3(new_n1069), .A4(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n734), .B1(new_n1062), .B2(new_n1072), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1056), .A2(new_n737), .A3(new_n1057), .A4(new_n1073), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT117), .Z(new_n1075));
  NAND2_X1  g0875(.A1(new_n695), .A2(new_n697), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n663), .B(new_n790), .C1(new_n1076), .C2(new_n703), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n876), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n884), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n873), .B1(new_n850), .B2(new_n859), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NOR3_X1   g0881(.A1(new_n721), .A2(new_n799), .A3(new_n883), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n873), .B1(new_n877), .B2(new_n884), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1081), .B(new_n1082), .C1(new_n1083), .C2(new_n872), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n873), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n794), .A2(KEYINPUT104), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n685), .A2(new_n796), .A3(new_n790), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n875), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1085), .B1(new_n1088), .B2(new_n883), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n1055), .A2(new_n1089), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n799), .B1(new_n890), .B2(new_n895), .ZN(new_n1091));
  AND3_X1   g0891(.A1(new_n1091), .A2(G330), .A3(new_n884), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1084), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n884), .B1(new_n722), .B2(new_n800), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1094), .A2(new_n1092), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n884), .B1(new_n1091), .B2(G330), .ZN(new_n1096));
  OR2_X1    g0896(.A1(new_n1082), .A2(new_n1096), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n1095), .A2(new_n1088), .B1(new_n1097), .B2(new_n1078), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n906), .A2(G330), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1098), .A2(new_n888), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1093), .A2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1081), .B1(new_n1083), .B2(new_n872), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1092), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1105), .A2(new_n1084), .A3(new_n1100), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1102), .A2(new_n679), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1093), .A2(new_n965), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1075), .A2(new_n1107), .A3(new_n1108), .ZN(G378));
  OAI211_X1 g0909(.A(new_n800), .B(new_n884), .C1(new_n904), .C2(new_n720), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(new_n865), .B2(new_n850), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n901), .B(G330), .C1(new_n1111), .C2(KEYINPUT40), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n322), .A2(KEYINPUT119), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT119), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n313), .A2(new_n321), .A3(new_n320), .A4(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n303), .A2(new_n843), .ZN(new_n1118));
  AND3_X1   g0918(.A1(new_n1115), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1118), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1114), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1118), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1115), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1124), .A2(new_n1113), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1121), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1112), .A2(new_n1127), .ZN(new_n1128));
  AND2_X1   g0928(.A1(new_n1121), .A2(new_n1126), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1129), .A2(new_n899), .A3(G330), .A4(new_n901), .ZN(new_n1130));
  AND2_X1   g0930(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n887), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1133), .A2(new_n885), .A3(new_n874), .A4(new_n886), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT121), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1132), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  AND2_X1   g0936(.A1(new_n874), .A2(new_n886), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1137), .A2(KEYINPUT121), .A3(new_n885), .A4(new_n1133), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1136), .A2(KEYINPUT57), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT120), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1100), .B1(new_n1105), .B2(new_n1084), .ZN(new_n1141));
  AND2_X1   g0941(.A1(new_n888), .A2(new_n1099), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1140), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1102), .A2(KEYINPUT120), .A3(new_n1142), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1139), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(KEYINPUT122), .B1(new_n1146), .B2(new_n680), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n1136), .A2(KEYINPUT57), .A3(new_n1138), .ZN(new_n1148));
  AOI21_X1  g0948(.A(KEYINPUT120), .B1(new_n1102), .B2(new_n1142), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n1140), .B(new_n1143), .C1(new_n1093), .C2(new_n1101), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1148), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT122), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1151), .A2(new_n1152), .A3(new_n679), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1154), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT57), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1147), .A2(new_n1153), .A3(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1129), .A2(new_n725), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n828), .A2(new_n221), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n210), .A2(new_n750), .B1(new_n754), .B2(new_n226), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(G97), .A2(new_n758), .B1(new_n768), .B2(G116), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1162), .B1(new_n339), .B2(new_n747), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n1161), .B(new_n1163), .C1(new_n330), .C2(new_n765), .ZN(new_n1164));
  AOI21_X1  g0964(.A(G41), .B1(new_n738), .B2(G283), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1164), .A2(new_n270), .A3(new_n1003), .A4(new_n1165), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1166), .B(KEYINPUT58), .ZN(new_n1167));
  AOI21_X1  g0967(.A(G41), .B1(KEYINPUT3), .B2(G33), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n759), .A2(new_n824), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(G125), .A2(new_n768), .B1(new_n746), .B2(G128), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n1170), .B1(new_n816), .B2(new_n750), .C1(new_n743), .C2(new_n1066), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1169), .B(new_n1171), .C1(G137), .C2(new_n765), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT59), .ZN(new_n1173));
  AOI21_X1  g0973(.A(G33), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(G41), .B1(new_n738), .B2(G124), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1174), .B(new_n1175), .C1(new_n754), .C2(new_n740), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n1167), .B1(G50), .B2(new_n1168), .C1(new_n1176), .C2(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1178), .B(KEYINPUT118), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(new_n734), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1159), .A2(new_n737), .A3(new_n1160), .A4(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(new_n1154), .B2(new_n965), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1158), .A2(new_n1183), .ZN(G375));
  NOR2_X1   g0984(.A1(new_n1142), .A2(new_n1098), .ZN(new_n1185));
  OR3_X1    g0985(.A1(new_n1185), .A2(new_n1101), .A3(new_n945), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n578), .A2(new_n759), .B1(new_n747), .B2(new_n809), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1187), .A2(new_n997), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1188), .B1(new_n538), .B2(new_n812), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(G97), .B2(new_n974), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n1190), .B1(new_n339), .B2(new_n764), .C1(new_n773), .C2(new_n739), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n262), .B(new_n1191), .C1(G77), .C2(new_n755), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n747), .A2(new_n968), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n738), .A2(G128), .B1(G159), .B2(new_n974), .ZN(new_n1194));
  XOR2_X1   g0994(.A(new_n1194), .B(KEYINPUT123), .Z(new_n1195));
  OAI221_X1 g0995(.A(new_n262), .B1(new_n226), .B2(new_n754), .C1(new_n759), .C2(new_n1066), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n764), .A2(new_n816), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n750), .A2(new_n221), .ZN(new_n1198));
  OR4_X1    g0998(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .A4(new_n1198), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n1193), .B(new_n1199), .C1(G132), .C2(new_n768), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n734), .B1(new_n1192), .B2(new_n1200), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1201), .B(new_n737), .C1(new_n726), .C2(new_n884), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(new_n210), .B2(new_n828), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n1098), .B2(new_n965), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1186), .A2(new_n1204), .ZN(G381));
  XNOR2_X1  g1005(.A(G378), .B(KEYINPUT124), .ZN(new_n1206));
  AND3_X1   g1006(.A1(new_n1158), .A2(new_n1183), .A3(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(G384), .ZN(new_n1208));
  INV_X1    g1008(.A(G381), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n966), .A2(new_n995), .A3(new_n1053), .A4(new_n1033), .ZN(new_n1210));
  NOR3_X1   g1010(.A1(new_n1210), .A2(G396), .A3(G393), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .A4(new_n1211), .ZN(G407));
  INV_X1    g1012(.A(G213), .ZN(new_n1213));
  INV_X1    g1013(.A(G343), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1213), .B1(new_n1207), .B2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(G407), .ZN(G409));
  NAND2_X1  g1016(.A1(G387), .A2(G390), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT125), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1217), .A2(new_n1218), .A3(new_n1210), .ZN(new_n1219));
  XOR2_X1   g1019(.A(G393), .B(G396), .Z(new_n1220));
  OR2_X1    g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1213), .A2(G343), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1158), .A2(G378), .A3(new_n1183), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1136), .A2(new_n965), .A3(new_n1138), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1181), .B(new_n1226), .C1(new_n1155), .C2(new_n945), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1206), .A2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1224), .B1(new_n1225), .B2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1185), .A2(KEYINPUT60), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1230), .A2(new_n679), .A3(new_n1100), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1185), .A2(KEYINPUT60), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1204), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  OR2_X1    g1033(.A1(new_n1233), .A2(new_n1208), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  AND2_X1   g1035(.A1(new_n1233), .A2(new_n1208), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1229), .A2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(KEYINPUT62), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT61), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT62), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1229), .A2(new_n1241), .A3(new_n1237), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1239), .A2(new_n1240), .A3(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1224), .A2(G2897), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1237), .A2(new_n1244), .ZN(new_n1245));
  OAI211_X1 g1045(.A(G2897), .B(new_n1224), .C1(new_n1235), .C2(new_n1236), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1229), .A2(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1223), .B1(new_n1243), .B2(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1221), .A2(new_n1240), .A3(new_n1222), .ZN(new_n1250));
  OAI21_X1  g1050(.A(KEYINPUT63), .B1(new_n1229), .B2(new_n1247), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1250), .B1(new_n1251), .B2(new_n1238), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1225), .A2(new_n1228), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1224), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1253), .A2(KEYINPUT63), .A3(new_n1237), .A4(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(KEYINPUT126), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT126), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1229), .A2(new_n1257), .A3(KEYINPUT63), .A4(new_n1237), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1256), .A2(new_n1258), .ZN(new_n1259));
  AND3_X1   g1059(.A1(new_n1252), .A2(new_n1259), .A3(KEYINPUT127), .ZN(new_n1260));
  AOI21_X1  g1060(.A(KEYINPUT127), .B1(new_n1252), .B2(new_n1259), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1249), .B1(new_n1260), .B2(new_n1261), .ZN(G405));
  NAND2_X1  g1062(.A1(G375), .A2(new_n1206), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n1225), .ZN(new_n1264));
  XNOR2_X1  g1064(.A(new_n1264), .B(new_n1237), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(new_n1265), .B(new_n1223), .ZN(G402));
endmodule


