//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 0 0 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 0 0 1 1 0 1 1 0 0 1 1 0 1 1 1 0 1 0 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 0 0 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:48 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n545, new_n547, new_n548, new_n549, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n612, new_n614, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1180, new_n1181, new_n1182, new_n1183, new_n1185;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT65), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  OAI211_X1 g036(.A(G137), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G101), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g041(.A(G125), .B1(new_n460), .B2(new_n461), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI211_X1 g044(.A(KEYINPUT66), .B(G125), .C1(new_n460), .C2(new_n461), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(KEYINPUT67), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT67), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(G113), .A3(G2104), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n469), .A2(new_n470), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n466), .B1(new_n476), .B2(G2105), .ZN(G160));
  NOR2_X1   g052(.A1(new_n460), .A2(new_n461), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n478), .A2(new_n459), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  MUX2_X1   g057(.A(G100), .B(G112), .S(G2105), .Z(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G2104), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n480), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  OAI211_X1 g061(.A(G138), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  XNOR2_X1  g066(.A(KEYINPUT68), .B(G114), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n491), .B1(new_n492), .B2(new_n459), .ZN(new_n493));
  XNOR2_X1  g068(.A(KEYINPUT3), .B(G2104), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .A3(G138), .A4(new_n459), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n494), .A2(G126), .A3(G2105), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n489), .A2(new_n493), .A3(new_n495), .A4(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  INV_X1    g073(.A(KEYINPUT5), .ZN(new_n499));
  INV_X1    g074(.A(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n503), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g081(.A(KEYINPUT6), .B(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G88), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G50), .ZN(new_n511));
  OAI22_X1  g086(.A1(new_n508), .A2(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n506), .A2(new_n512), .ZN(G166));
  INV_X1    g088(.A(new_n510), .ZN(new_n514));
  NAND3_X1  g089(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(KEYINPUT7), .ZN(new_n516));
  OR2_X1    g091(.A1(new_n515), .A2(KEYINPUT7), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n514), .A2(G51), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AND2_X1   g093(.A1(new_n507), .A2(G89), .ZN(new_n519));
  AND2_X1   g094(.A1(G63), .A2(G651), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n503), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n518), .A2(new_n521), .ZN(G286));
  INV_X1    g097(.A(G286), .ZN(G168));
  INV_X1    g098(.A(G90), .ZN(new_n524));
  INV_X1    g099(.A(G52), .ZN(new_n525));
  OAI22_X1  g100(.A1(new_n508), .A2(new_n524), .B1(new_n510), .B2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(new_n502), .ZN(new_n527));
  NOR2_X1   g102(.A1(KEYINPUT5), .A2(G543), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(G64), .ZN(new_n530));
  INV_X1    g105(.A(G77), .ZN(new_n531));
  OAI22_X1  g106(.A1(new_n529), .A2(new_n530), .B1(new_n531), .B2(new_n500), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n532), .A2(KEYINPUT69), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n505), .B1(new_n532), .B2(KEYINPUT69), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n526), .B1(new_n533), .B2(new_n534), .ZN(G171));
  AOI22_X1  g110(.A1(new_n503), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n536), .A2(new_n505), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n514), .A2(G43), .ZN(new_n538));
  INV_X1    g113(.A(new_n508), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G81), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n537), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(G860), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT70), .ZN(G153));
  AND3_X1   g119(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G36), .ZN(G176));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT71), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n545), .A2(new_n549), .ZN(G188));
  INV_X1    g125(.A(G65), .ZN(new_n551));
  OAI21_X1  g126(.A(KEYINPUT72), .B1(new_n527), .B2(new_n528), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT72), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n501), .A2(new_n553), .A3(new_n502), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n551), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(G78), .A2(G543), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  OR2_X1    g132(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g133(.A(KEYINPUT73), .B1(new_n558), .B2(G651), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n507), .A2(G53), .A3(G543), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(KEYINPUT9), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT9), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n507), .A2(new_n562), .A3(G53), .A4(G543), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n561), .A2(new_n563), .B1(new_n539), .B2(G91), .ZN(new_n564));
  OAI211_X1 g139(.A(KEYINPUT73), .B(G651), .C1(new_n555), .C2(new_n557), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OR2_X1    g141(.A1(new_n559), .A2(new_n566), .ZN(G299));
  INV_X1    g142(.A(G171), .ZN(G301));
  OR2_X1    g143(.A1(new_n506), .A2(new_n512), .ZN(G303));
  NAND3_X1  g144(.A1(new_n503), .A2(new_n507), .A3(G87), .ZN(new_n570));
  INV_X1    g145(.A(G74), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n501), .A2(new_n571), .A3(new_n502), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G651), .ZN(new_n573));
  AND2_X1   g148(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n507), .A2(G49), .A3(G543), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(G288));
  NAND2_X1  g151(.A1(new_n503), .A2(G61), .ZN(new_n577));
  NAND2_X1  g152(.A1(G73), .A2(G543), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT74), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n505), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n539), .A2(G86), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n507), .A2(G48), .A3(G543), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(G305));
  AOI22_X1  g159(.A1(new_n503), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n585), .A2(new_n505), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n586), .B(KEYINPUT75), .ZN(new_n587));
  AOI22_X1  g162(.A1(G85), .A2(new_n539), .B1(new_n514), .B2(G47), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(G290));
  INV_X1    g164(.A(G66), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n590), .B1(new_n552), .B2(new_n554), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT78), .ZN(new_n593));
  NAND2_X1  g168(.A1(G79), .A2(G543), .ZN(new_n594));
  XOR2_X1   g169(.A(new_n594), .B(KEYINPUT77), .Z(new_n595));
  NAND3_X1  g170(.A1(new_n592), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n595), .ZN(new_n597));
  OAI21_X1  g172(.A(KEYINPUT78), .B1(new_n597), .B2(new_n591), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n596), .A2(G651), .A3(new_n598), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n510), .B(KEYINPUT76), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n539), .A2(KEYINPUT10), .A3(G92), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT10), .ZN(new_n602));
  INV_X1    g177(.A(G92), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n508), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n600), .A2(G54), .B1(new_n601), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n599), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(G868), .ZN(new_n607));
  MUX2_X1   g182(.A(G301), .B(new_n606), .S(new_n607), .Z(G284));
  MUX2_X1   g183(.A(G301), .B(new_n606), .S(new_n607), .Z(G321));
  MUX2_X1   g184(.A(G286), .B(G299), .S(new_n607), .Z(G297));
  MUX2_X1   g185(.A(G286), .B(G299), .S(new_n607), .Z(G280));
  AOI21_X1  g186(.A(new_n606), .B1(G559), .B2(new_n542), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT79), .ZN(G148));
  INV_X1    g188(.A(new_n606), .ZN(new_n614));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  MUX2_X1   g191(.A(new_n541), .B(new_n616), .S(G868), .Z(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g193(.A(KEYINPUT12), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n479), .A2(new_n619), .A3(G2104), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n494), .A2(new_n459), .ZN(new_n621));
  OAI21_X1  g196(.A(KEYINPUT12), .B1(new_n621), .B2(new_n463), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT13), .ZN(new_n624));
  INV_X1    g199(.A(G2100), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n479), .A2(G135), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n481), .A2(G123), .ZN(new_n629));
  AND2_X1   g204(.A1(G111), .A2(G2105), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n630), .B1(G99), .B2(new_n459), .ZN(new_n631));
  OAI211_X1 g206(.A(new_n628), .B(new_n629), .C1(new_n463), .C2(new_n631), .ZN(new_n632));
  INV_X1    g207(.A(G2096), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n626), .A2(new_n627), .A3(new_n634), .ZN(G156));
  XOR2_X1   g210(.A(G2443), .B(G2446), .Z(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT15), .B(G2435), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT81), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2427), .B(G2430), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(KEYINPUT80), .B(KEYINPUT14), .Z(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT82), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2451), .B(G2454), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT16), .Z(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n639), .A2(new_n640), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n644), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n647), .B1(new_n644), .B2(new_n648), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n636), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(new_n651), .ZN(new_n653));
  INV_X1    g228(.A(new_n636), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n653), .A2(new_n649), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1341), .B(G1348), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(new_n657), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n652), .A2(new_n655), .A3(new_n659), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n658), .A2(G14), .A3(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(G401));
  XOR2_X1   g237(.A(G2084), .B(G2090), .Z(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2072), .B(G2078), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n665), .A2(KEYINPUT17), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n663), .A2(new_n668), .ZN(new_n670));
  AND2_X1   g245(.A1(new_n670), .A2(KEYINPUT17), .ZN(new_n671));
  OAI221_X1 g246(.A(new_n669), .B1(new_n664), .B2(new_n666), .C1(new_n671), .C2(new_n665), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n663), .A2(new_n665), .A3(new_n668), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT18), .Z(new_n674));
  NAND3_X1  g249(.A1(new_n672), .A2(KEYINPUT83), .A3(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  AOI21_X1  g251(.A(KEYINPUT83), .B1(new_n672), .B2(new_n674), .ZN(new_n677));
  OAI21_X1  g252(.A(G2096), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(new_n677), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n679), .A2(new_n633), .A3(new_n675), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n681), .A2(new_n625), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n678), .A2(new_n680), .A3(G2100), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(G227));
  XOR2_X1   g259(.A(G1956), .B(G2474), .Z(new_n685));
  XOR2_X1   g260(.A(G1961), .B(G1966), .Z(new_n686));
  NAND2_X1  g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT84), .ZN(new_n688));
  XOR2_X1   g263(.A(G1971), .B(G1976), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT19), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT85), .B(KEYINPUT20), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  OR2_X1    g268(.A1(new_n685), .A2(new_n686), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(new_n690), .B2(new_n687), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n690), .A2(KEYINPUT86), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n693), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(KEYINPUT87), .Z(new_n700));
  NAND2_X1  g275(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n700), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n693), .A2(new_n702), .A3(new_n697), .ZN(new_n703));
  XNOR2_X1  g278(.A(G1991), .B(G1996), .ZN(new_n704));
  XNOR2_X1  g279(.A(G1981), .B(G1986), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  AND3_X1   g281(.A1(new_n701), .A2(new_n703), .A3(new_n706), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n706), .B1(new_n701), .B2(new_n703), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n707), .A2(new_n708), .ZN(G229));
  NAND2_X1  g284(.A1(new_n481), .A2(G128), .ZN(new_n710));
  MUX2_X1   g285(.A(G104), .B(G116), .S(G2105), .Z(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G2104), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n479), .A2(G140), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n714), .A2(KEYINPUT92), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(KEYINPUT92), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n713), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G29), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT93), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n718), .A2(G26), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT28), .ZN(new_n722));
  AND3_X1   g297(.A1(new_n720), .A2(G2067), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(G2067), .B1(new_n720), .B2(new_n722), .ZN(new_n724));
  INV_X1    g299(.A(G1348), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n614), .A2(G16), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G4), .B2(G16), .ZN(new_n727));
  OAI22_X1  g302(.A1(new_n723), .A2(new_n724), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n725), .B2(new_n727), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n632), .A2(new_n718), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT98), .Z(new_n731));
  AND2_X1   g306(.A1(KEYINPUT30), .A2(G28), .ZN(new_n732));
  NOR2_X1   g307(.A1(KEYINPUT30), .A2(G28), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n718), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  XOR2_X1   g309(.A(KEYINPUT31), .B(G11), .Z(new_n735));
  INV_X1    g310(.A(new_n735), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n736), .A2(KEYINPUT97), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n736), .A2(KEYINPUT97), .ZN(new_n738));
  NAND4_X1  g313(.A1(new_n731), .A2(new_n734), .A3(new_n737), .A4(new_n738), .ZN(new_n739));
  AND2_X1   g314(.A1(new_n739), .A2(KEYINPUT99), .ZN(new_n740));
  NOR2_X1   g315(.A1(G29), .A2(G35), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G162), .B2(G29), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT29), .ZN(new_n743));
  OAI22_X1  g318(.A1(new_n739), .A2(KEYINPUT99), .B1(G2090), .B2(new_n743), .ZN(new_n744));
  XOR2_X1   g319(.A(KEYINPUT89), .B(G16), .Z(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n746), .A2(G19), .ZN(new_n747));
  INV_X1    g322(.A(new_n541), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n747), .B1(new_n748), .B2(new_n746), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(G1341), .Z(new_n750));
  NAND2_X1  g325(.A1(G164), .A2(G29), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G27), .B2(G29), .ZN(new_n752));
  INV_X1    g327(.A(G2078), .ZN(new_n753));
  OR2_X1    g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n752), .A2(new_n753), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n750), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n743), .A2(G2090), .ZN(new_n757));
  NOR4_X1   g332(.A1(new_n740), .A2(new_n744), .A3(new_n756), .A4(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n745), .A2(G20), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT100), .Z(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT23), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G299), .B2(G16), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G1956), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n464), .A2(G103), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT94), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT25), .ZN(new_n766));
  NAND2_X1  g341(.A1(G115), .A2(G2104), .ZN(new_n767));
  INV_X1    g342(.A(G127), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n767), .B1(new_n478), .B2(new_n768), .ZN(new_n769));
  AOI22_X1  g344(.A1(new_n769), .A2(G2105), .B1(new_n479), .B2(G139), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n766), .A2(new_n770), .ZN(new_n771));
  MUX2_X1   g346(.A(G33), .B(new_n771), .S(G29), .Z(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G2072), .ZN(new_n773));
  NOR2_X1   g348(.A1(G29), .A2(G32), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n464), .A2(G105), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n479), .A2(G141), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n481), .A2(G129), .ZN(new_n777));
  NAND3_X1  g352(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT26), .Z(new_n779));
  AND4_X1   g354(.A1(new_n775), .A2(new_n776), .A3(new_n777), .A4(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n774), .B1(new_n780), .B2(G29), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT95), .ZN(new_n782));
  XOR2_X1   g357(.A(KEYINPUT27), .B(G1996), .Z(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  XOR2_X1   g359(.A(KEYINPUT24), .B(G34), .Z(new_n785));
  NOR2_X1   g360(.A1(new_n785), .A2(G29), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G160), .B2(G29), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n787), .A2(G2084), .ZN(new_n788));
  INV_X1    g363(.A(G16), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n789), .A2(G5), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G171), .B2(new_n789), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n791), .A2(G1961), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(G1961), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n784), .A2(new_n788), .A3(new_n792), .A4(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(G286), .A2(new_n789), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n795), .A2(KEYINPUT96), .ZN(new_n796));
  OAI21_X1  g371(.A(KEYINPUT96), .B1(G16), .B2(G21), .ZN(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n796), .B1(new_n795), .B2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(G1966), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  OAI22_X1  g376(.A1(new_n782), .A2(new_n783), .B1(G2084), .B2(new_n787), .ZN(new_n802));
  NOR4_X1   g377(.A1(new_n773), .A2(new_n794), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n729), .A2(new_n758), .A3(new_n763), .A4(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT90), .ZN(new_n805));
  XNOR2_X1  g380(.A(G290), .B(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n806), .A2(new_n746), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n745), .A2(G24), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(G1986), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n789), .A2(G23), .ZN(new_n812));
  INV_X1    g387(.A(G288), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n812), .B1(new_n813), .B2(new_n789), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT33), .B(G1976), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n746), .A2(G22), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(G166), .B2(new_n746), .ZN(new_n818));
  INV_X1    g393(.A(G1971), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n816), .A2(new_n820), .ZN(new_n821));
  OR2_X1    g396(.A1(G6), .A2(G16), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(G305), .B2(new_n789), .ZN(new_n823));
  XOR2_X1   g398(.A(KEYINPUT32), .B(G1981), .Z(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n821), .A2(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT34), .ZN(new_n827));
  OAI21_X1  g402(.A(KEYINPUT91), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT91), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n829), .B(KEYINPUT34), .C1(new_n821), .C2(new_n825), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n479), .A2(G131), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n481), .A2(G119), .ZN(new_n833));
  AND2_X1   g408(.A1(G107), .A2(G2105), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(G95), .B2(new_n459), .ZN(new_n835));
  OAI211_X1 g410(.A(new_n832), .B(new_n833), .C1(new_n463), .C2(new_n835), .ZN(new_n836));
  MUX2_X1   g411(.A(G25), .B(new_n836), .S(G29), .Z(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT88), .ZN(new_n838));
  XOR2_X1   g413(.A(KEYINPUT35), .B(G1991), .Z(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n838), .B(new_n840), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n841), .B1(new_n827), .B2(new_n826), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n811), .A2(new_n831), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n843), .A2(KEYINPUT36), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT36), .ZN(new_n845));
  NAND4_X1  g420(.A1(new_n811), .A2(new_n831), .A3(new_n845), .A4(new_n842), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n804), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT101), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(G311));
  INV_X1    g424(.A(new_n847), .ZN(G150));
  AOI22_X1  g425(.A1(new_n503), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n851), .A2(new_n505), .ZN(new_n852));
  INV_X1    g427(.A(G93), .ZN(new_n853));
  INV_X1    g428(.A(G55), .ZN(new_n854));
  OAI22_X1  g429(.A1(new_n508), .A2(new_n853), .B1(new_n510), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT102), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  OAI21_X1  g433(.A(KEYINPUT102), .B1(new_n852), .B2(new_n855), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(G860), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n861), .B(KEYINPUT37), .Z(new_n862));
  INV_X1    g437(.A(KEYINPUT103), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n863), .B1(new_n541), .B2(new_n856), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n864), .B1(new_n860), .B2(new_n748), .ZN(new_n865));
  NAND4_X1  g440(.A1(new_n858), .A2(new_n863), .A3(new_n541), .A4(new_n859), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT38), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n614), .A2(G559), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n868), .B(new_n869), .ZN(new_n870));
  OR2_X1    g445(.A1(new_n870), .A2(KEYINPUT39), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT104), .ZN(new_n872));
  AND2_X1   g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(G860), .B1(new_n870), .B2(KEYINPUT39), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n874), .B1(new_n871), .B2(new_n872), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n862), .B1(new_n873), .B2(new_n875), .ZN(G145));
  XNOR2_X1  g451(.A(G162), .B(new_n632), .ZN(new_n877));
  XNOR2_X1  g452(.A(G160), .B(KEYINPUT105), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n877), .B(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n481), .A2(G130), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT106), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n881), .B(new_n882), .ZN(new_n883));
  MUX2_X1   g458(.A(G106), .B(G118), .S(G2105), .Z(new_n884));
  AOI22_X1  g459(.A1(new_n479), .A2(G142), .B1(G2104), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n836), .B(new_n623), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  OR2_X1    g464(.A1(new_n836), .A2(new_n623), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n836), .A2(new_n623), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n886), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  OR2_X1    g467(.A1(new_n717), .A2(G164), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n717), .A2(G164), .ZN(new_n894));
  AND4_X1   g469(.A1(new_n889), .A2(new_n892), .A3(new_n893), .A4(new_n894), .ZN(new_n895));
  AOI22_X1  g470(.A1(new_n889), .A2(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n771), .B(new_n780), .ZN(new_n897));
  NOR3_X1   g472(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  XOR2_X1   g473(.A(new_n771), .B(new_n780), .Z(new_n899));
  NAND2_X1  g474(.A1(new_n889), .A2(new_n892), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n893), .A2(new_n894), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n889), .A2(new_n892), .A3(new_n893), .A4(new_n894), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n899), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n880), .B1(new_n898), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n897), .B1(new_n895), .B2(new_n896), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n902), .A2(new_n899), .A3(new_n903), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n906), .A2(new_n907), .A3(new_n879), .ZN(new_n908));
  XOR2_X1   g483(.A(KEYINPUT107), .B(G37), .Z(new_n909));
  NAND3_X1  g484(.A1(new_n905), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g486(.A1(new_n860), .A2(G868), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT108), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n616), .B(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(new_n867), .ZN(new_n915));
  OR2_X1    g490(.A1(G299), .A2(new_n606), .ZN(new_n916));
  NAND2_X1  g491(.A1(G299), .A2(new_n606), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT41), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n916), .A2(KEYINPUT41), .A3(new_n917), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n915), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n867), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n914), .B(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n918), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(G290), .B(G288), .ZN(new_n927));
  XNOR2_X1  g502(.A(G303), .B(G305), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n927), .B(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n929), .B1(KEYINPUT109), .B2(KEYINPUT42), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n922), .A2(new_n926), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n930), .B1(new_n922), .B2(new_n926), .ZN(new_n932));
  OAI22_X1  g507(.A1(new_n931), .A2(new_n932), .B1(KEYINPUT109), .B2(KEYINPUT42), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n922), .A2(new_n926), .ZN(new_n934));
  INV_X1    g509(.A(new_n930), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g511(.A1(KEYINPUT109), .A2(KEYINPUT42), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n922), .A2(new_n926), .A3(new_n930), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n933), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n912), .B1(new_n940), .B2(G868), .ZN(G295));
  AOI21_X1  g516(.A(new_n912), .B1(new_n940), .B2(G868), .ZN(G331));
  OR3_X1    g517(.A1(G171), .A2(KEYINPUT110), .A3(G286), .ZN(new_n943));
  OAI21_X1  g518(.A(KEYINPUT110), .B1(G171), .B2(G286), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(KEYINPUT111), .B1(G301), .B2(G168), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT111), .ZN(new_n947));
  NAND3_X1  g522(.A1(G171), .A2(new_n947), .A3(G286), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n945), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n949), .A2(new_n867), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n946), .A2(new_n948), .ZN(new_n951));
  AOI22_X1  g526(.A1(new_n951), .A2(new_n945), .B1(new_n865), .B2(new_n866), .ZN(new_n952));
  OAI211_X1 g527(.A(new_n920), .B(new_n921), .C1(new_n950), .C2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n923), .A2(new_n945), .A3(new_n951), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n949), .A2(new_n867), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n954), .A2(new_n925), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n929), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n953), .A2(new_n929), .A3(new_n956), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n959), .A2(new_n909), .A3(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT43), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(G37), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n959), .A2(KEYINPUT43), .A3(new_n964), .A4(new_n960), .ZN(new_n965));
  AOI21_X1  g540(.A(KEYINPUT44), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n959), .A2(new_n962), .A3(new_n964), .A4(new_n960), .ZN(new_n967));
  AND3_X1   g542(.A1(new_n953), .A2(new_n929), .A3(new_n956), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n929), .B1(new_n953), .B2(new_n956), .ZN(new_n969));
  INV_X1    g544(.A(new_n909), .ZN(new_n970));
  NOR3_X1   g545(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n967), .B1(new_n971), .B2(new_n962), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n966), .B1(KEYINPUT44), .B2(new_n972), .ZN(G397));
  XNOR2_X1  g548(.A(G290), .B(new_n810), .ZN(new_n974));
  INV_X1    g549(.A(G1384), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n497), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT45), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n475), .A2(new_n470), .ZN(new_n979));
  AOI21_X1  g554(.A(KEYINPUT66), .B1(new_n494), .B2(G125), .ZN(new_n980));
  OAI21_X1  g555(.A(G2105), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(new_n466), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n981), .A2(G40), .A3(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n978), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n974), .A2(new_n985), .ZN(new_n986));
  XOR2_X1   g561(.A(new_n986), .B(KEYINPUT112), .Z(new_n987));
  INV_X1    g562(.A(G1996), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n780), .B(new_n988), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n717), .B(G2067), .ZN(new_n990));
  OR2_X1    g565(.A1(new_n990), .A2(KEYINPUT113), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(KEYINPUT113), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n989), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n836), .B(new_n839), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n985), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n987), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G8), .ZN(new_n997));
  INV_X1    g572(.A(G40), .ZN(new_n998));
  AOI211_X1 g573(.A(new_n998), .B(new_n466), .C1(new_n476), .C2(G2105), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n497), .A2(KEYINPUT45), .A3(new_n975), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n978), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n800), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT50), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1003), .B1(new_n497), .B2(new_n975), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1004), .A2(new_n983), .ZN(new_n1005));
  INV_X1    g580(.A(G2084), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n497), .A2(new_n1003), .A3(new_n975), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1002), .A2(new_n1008), .A3(G168), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT124), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1010), .A2(KEYINPUT51), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(G168), .B1(new_n1002), .B2(new_n1008), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n997), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT51), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1010), .A2(new_n997), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1016), .B1(new_n1009), .B2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT62), .B1(new_n1015), .B2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT55), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1021), .B1(G166), .B2(new_n997), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n976), .A2(KEYINPUT50), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1024), .A2(new_n999), .A3(new_n1007), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1025), .A2(G2090), .ZN(new_n1026));
  AOI21_X1  g601(.A(KEYINPUT45), .B1(new_n497), .B2(new_n975), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1027), .A2(new_n983), .ZN(new_n1028));
  AOI21_X1  g603(.A(G1971), .B1(new_n1028), .B2(new_n1000), .ZN(new_n1029));
  OAI211_X1 g604(.A(G8), .B(new_n1023), .C1(new_n1026), .C2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G2090), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT118), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1007), .A2(new_n1032), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n497), .A2(KEYINPUT118), .A3(new_n1003), .A4(new_n975), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1005), .A2(new_n1031), .A3(new_n1033), .A4(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1001), .A2(new_n819), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n997), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1030), .B1(new_n1037), .B2(new_n1023), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n570), .A2(new_n573), .A3(new_n575), .A4(G1976), .ZN(new_n1039));
  XNOR2_X1  g614(.A(new_n1039), .B(KEYINPUT114), .ZN(new_n1040));
  NAND4_X1  g615(.A1(G160), .A2(G40), .A3(new_n975), .A4(new_n497), .ZN(new_n1041));
  XNOR2_X1  g616(.A(KEYINPUT115), .B(G1976), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1042), .B1(new_n574), .B2(new_n575), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1040), .A2(new_n1041), .A3(G8), .A4(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1040), .A2(new_n1041), .A3(KEYINPUT116), .A4(G8), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n1040), .A2(new_n1041), .A3(G8), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1049), .A2(new_n1044), .A3(KEYINPUT116), .A4(new_n1045), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1041), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1051), .A2(new_n997), .ZN(new_n1052));
  INV_X1    g627(.A(G1981), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n581), .A2(new_n582), .A3(new_n1053), .A4(new_n583), .ZN(new_n1054));
  XOR2_X1   g629(.A(KEYINPUT117), .B(G86), .Z(new_n1055));
  OAI21_X1  g630(.A(new_n583), .B1(new_n508), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(G1981), .B1(new_n1056), .B2(new_n580), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1054), .A2(KEYINPUT49), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1054), .A2(new_n1057), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT49), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1052), .A2(new_n1058), .A3(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1048), .A2(new_n1050), .A3(new_n1062), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n978), .A2(new_n999), .A3(new_n753), .A4(new_n1000), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT53), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1028), .A2(KEYINPUT53), .A3(new_n753), .A4(new_n1000), .ZN(new_n1067));
  INV_X1    g642(.A(G1961), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1025), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1066), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(G171), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n1038), .A2(new_n1063), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT62), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1009), .A2(new_n1017), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT51), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1013), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1073), .B(new_n1075), .C1(new_n1076), .C2(new_n997), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1019), .A2(new_n1072), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(G1976), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1062), .A2(new_n1079), .A3(new_n813), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(new_n1054), .ZN(new_n1081));
  AND3_X1   g656(.A1(new_n1048), .A2(new_n1050), .A3(new_n1062), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1030), .ZN(new_n1083));
  AOI22_X1  g658(.A1(new_n1052), .A2(new_n1081), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1033), .A2(new_n1024), .A3(new_n999), .A4(new_n1034), .ZN(new_n1085));
  INV_X1    g660(.A(G1956), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  XNOR2_X1  g662(.A(KEYINPUT56), .B(G2072), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1028), .A2(new_n1000), .A3(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT120), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1091), .B1(new_n559), .B2(new_n566), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT57), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1091), .B(KEYINPUT57), .C1(new_n559), .C2(new_n566), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1090), .A2(new_n1096), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1087), .A2(new_n1094), .A3(new_n1095), .A4(new_n1089), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(G1348), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1041), .A2(G2067), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n614), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1097), .B1(new_n1099), .B2(new_n1102), .ZN(new_n1103));
  AOI22_X1  g678(.A1(new_n1087), .A2(new_n1089), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1104));
  OAI21_X1  g679(.A(KEYINPUT61), .B1(new_n1099), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT61), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1097), .A2(new_n1106), .A3(new_n1098), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  XOR2_X1   g683(.A(KEYINPUT121), .B(G1996), .Z(new_n1109));
  NAND4_X1  g684(.A1(new_n978), .A2(new_n999), .A3(new_n1000), .A4(new_n1109), .ZN(new_n1110));
  XOR2_X1   g685(.A(KEYINPUT58), .B(G1341), .Z(new_n1111));
  OAI21_X1  g686(.A(new_n1111), .B1(new_n983), .B2(new_n976), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n541), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT122), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT123), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n1114), .A2(new_n1115), .A3(KEYINPUT59), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1113), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1025), .A2(new_n725), .ZN(new_n1118));
  INV_X1    g693(.A(G2067), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1051), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT60), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1118), .A2(new_n1120), .A3(new_n1121), .A4(new_n614), .ZN(new_n1122));
  OAI211_X1 g697(.A(new_n1117), .B(new_n1122), .C1(new_n1114), .C2(new_n1113), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1118), .A2(new_n1120), .A3(new_n606), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1121), .B1(new_n1102), .B2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(KEYINPUT59), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1126));
  NOR3_X1   g701(.A1(new_n1123), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1103), .B1(new_n1108), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT125), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n497), .A2(new_n1003), .A3(new_n975), .ZN(new_n1130));
  NOR3_X1   g705(.A1(new_n1130), .A2(new_n1004), .A3(new_n983), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1129), .B1(new_n1131), .B2(G1961), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1025), .A2(KEYINPUT125), .A3(new_n1068), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1132), .A2(new_n1066), .A3(new_n1067), .A4(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1071), .B1(new_n1134), .B2(G171), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT54), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1075), .B1(new_n1076), .B2(new_n997), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1038), .A2(new_n1063), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1134), .A2(G171), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1066), .A2(new_n1067), .A3(new_n1069), .A4(G301), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1140), .A2(KEYINPUT54), .A3(new_n1141), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1137), .A2(new_n1138), .A3(new_n1139), .A4(new_n1142), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1078), .B(new_n1084), .C1(new_n1128), .C2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT119), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1002), .A2(new_n1008), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1146), .A2(G8), .A3(G168), .ZN(new_n1147));
  NOR3_X1   g722(.A1(new_n1038), .A2(new_n1063), .A3(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1145), .B1(new_n1148), .B2(KEYINPUT63), .ZN(new_n1149));
  OR2_X1    g724(.A1(new_n1037), .A2(new_n1023), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1147), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1082), .A2(new_n1150), .A3(new_n1030), .A4(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT63), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1152), .A2(KEYINPUT119), .A3(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1151), .A2(KEYINPUT63), .A3(new_n1030), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1023), .ZN(new_n1156));
  OAI21_X1  g731(.A(G8), .B1(new_n1026), .B2(new_n1029), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1155), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  AOI22_X1  g733(.A1(new_n1149), .A2(new_n1154), .B1(new_n1158), .B2(new_n1082), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n996), .B1(new_n1144), .B2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n836), .A2(new_n840), .ZN(new_n1161));
  AOI22_X1  g736(.A1(new_n993), .A2(new_n1161), .B1(new_n1119), .B2(new_n717), .ZN(new_n1162));
  NOR3_X1   g737(.A1(new_n985), .A2(G1986), .A3(G290), .ZN(new_n1163));
  XNOR2_X1  g738(.A(new_n1163), .B(KEYINPUT48), .ZN(new_n1164));
  OAI22_X1  g739(.A1(new_n1162), .A2(new_n985), .B1(new_n995), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n991), .A2(new_n992), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n985), .B1(new_n1166), .B2(new_n780), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n984), .A2(new_n988), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n1168), .B(KEYINPUT46), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1169), .ZN(new_n1170));
  OAI21_X1  g745(.A(KEYINPUT47), .B1(new_n1167), .B2(new_n1170), .ZN(new_n1171));
  OR3_X1    g746(.A1(new_n1167), .A2(KEYINPUT47), .A3(new_n1170), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1165), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1160), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1174), .A2(KEYINPUT126), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT126), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1160), .A2(new_n1176), .A3(new_n1173), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1175), .A2(new_n1177), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g753(.A(G319), .B1(new_n707), .B2(new_n708), .ZN(new_n1180));
  NOR2_X1   g754(.A1(new_n1180), .A2(G227), .ZN(new_n1181));
  AND3_X1   g755(.A1(new_n1181), .A2(new_n910), .A3(new_n661), .ZN(new_n1182));
  OAI211_X1 g756(.A(new_n1182), .B(new_n965), .C1(new_n971), .C2(KEYINPUT43), .ZN(new_n1183));
  XNOR2_X1  g757(.A(new_n1183), .B(KEYINPUT127), .ZN(G308));
  INV_X1    g758(.A(KEYINPUT127), .ZN(new_n1185));
  XNOR2_X1  g759(.A(new_n1183), .B(new_n1185), .ZN(G225));
endmodule


