//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 1 1 0 1 0 0 1 1 0 0 1 0 0 1 0 0 0 1 1 0 1 0 0 0 0 0 1 0 1 1 1 1 0 1 0 1 0 1 0 0 0 1 0 1 0 0 1 0 0 1 0 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n791, new_n792,
    new_n793, new_n794, new_n796, new_n797, new_n798, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n849, new_n850, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n864, new_n865, new_n867, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913;
  XOR2_X1   g000(.A(KEYINPUT70), .B(KEYINPUT36), .Z(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g002(.A1(G227gat), .A2(G233gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT23), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT64), .ZN(new_n209));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210));
  AOI22_X1  g009(.A1(new_n207), .A2(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G183gat), .ZN(new_n212));
  INV_X1    g011(.A(G190gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(G183gat), .A2(G190gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n214), .A2(KEYINPUT24), .A3(new_n215), .ZN(new_n216));
  OR2_X1    g015(.A1(new_n215), .A2(KEYINPUT24), .ZN(new_n217));
  NAND3_X1  g016(.A1(KEYINPUT64), .A2(G169gat), .A3(G176gat), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n211), .A2(new_n216), .A3(new_n217), .A4(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(KEYINPUT25), .ZN(new_n220));
  XNOR2_X1  g019(.A(KEYINPUT27), .B(G183gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(new_n213), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n222), .A2(KEYINPUT65), .A3(KEYINPUT28), .ZN(new_n223));
  XOR2_X1   g022(.A(KEYINPUT65), .B(KEYINPUT28), .Z(new_n224));
  NAND3_X1  g023(.A1(new_n224), .A2(new_n213), .A3(new_n221), .ZN(new_n225));
  AND2_X1   g024(.A1(new_n205), .A2(KEYINPUT26), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n205), .A2(KEYINPUT26), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n210), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n223), .A2(new_n225), .A3(new_n215), .A4(new_n228), .ZN(new_n229));
  AND3_X1   g028(.A1(new_n216), .A2(new_n210), .A3(new_n217), .ZN(new_n230));
  AOI21_X1  g029(.A(KEYINPUT25), .B1(new_n207), .B2(new_n208), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n220), .A2(new_n229), .A3(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(G127gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(G134gat), .ZN(new_n235));
  INV_X1    g034(.A(G134gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(G127gat), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT66), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n235), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n234), .A2(KEYINPUT66), .A3(G134gat), .ZN(new_n240));
  XNOR2_X1  g039(.A(G113gat), .B(G120gat), .ZN(new_n241));
  OAI211_X1 g040(.A(new_n239), .B(new_n240), .C1(KEYINPUT1), .C2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT67), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT1), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(G127gat), .B(G134gat), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n247), .B1(new_n241), .B2(new_n243), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n242), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n249), .ZN(new_n250));
  AOI22_X1  g049(.A1(new_n219), .A2(KEYINPUT25), .B1(new_n231), .B2(new_n230), .ZN(new_n251));
  INV_X1    g050(.A(new_n249), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n251), .A2(new_n252), .A3(new_n229), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n204), .B1(new_n250), .B2(new_n253), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n254), .A2(KEYINPUT68), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT68), .ZN(new_n256));
  AOI211_X1 g055(.A(new_n256), .B(new_n204), .C1(new_n250), .C2(new_n253), .ZN(new_n257));
  OAI21_X1  g056(.A(KEYINPUT32), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT33), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n259), .B1(new_n255), .B2(new_n257), .ZN(new_n260));
  XNOR2_X1  g059(.A(G15gat), .B(G43gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(G71gat), .B(G99gat), .ZN(new_n262));
  XOR2_X1   g061(.A(new_n261), .B(new_n262), .Z(new_n263));
  NAND3_X1  g062(.A1(new_n258), .A2(new_n260), .A3(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n263), .ZN(new_n265));
  OAI221_X1 g064(.A(KEYINPUT32), .B1(new_n259), .B2(new_n265), .C1(new_n255), .C2(new_n257), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n250), .A2(new_n204), .A3(new_n253), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n268), .B(KEYINPUT34), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n269), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n264), .A2(new_n271), .A3(new_n266), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n203), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n270), .A2(KEYINPUT69), .A3(new_n272), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT69), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n267), .A2(new_n275), .A3(new_n269), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n273), .B1(new_n277), .B2(KEYINPUT36), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT3), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT22), .ZN(new_n280));
  INV_X1    g079(.A(G211gat), .ZN(new_n281));
  INV_X1    g080(.A(G218gat), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT71), .ZN(new_n284));
  XNOR2_X1  g083(.A(G197gat), .B(G204gat), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT71), .ZN(new_n286));
  OAI211_X1 g085(.A(new_n286), .B(new_n280), .C1(new_n281), .C2(new_n282), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n284), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(G211gat), .B(G218gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n288), .B(new_n289), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n279), .B1(new_n290), .B2(KEYINPUT29), .ZN(new_n291));
  XOR2_X1   g090(.A(G141gat), .B(G148gat), .Z(new_n292));
  NAND2_X1  g091(.A1(G155gat), .A2(G162gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT2), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT77), .ZN(new_n295));
  INV_X1    g094(.A(G155gat), .ZN(new_n296));
  INV_X1    g095(.A(G162gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(new_n293), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT77), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n293), .A2(new_n300), .A3(KEYINPUT2), .ZN(new_n301));
  NAND4_X1  g100(.A1(new_n292), .A2(new_n295), .A3(new_n299), .A4(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(G141gat), .B(G148gat), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n293), .B(new_n298), .C1(new_n303), .C2(KEYINPUT2), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n291), .A2(new_n305), .ZN(new_n306));
  AND2_X1   g105(.A1(new_n302), .A2(new_n304), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(new_n279), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT29), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(new_n290), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n306), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(G50gat), .ZN(new_n313));
  INV_X1    g112(.A(G50gat), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n306), .A2(new_n314), .A3(new_n311), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(KEYINPUT31), .B(G22gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(G228gat), .A2(G233gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n317), .B(new_n318), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  XNOR2_X1  g120(.A(G78gat), .B(G106gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n316), .A2(new_n319), .ZN(new_n323));
  AND3_X1   g122(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n322), .B1(new_n321), .B2(new_n323), .ZN(new_n325));
  OR2_X1    g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(KEYINPUT0), .B(G57gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n327), .B(G85gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(G1gat), .B(G29gat), .ZN(new_n329));
  XOR2_X1   g128(.A(new_n328), .B(new_n329), .Z(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT5), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT1), .B1(new_n241), .B2(new_n243), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n333), .B(new_n247), .C1(new_n243), .C2(new_n241), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n307), .A2(KEYINPUT79), .A3(new_n242), .A4(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT79), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n336), .B1(new_n249), .B2(new_n305), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n335), .B(new_n337), .C1(new_n252), .C2(new_n307), .ZN(new_n338));
  NAND2_X1  g137(.A1(G225gat), .A2(G233gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n339), .B(KEYINPUT78), .ZN(new_n340));
  AND2_X1   g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT80), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT4), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n335), .A2(new_n337), .A3(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n252), .A2(KEYINPUT4), .A3(new_n307), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n305), .A2(KEYINPUT3), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n308), .A2(new_n249), .A3(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n340), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n342), .B1(new_n346), .B2(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n305), .B(new_n279), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n340), .B1(new_n352), .B2(new_n249), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n353), .A2(KEYINPUT80), .A3(new_n344), .A4(new_n345), .ZN(new_n354));
  AOI211_X1 g153(.A(new_n332), .B(new_n341), .C1(new_n351), .C2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n335), .A2(new_n337), .A3(KEYINPUT4), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT81), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n252), .A2(new_n343), .A3(new_n307), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT81), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n335), .A2(new_n337), .A3(new_n359), .A4(KEYINPUT4), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n357), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n350), .A2(KEYINPUT5), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n331), .B1(new_n355), .B2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT6), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n351), .A2(new_n354), .ZN(new_n367));
  INV_X1    g166(.A(new_n341), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n367), .A2(KEYINPUT5), .A3(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n369), .A2(new_n330), .A3(new_n363), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n365), .A2(new_n366), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT82), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n365), .A2(KEYINPUT82), .A3(new_n370), .A4(new_n366), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n330), .B1(new_n369), .B2(new_n363), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT6), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n373), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n233), .A2(new_n309), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT74), .ZN(new_n379));
  NAND2_X1  g178(.A1(G226gat), .A2(G233gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n380), .B(KEYINPUT72), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n378), .A2(new_n379), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(KEYINPUT29), .B1(new_n251), .B2(new_n229), .ZN(new_n383));
  INV_X1    g182(.A(new_n381), .ZN(new_n384));
  OAI21_X1  g183(.A(KEYINPUT74), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n290), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n381), .B(KEYINPUT73), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n233), .A2(new_n387), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n382), .A2(new_n385), .A3(new_n386), .A4(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(G8gat), .B(G36gat), .ZN(new_n390));
  INV_X1    g189(.A(G64gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n390), .B(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n392), .B(G92gat), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n233), .A2(new_n384), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n394), .B1(new_n383), .B2(new_n387), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(new_n290), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n389), .A2(new_n393), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(KEYINPUT76), .ZN(new_n398));
  OR2_X1    g197(.A1(new_n398), .A2(KEYINPUT30), .ZN(new_n399));
  AND2_X1   g198(.A1(new_n389), .A2(new_n396), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n393), .B(KEYINPUT75), .ZN(new_n401));
  OR2_X1    g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n398), .A2(KEYINPUT30), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n399), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n326), .B1(new_n377), .B2(new_n405), .ZN(new_n406));
  AND2_X1   g205(.A1(new_n371), .A2(new_n376), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT86), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT37), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n389), .A2(new_n409), .A3(new_n396), .ZN(new_n410));
  XOR2_X1   g209(.A(KEYINPUT84), .B(KEYINPUT38), .Z(new_n411));
  NOR2_X1   g210(.A1(new_n401), .A2(new_n411), .ZN(new_n412));
  AND2_X1   g211(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT85), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n382), .A2(new_n385), .A3(new_n290), .A4(new_n388), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n409), .B1(new_n395), .B2(new_n386), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT83), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  AND3_X1   g216(.A1(new_n415), .A2(new_n416), .A3(KEYINPUT83), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n413), .B(new_n414), .C1(new_n417), .C2(new_n418), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n410), .B(new_n412), .C1(new_n418), .C2(new_n417), .ZN(new_n420));
  AOI22_X1  g219(.A1(new_n420), .A2(KEYINPUT85), .B1(new_n393), .B2(new_n400), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n407), .A2(new_n408), .A3(new_n419), .A4(new_n421), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n421), .A2(new_n371), .A3(new_n376), .A4(new_n419), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT86), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n400), .A2(new_n409), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n425), .A2(new_n393), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(new_n410), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(new_n411), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n422), .A2(new_n424), .A3(new_n428), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n324), .A2(new_n325), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n349), .B1(new_n361), .B2(new_n348), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT39), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n331), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n338), .A2(new_n340), .ZN(new_n434));
  OR2_X1    g233(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n433), .B1(new_n435), .B2(new_n432), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT40), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n405), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n375), .B1(new_n436), .B2(new_n437), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n430), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  AOI211_X1 g240(.A(new_n278), .B(new_n406), .C1(new_n429), .C2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT35), .ZN(new_n443));
  INV_X1    g242(.A(new_n270), .ZN(new_n444));
  INV_X1    g243(.A(new_n272), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n446), .A2(new_n326), .A3(new_n405), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n443), .B1(new_n447), .B2(new_n407), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n430), .B1(new_n274), .B2(new_n276), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n449), .A2(new_n377), .A3(KEYINPUT35), .A4(new_n405), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(KEYINPUT87), .B1(new_n442), .B2(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n278), .B1(new_n429), .B2(new_n441), .ZN(new_n453));
  INV_X1    g252(.A(new_n406), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT87), .ZN(new_n456));
  INV_X1    g255(.A(new_n451), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n452), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(G127gat), .B(G155gat), .ZN(new_n460));
  XOR2_X1   g259(.A(new_n460), .B(KEYINPUT96), .Z(new_n461));
  XNOR2_X1  g260(.A(G15gat), .B(G22gat), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n462), .A2(KEYINPUT89), .A3(G1gat), .ZN(new_n463));
  INV_X1    g262(.A(new_n462), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n463), .B1(KEYINPUT16), .B2(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(G1gat), .B1(new_n462), .B2(KEYINPUT89), .ZN(new_n466));
  OR3_X1    g265(.A1(new_n465), .A2(G8gat), .A3(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(G8gat), .B1(new_n465), .B2(new_n466), .ZN(new_n468));
  AND3_X1   g267(.A1(new_n467), .A2(KEYINPUT90), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(KEYINPUT90), .B1(new_n467), .B2(new_n468), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT93), .ZN(new_n472));
  INV_X1    g271(.A(G57gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(KEYINPUT93), .A2(G57gat), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n391), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n473), .A2(G64gat), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT94), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(G71gat), .A2(G78gat), .ZN(new_n479));
  OR2_X1    g278(.A1(G71gat), .A2(G78gat), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT9), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n475), .ZN(new_n483));
  NOR2_X1   g282(.A1(KEYINPUT93), .A2(G57gat), .ZN(new_n484));
  OAI21_X1  g283(.A(G64gat), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT94), .ZN(new_n486));
  INV_X1    g285(.A(new_n477), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n478), .A2(new_n482), .A3(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(G57gat), .B(G64gat), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n480), .B(new_n479), .C1(new_n490), .C2(new_n481), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT95), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n489), .A2(KEYINPUT95), .A3(new_n491), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(KEYINPUT21), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n471), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(G183gat), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n471), .A2(new_n212), .A3(new_n497), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(G231gat), .A2(G233gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n501), .A2(new_n502), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n461), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n505), .ZN(new_n507));
  INV_X1    g306(.A(new_n461), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n507), .A2(new_n503), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  OR2_X1    g309(.A1(new_n496), .A2(KEYINPUT21), .ZN(new_n511));
  XNOR2_X1  g310(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n512), .B(G211gat), .ZN(new_n513));
  XOR2_X1   g312(.A(new_n511), .B(new_n513), .Z(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n510), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n506), .A2(new_n509), .A3(new_n514), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(G134gat), .B(G162gat), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n519), .B(KEYINPUT97), .ZN(new_n520));
  AND2_X1   g319(.A1(G232gat), .A2(G233gat), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n521), .A2(KEYINPUT41), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n520), .B(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(G99gat), .A2(G106gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(KEYINPUT8), .ZN(new_n525));
  NAND2_X1  g324(.A1(G85gat), .A2(G92gat), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT7), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(G85gat), .ZN(new_n529));
  INV_X1    g328(.A(G92gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n525), .A2(new_n528), .A3(new_n531), .A4(new_n532), .ZN(new_n533));
  AND2_X1   g332(.A1(G99gat), .A2(G106gat), .ZN(new_n534));
  NOR2_X1   g333(.A1(G99gat), .A2(G106gat), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n533), .B(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  NOR2_X1   g337(.A1(G29gat), .A2(G36gat), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT14), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n539), .B(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(G29gat), .A2(G36gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(G43gat), .B(G50gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(KEYINPUT15), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  XOR2_X1   g346(.A(G43gat), .B(G50gat), .Z(new_n548));
  INV_X1    g347(.A(KEYINPUT15), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT88), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n542), .B(new_n551), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n550), .A2(new_n541), .A3(new_n545), .A4(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n547), .A2(new_n553), .ZN(new_n554));
  AOI22_X1  g353(.A1(new_n538), .A2(new_n554), .B1(KEYINPUT41), .B2(new_n521), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT17), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n554), .B(new_n556), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n555), .B1(new_n557), .B2(new_n538), .ZN(new_n558));
  XNOR2_X1  g357(.A(G190gat), .B(G218gat), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n523), .B1(new_n560), .B2(KEYINPUT98), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n558), .B(new_n559), .ZN(new_n562));
  AND2_X1   g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n561), .A2(new_n562), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n518), .A2(new_n566), .ZN(new_n567));
  XOR2_X1   g366(.A(new_n471), .B(new_n554), .Z(new_n568));
  NAND2_X1  g367(.A1(G229gat), .A2(G233gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(KEYINPUT92), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(KEYINPUT13), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n467), .A2(new_n468), .ZN(new_n573));
  OR2_X1    g372(.A1(new_n557), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n554), .B1(new_n469), .B2(new_n470), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n574), .A2(new_n575), .A3(new_n569), .ZN(new_n576));
  NOR2_X1   g375(.A1(KEYINPUT91), .A2(KEYINPUT18), .ZN(new_n577));
  OR2_X1    g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n577), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n572), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(KEYINPUT11), .B(G169gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(G197gat), .ZN(new_n582));
  XOR2_X1   g381(.A(G113gat), .B(G141gat), .Z(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(KEYINPUT12), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n580), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n572), .A2(new_n585), .A3(new_n578), .A4(new_n579), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(G230gat), .A2(G233gat), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n494), .A2(new_n537), .A3(new_n495), .ZN(new_n592));
  INV_X1    g391(.A(new_n535), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n593), .A2(KEYINPUT99), .A3(new_n524), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n533), .A2(new_n594), .ZN(new_n595));
  AND3_X1   g394(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n596));
  AOI21_X1  g395(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AOI22_X1  g397(.A1(KEYINPUT8), .A2(new_n524), .B1(new_n529), .B2(new_n530), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n598), .A2(new_n599), .A3(new_n536), .A4(KEYINPUT99), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n595), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n489), .A2(new_n491), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(KEYINPUT100), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT100), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n489), .A2(new_n604), .A3(new_n601), .A4(new_n491), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT10), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n592), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n496), .A2(KEYINPUT10), .A3(new_n538), .ZN(new_n609));
  AND3_X1   g408(.A1(new_n608), .A2(KEYINPUT101), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(KEYINPUT101), .B1(new_n608), .B2(new_n609), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n591), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  XOR2_X1   g411(.A(G120gat), .B(G148gat), .Z(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(G176gat), .ZN(new_n614));
  INV_X1    g413(.A(G204gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  AND2_X1   g416(.A1(new_n592), .A2(new_n606), .ZN(new_n618));
  OAI211_X1 g417(.A(new_n612), .B(new_n617), .C1(new_n591), .C2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n591), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n620), .B1(new_n608), .B2(new_n609), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n618), .A2(new_n591), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n616), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n619), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n590), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n459), .A2(new_n567), .A3(new_n625), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n626), .A2(new_n377), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n627), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g427(.A1(new_n626), .A2(new_n405), .ZN(new_n629));
  NAND2_X1  g428(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n630));
  OR2_X1    g429(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT42), .ZN(new_n633));
  OR2_X1    g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  INV_X1    g434(.A(G8gat), .ZN(new_n636));
  OAI211_X1 g435(.A(new_n634), .B(new_n635), .C1(new_n636), .C2(new_n629), .ZN(G1325gat));
  INV_X1    g436(.A(G15gat), .ZN(new_n638));
  INV_X1    g437(.A(new_n278), .ZN(new_n639));
  NOR3_X1   g438(.A1(new_n626), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n446), .ZN(new_n641));
  OR2_X1    g440(.A1(new_n626), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n640), .B1(new_n638), .B2(new_n642), .ZN(G1326gat));
  NOR2_X1   g442(.A1(new_n626), .A2(new_n326), .ZN(new_n644));
  XOR2_X1   g443(.A(KEYINPUT43), .B(G22gat), .Z(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(G1327gat));
  AOI21_X1  g445(.A(new_n565), .B1(new_n452), .B2(new_n458), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n647), .A2(new_n518), .A3(new_n625), .ZN(new_n648));
  NOR3_X1   g447(.A1(new_n648), .A2(G29gat), .A3(new_n377), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n649), .B(KEYINPUT45), .Z(new_n650));
  AOI21_X1  g449(.A(new_n451), .B1(new_n453), .B2(new_n454), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT44), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n652), .A2(new_n653), .A3(new_n566), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n654), .B1(new_n647), .B2(new_n653), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n625), .A2(new_n518), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(KEYINPUT102), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(G29gat), .B1(new_n659), .B2(new_n377), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n650), .A2(new_n660), .ZN(G1328gat));
  OR3_X1    g460(.A1(new_n648), .A2(G36gat), .A3(new_n405), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT46), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n663), .A2(KEYINPUT103), .ZN(new_n664));
  AND2_X1   g463(.A1(new_n663), .A2(KEYINPUT103), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n662), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(G36gat), .B1(new_n659), .B2(new_n405), .ZN(new_n667));
  OAI211_X1 g466(.A(new_n666), .B(new_n667), .C1(new_n664), .C2(new_n662), .ZN(G1329gat));
  NAND4_X1  g467(.A1(new_n655), .A2(G43gat), .A3(new_n278), .A4(new_n658), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT104), .ZN(new_n670));
  INV_X1    g469(.A(G43gat), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n671), .B1(new_n648), .B2(new_n641), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n669), .A2(new_n670), .A3(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n670), .B1(new_n669), .B2(new_n672), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT47), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n669), .A2(new_n672), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(KEYINPUT104), .ZN(new_n679));
  AOI21_X1  g478(.A(KEYINPUT47), .B1(new_n679), .B2(new_n673), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n677), .A2(new_n680), .ZN(G1330gat));
  OAI21_X1  g480(.A(G50gat), .B1(new_n659), .B2(new_n326), .ZN(new_n682));
  OR3_X1    g481(.A1(new_n648), .A2(G50gat), .A3(new_n326), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g483(.A(KEYINPUT48), .B1(new_n683), .B2(KEYINPUT105), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1331gat));
  INV_X1    g485(.A(new_n624), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n516), .A2(new_n590), .A3(new_n565), .A4(new_n517), .ZN(new_n688));
  OR3_X1    g487(.A1(new_n651), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n689), .A2(new_n377), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n474), .A2(new_n475), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(G1332gat));
  AOI21_X1  g491(.A(new_n689), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(new_n404), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT106), .ZN(new_n695));
  OR2_X1    g494(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(G1333gat));
  INV_X1    g496(.A(G71gat), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n689), .A2(new_n698), .A3(new_n639), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT107), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n698), .B1(new_n689), .B2(new_n641), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g502(.A1(new_n689), .A2(new_n326), .ZN(new_n704));
  XOR2_X1   g503(.A(KEYINPUT108), .B(G78gat), .Z(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT109), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n704), .B(new_n706), .ZN(G1335gat));
  NAND2_X1  g506(.A1(new_n518), .A2(new_n590), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n708), .A2(new_n687), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT110), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n655), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(G85gat), .B1(new_n711), .B2(new_n377), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT111), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n713), .B1(new_n651), .B2(new_n565), .ZN(new_n714));
  INV_X1    g513(.A(new_n708), .ZN(new_n715));
  OAI211_X1 g514(.A(KEYINPUT111), .B(new_n566), .C1(new_n442), .C2(new_n451), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  OR2_X1    g517(.A1(new_n718), .A2(KEYINPUT51), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(KEYINPUT51), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(new_n624), .ZN(new_n722));
  INV_X1    g521(.A(new_n377), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(new_n529), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n712), .B1(new_n722), .B2(new_n724), .ZN(G1336gat));
  XOR2_X1   g524(.A(KEYINPUT112), .B(KEYINPUT51), .Z(new_n726));
  NAND2_X1  g525(.A1(new_n717), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(KEYINPUT113), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT113), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n717), .A2(new_n729), .A3(new_n726), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n728), .A2(new_n720), .A3(new_n730), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n405), .A2(G92gat), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n731), .A2(new_n624), .A3(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(G92gat), .B1(new_n711), .B2(new_n405), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(KEYINPUT52), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n721), .A2(new_n624), .A3(new_n732), .ZN(new_n737));
  XNOR2_X1  g536(.A(KEYINPUT114), .B(KEYINPUT52), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n737), .A2(new_n734), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n736), .A2(new_n739), .ZN(G1337gat));
  OAI21_X1  g539(.A(G99gat), .B1(new_n711), .B2(new_n639), .ZN(new_n741));
  INV_X1    g540(.A(G99gat), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n721), .A2(new_n742), .A3(new_n624), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n741), .B1(new_n743), .B2(new_n641), .ZN(G1338gat));
  NOR3_X1   g543(.A1(new_n326), .A2(G106gat), .A3(new_n687), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n721), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n655), .A2(new_n430), .A3(new_n710), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(G106gat), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT53), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n746), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  AOI22_X1  g549(.A1(new_n731), .A2(new_n745), .B1(new_n747), .B2(G106gat), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n750), .B1(new_n751), .B2(new_n749), .ZN(G1339gat));
  INV_X1    g551(.A(KEYINPUT54), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n617), .B1(new_n621), .B2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT115), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n608), .A2(new_n620), .A3(new_n609), .ZN(new_n756));
  AND2_X1   g555(.A1(new_n756), .A2(KEYINPUT54), .ZN(new_n757));
  AND3_X1   g556(.A1(new_n612), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n755), .B1(new_n612), .B2(new_n757), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n754), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT55), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  OAI211_X1 g561(.A(KEYINPUT55), .B(new_n754), .C1(new_n758), .C2(new_n759), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n762), .A2(new_n589), .A3(new_n619), .A4(new_n763), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n568), .A2(new_n571), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n569), .B1(new_n574), .B2(new_n575), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n584), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n624), .A2(new_n588), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n764), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n565), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT116), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n767), .B(new_n588), .C1(new_n564), .C2(new_n563), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n773), .A2(new_n619), .A3(new_n762), .A4(new_n763), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n770), .A2(new_n771), .A3(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n566), .B1(new_n764), .B2(new_n768), .ZN(new_n776));
  INV_X1    g575(.A(new_n774), .ZN(new_n777));
  OAI21_X1  g576(.A(KEYINPUT116), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n775), .A2(new_n518), .A3(new_n778), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n688), .A2(new_n624), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n377), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  AND2_X1   g581(.A1(new_n782), .A2(new_n449), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n783), .A2(new_n405), .ZN(new_n784));
  INV_X1    g583(.A(G113gat), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n784), .A2(new_n785), .A3(new_n589), .ZN(new_n786));
  INV_X1    g585(.A(new_n447), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n782), .A2(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(G113gat), .B1(new_n788), .B2(new_n590), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n786), .A2(new_n789), .ZN(G1340gat));
  INV_X1    g589(.A(G120gat), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n784), .A2(new_n791), .A3(new_n624), .ZN(new_n792));
  OAI21_X1  g591(.A(G120gat), .B1(new_n788), .B2(new_n687), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  XOR2_X1   g593(.A(new_n794), .B(KEYINPUT117), .Z(G1341gat));
  NOR3_X1   g594(.A1(new_n788), .A2(new_n234), .A3(new_n518), .ZN(new_n796));
  INV_X1    g595(.A(new_n518), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n784), .A2(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n796), .B1(new_n798), .B2(new_n234), .ZN(G1342gat));
  NOR2_X1   g598(.A1(new_n404), .A2(new_n565), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n783), .A2(new_n236), .A3(new_n800), .ZN(new_n801));
  XOR2_X1   g600(.A(new_n801), .B(KEYINPUT56), .Z(new_n802));
  OAI21_X1  g601(.A(G134gat), .B1(new_n788), .B2(new_n565), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n803), .B(KEYINPUT118), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(G1343gat));
  NAND2_X1  g604(.A1(new_n779), .A2(new_n781), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n430), .ZN(new_n807));
  XOR2_X1   g606(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n807), .A2(KEYINPUT120), .A3(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n518), .B1(new_n776), .B2(new_n777), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n326), .B1(new_n811), .B2(new_n781), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(KEYINPUT57), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT120), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n326), .B1(new_n779), .B2(new_n781), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n814), .B1(new_n815), .B2(new_n808), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n810), .A2(new_n813), .A3(new_n816), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n278), .A2(new_n377), .A3(new_n404), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(G141gat), .B1(new_n819), .B2(new_n590), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT121), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n278), .A2(new_n326), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n782), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n823), .A2(new_n404), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n590), .A2(G141gat), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n821), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n820), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(KEYINPUT58), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT58), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n820), .A2(new_n829), .A3(new_n826), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n828), .A2(new_n830), .ZN(G1344gat));
  INV_X1    g630(.A(KEYINPUT59), .ZN(new_n832));
  OAI211_X1 g631(.A(new_n832), .B(G148gat), .C1(new_n819), .C2(new_n687), .ZN(new_n833));
  INV_X1    g632(.A(G148gat), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n806), .A2(new_n430), .A3(new_n808), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT122), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n797), .B1(new_n770), .B2(new_n774), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n430), .B1(new_n837), .B2(new_n780), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT57), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n836), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n812), .A2(KEYINPUT122), .A3(KEYINPUT57), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n835), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n843), .A2(new_n687), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n834), .B1(new_n844), .B2(new_n818), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n833), .B1(new_n845), .B2(new_n832), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n824), .A2(new_n834), .A3(new_n624), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(G1345gat));
  AOI21_X1  g647(.A(G155gat), .B1(new_n824), .B2(new_n797), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n819), .A2(new_n296), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n849), .B1(new_n850), .B2(new_n797), .ZN(G1346gat));
  OAI21_X1  g650(.A(G162gat), .B1(new_n819), .B2(new_n565), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n800), .A2(new_n297), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n852), .B1(new_n823), .B2(new_n853), .ZN(G1347gat));
  AOI21_X1  g653(.A(new_n723), .B1(new_n779), .B2(new_n781), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n449), .A2(new_n404), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(G169gat), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n857), .A2(new_n858), .A3(new_n589), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n723), .A2(new_n405), .ZN(new_n860));
  AND4_X1   g659(.A1(new_n326), .A2(new_n806), .A3(new_n446), .A4(new_n860), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n861), .A2(new_n589), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n859), .B1(new_n862), .B2(new_n858), .ZN(G1348gat));
  AOI21_X1  g662(.A(G176gat), .B1(new_n857), .B2(new_n624), .ZN(new_n864));
  AND2_X1   g663(.A1(new_n861), .A2(new_n624), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n864), .B1(new_n865), .B2(G176gat), .ZN(G1349gat));
  AOI21_X1  g665(.A(new_n212), .B1(new_n861), .B2(new_n797), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n857), .A2(new_n221), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n867), .B1(new_n797), .B2(new_n868), .ZN(new_n869));
  XOR2_X1   g668(.A(new_n869), .B(KEYINPUT60), .Z(G1350gat));
  NAND3_X1  g669(.A1(new_n857), .A2(new_n213), .A3(new_n566), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT61), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n861), .A2(new_n566), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n872), .B1(new_n873), .B2(G190gat), .ZN(new_n874));
  AOI211_X1 g673(.A(KEYINPUT61), .B(new_n213), .C1(new_n861), .C2(new_n566), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n871), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  XNOR2_X1  g675(.A(new_n876), .B(KEYINPUT123), .ZN(G1351gat));
  NAND2_X1  g676(.A1(new_n822), .A2(new_n404), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(KEYINPUT124), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n855), .A2(new_n880), .ZN(new_n881));
  OR2_X1    g680(.A1(new_n879), .A2(KEYINPUT124), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(G197gat), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n884), .A2(new_n885), .A3(new_n589), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n639), .A2(new_n860), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n838), .A2(new_n836), .A3(new_n839), .ZN(new_n888));
  OAI21_X1  g687(.A(KEYINPUT122), .B1(new_n812), .B2(KEYINPUT57), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n887), .B1(new_n890), .B2(new_n835), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n891), .A2(new_n589), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n886), .B1(new_n892), .B2(new_n885), .ZN(G1352gat));
  NOR3_X1   g692(.A1(new_n883), .A2(G204gat), .A3(new_n687), .ZN(new_n894));
  NAND2_X1  g693(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  XOR2_X1   g695(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n897));
  NOR3_X1   g696(.A1(new_n843), .A2(new_n687), .A3(new_n887), .ZN(new_n898));
  OAI221_X1 g697(.A(new_n896), .B1(new_n894), .B2(new_n897), .C1(new_n615), .C2(new_n898), .ZN(G1353gat));
  NAND3_X1  g698(.A1(new_n884), .A2(new_n281), .A3(new_n797), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT63), .ZN(new_n901));
  AOI211_X1 g700(.A(new_n901), .B(new_n281), .C1(new_n891), .C2(new_n797), .ZN(new_n902));
  INV_X1    g701(.A(new_n887), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n842), .A2(new_n797), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(KEYINPUT63), .B1(new_n904), .B2(G211gat), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n900), .B1(new_n902), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(KEYINPUT126), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT126), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n908), .B(new_n900), .C1(new_n902), .C2(new_n905), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n907), .A2(new_n909), .ZN(G1354gat));
  NAND3_X1  g709(.A1(new_n884), .A2(new_n282), .A3(new_n566), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n891), .A2(new_n566), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n911), .B1(new_n912), .B2(new_n282), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n913), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


