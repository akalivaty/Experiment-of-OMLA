//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 1 0 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 0 1 0 1 1 1 1 0 0 0 1 0 0 1 0 1 1 0 0 1 1 0 1 1 0 0 0 1 0 0 0 1 1 1 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:13 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  OR2_X1    g001(.A1(KEYINPUT2), .A2(G113), .ZN(new_n188));
  NAND2_X1  g002(.A1(KEYINPUT2), .A2(G113), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT67), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  AOI21_X1  g005(.A(KEYINPUT67), .B1(KEYINPUT2), .B2(G113), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n188), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G119), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G116), .ZN(new_n195));
  INV_X1    g009(.A(G116), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G119), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n193), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT68), .ZN(new_n200));
  OAI211_X1 g014(.A(new_n200), .B(new_n188), .C1(new_n191), .C2(new_n192), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT69), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n198), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g017(.A(G116), .B(G119), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT69), .ZN(new_n205));
  AND3_X1   g019(.A1(new_n201), .A2(new_n203), .A3(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n193), .A2(KEYINPUT68), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n199), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT64), .ZN(new_n209));
  INV_X1    g023(.A(G137), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n209), .B1(new_n210), .B2(G134), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT11), .ZN(new_n212));
  INV_X1    g026(.A(G134), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n212), .B1(new_n213), .B2(G137), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(KEYINPUT64), .A3(G137), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n210), .A2(KEYINPUT11), .A3(G134), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n211), .A2(new_n214), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G131), .ZN(new_n218));
  AND4_X1   g032(.A1(new_n211), .A2(new_n214), .A3(new_n215), .A4(new_n216), .ZN(new_n219));
  INV_X1    g033(.A(G131), .ZN(new_n220));
  AOI21_X1  g034(.A(KEYINPUT65), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT65), .ZN(new_n222));
  NOR3_X1   g036(.A1(new_n217), .A2(new_n222), .A3(G131), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n218), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g038(.A(G143), .B(G146), .ZN(new_n225));
  NAND2_X1  g039(.A1(KEYINPUT0), .A2(G128), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  XOR2_X1   g041(.A(KEYINPUT0), .B(G128), .Z(new_n228));
  OAI21_X1  g042(.A(new_n227), .B1(new_n228), .B2(new_n225), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n224), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G146), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G143), .ZN(new_n232));
  INV_X1    g046(.A(G143), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G146), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n232), .A2(KEYINPUT1), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n235), .A2(new_n236), .A3(G128), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n210), .A2(G134), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n213), .A2(G137), .ZN(new_n239));
  OAI21_X1  g053(.A(G131), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G128), .ZN(new_n241));
  OAI211_X1 g055(.A(new_n232), .B(new_n234), .C1(KEYINPUT1), .C2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n237), .A2(new_n240), .A3(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n244), .B1(new_n221), .B2(new_n223), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n208), .B1(new_n230), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n229), .ZN(new_n247));
  AND2_X1   g061(.A1(new_n211), .A2(new_n215), .ZN(new_n248));
  AND2_X1   g062(.A1(new_n214), .A2(new_n216), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n248), .A2(new_n249), .A3(KEYINPUT65), .A4(new_n220), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n222), .B1(new_n217), .B2(G131), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n247), .B1(new_n252), .B2(new_n218), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n189), .B(new_n190), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n254), .A2(new_n188), .A3(new_n204), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n201), .A2(new_n203), .A3(new_n205), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n200), .B1(new_n254), .B2(new_n188), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n243), .B1(new_n251), .B2(new_n250), .ZN(new_n259));
  NOR3_X1   g073(.A1(new_n253), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  OAI21_X1  g074(.A(KEYINPUT28), .B1(new_n246), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT74), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AOI22_X1  g077(.A1(new_n250), .A2(new_n251), .B1(G131), .B2(new_n217), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n245), .B(new_n208), .C1(new_n264), .C2(new_n247), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT73), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT28), .ZN(new_n267));
  AND3_X1   g081(.A1(new_n265), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n266), .B1(new_n265), .B2(new_n267), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  XOR2_X1   g084(.A(KEYINPUT26), .B(G101), .Z(new_n271));
  NOR2_X1   g085(.A1(G237), .A2(G953), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G210), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT27), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n273), .B(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT70), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n273), .B(KEYINPUT27), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n278), .A2(KEYINPUT70), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n271), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(KEYINPUT70), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n275), .A2(new_n276), .ZN(new_n282));
  INV_X1    g096(.A(new_n271), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n281), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n280), .A2(new_n284), .ZN(new_n285));
  OAI211_X1 g099(.A(KEYINPUT74), .B(KEYINPUT28), .C1(new_n246), .C2(new_n260), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n263), .A2(new_n270), .A3(new_n285), .A4(new_n286), .ZN(new_n287));
  AND2_X1   g101(.A1(new_n287), .A2(KEYINPUT29), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n224), .A2(KEYINPUT66), .A3(new_n229), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT66), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n290), .B1(new_n264), .B2(new_n247), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT30), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n289), .A2(new_n291), .A3(new_n292), .A4(new_n245), .ZN(new_n293));
  OAI21_X1  g107(.A(KEYINPUT30), .B1(new_n253), .B2(new_n259), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n208), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n284), .B(new_n280), .C1(new_n295), .C2(new_n260), .ZN(new_n296));
  INV_X1    g110(.A(new_n268), .ZN(new_n297));
  INV_X1    g111(.A(new_n269), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n289), .A2(new_n291), .A3(new_n245), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n260), .B1(new_n299), .B2(new_n258), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n297), .B(new_n298), .C1(new_n300), .C2(new_n267), .ZN(new_n301));
  XNOR2_X1  g115(.A(new_n285), .B(KEYINPUT72), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT29), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n296), .B1(new_n301), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n187), .B1(new_n288), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G472), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT32), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT71), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n265), .A2(new_n285), .A3(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n309), .B1(new_n265), .B2(new_n285), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n293), .A2(new_n294), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(new_n258), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n313), .A2(new_n315), .A3(KEYINPUT31), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT31), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n265), .A2(new_n285), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(KEYINPUT71), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(new_n310), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n317), .B1(new_n320), .B2(new_n295), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n316), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n302), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n301), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g138(.A(G902), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G472), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n308), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  AOI22_X1  g141(.A1(new_n316), .A2(new_n321), .B1(new_n301), .B2(new_n323), .ZN(new_n328));
  NOR4_X1   g142(.A1(new_n328), .A2(KEYINPUT32), .A3(G472), .A4(G902), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n307), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(KEYINPUT75), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT79), .ZN(new_n332));
  XNOR2_X1  g146(.A(G125), .B(G140), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n332), .B1(new_n333), .B2(new_n231), .ZN(new_n334));
  INV_X1    g148(.A(G125), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G140), .ZN(new_n336));
  INV_X1    g150(.A(G140), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G125), .ZN(new_n338));
  AND4_X1   g152(.A1(new_n332), .A2(new_n336), .A3(new_n338), .A4(new_n231), .ZN(new_n339));
  OR2_X1    g153(.A1(new_n334), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT92), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT77), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n336), .A2(new_n338), .A3(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n335), .A2(KEYINPUT77), .A3(G140), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n341), .B1(new_n345), .B2(new_n231), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n343), .A2(KEYINPUT92), .A3(G146), .A4(new_n344), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n340), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(G214), .ZN(new_n349));
  NOR3_X1   g163(.A1(new_n349), .A2(G237), .A3(G953), .ZN(new_n350));
  OAI21_X1  g164(.A(KEYINPUT90), .B1(new_n350), .B2(G143), .ZN(new_n351));
  INV_X1    g165(.A(G237), .ZN(new_n352));
  INV_X1    g166(.A(G953), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n352), .A2(new_n353), .A3(G214), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT90), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(new_n355), .A3(new_n233), .ZN(new_n356));
  AOI22_X1  g170(.A1(new_n351), .A2(new_n356), .B1(G143), .B2(new_n350), .ZN(new_n357));
  NAND2_X1  g171(.A1(KEYINPUT18), .A2(G131), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NOR3_X1   g173(.A1(new_n357), .A2(KEYINPUT91), .A3(new_n358), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT91), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n350), .A2(G143), .ZN(new_n362));
  AOI211_X1 g176(.A(KEYINPUT90), .B(G143), .C1(new_n272), .C2(G214), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n355), .B1(new_n354), .B2(new_n233), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n362), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n358), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n361), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n348), .B(new_n359), .C1(new_n360), .C2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n365), .A2(G131), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT17), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n220), .B(new_n362), .C1(new_n363), .C2(new_n364), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n365), .A2(KEYINPUT17), .A3(G131), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT78), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n338), .A2(KEYINPUT16), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n376), .B1(new_n345), .B2(KEYINPUT16), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n375), .B1(new_n377), .B2(G146), .ZN(new_n378));
  INV_X1    g192(.A(new_n376), .ZN(new_n379));
  AND3_X1   g193(.A1(new_n335), .A2(KEYINPUT77), .A3(G140), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n380), .B1(new_n333), .B2(new_n342), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT16), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n379), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n383), .A2(KEYINPUT78), .A3(new_n231), .ZN(new_n384));
  OAI211_X1 g198(.A(G146), .B(new_n379), .C1(new_n381), .C2(new_n382), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n378), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n368), .B1(new_n374), .B2(new_n386), .ZN(new_n387));
  XNOR2_X1  g201(.A(G113), .B(G122), .ZN(new_n388));
  INV_X1    g202(.A(G104), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n388), .B(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n387), .A2(new_n391), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n368), .B(new_n390), .C1(new_n374), .C2(new_n386), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(new_n187), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G475), .ZN(new_n396));
  NAND2_X1  g210(.A1(KEYINPUT94), .A2(KEYINPUT15), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  NOR2_X1   g212(.A1(KEYINPUT94), .A2(KEYINPUT15), .ZN(new_n399));
  OAI21_X1  g213(.A(G478), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(G107), .ZN(new_n401));
  OR2_X1    g215(.A1(new_n196), .A2(G122), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n401), .B1(new_n402), .B2(KEYINPUT14), .ZN(new_n403));
  XNOR2_X1  g217(.A(G116), .B(G122), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  OR2_X1    g219(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n403), .A2(new_n405), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n241), .A2(G143), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n409), .B(KEYINPUT93), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n233), .A2(G128), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(G134), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n410), .A2(new_n213), .A3(new_n411), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n408), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n404), .B(new_n401), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n411), .B(KEYINPUT13), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n213), .B1(new_n410), .B2(new_n419), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  XOR2_X1   g236(.A(KEYINPUT76), .B(G217), .Z(new_n423));
  XNOR2_X1  g237(.A(KEYINPUT9), .B(G234), .ZN(new_n424));
  NOR3_X1   g238(.A1(new_n423), .A2(G953), .A3(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n416), .A2(new_n422), .A3(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n425), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n427), .B1(new_n415), .B2(new_n421), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n400), .B1(new_n429), .B2(new_n187), .ZN(new_n430));
  INV_X1    g244(.A(new_n400), .ZN(new_n431));
  AOI211_X1 g245(.A(G902), .B(new_n431), .C1(new_n426), .C2(new_n428), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT20), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n347), .B1(new_n334), .B2(new_n339), .ZN(new_n435));
  AOI21_X1  g249(.A(KEYINPUT92), .B1(new_n381), .B2(G146), .ZN(new_n436));
  OAI22_X1  g250(.A1(new_n435), .A2(new_n436), .B1(new_n365), .B2(new_n366), .ZN(new_n437));
  INV_X1    g251(.A(new_n367), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n365), .A2(new_n361), .A3(new_n366), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n437), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT19), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n333), .A2(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n442), .B1(new_n345), .B2(new_n441), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n385), .B1(G146), .B2(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n444), .B1(new_n369), .B2(new_n371), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n391), .B1(new_n440), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n393), .ZN(new_n447));
  NOR2_X1   g261(.A1(G475), .A2(G902), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n434), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n448), .ZN(new_n450));
  AOI211_X1 g264(.A(KEYINPUT20), .B(new_n450), .C1(new_n446), .C2(new_n393), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n396), .B(new_n433), .C1(new_n449), .C2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n353), .A2(G952), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n453), .B1(G234), .B2(G237), .ZN(new_n454));
  NAND2_X1  g268(.A1(G234), .A2(G237), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n455), .A2(G902), .A3(G953), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(KEYINPUT21), .B(G898), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n454), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(KEYINPUT95), .B1(new_n452), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(G475), .ZN(new_n461));
  AOI21_X1  g275(.A(G902), .B1(new_n392), .B2(new_n393), .ZN(new_n462));
  OAI22_X1  g276(.A1(new_n449), .A2(new_n451), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT95), .ZN(new_n465));
  INV_X1    g279(.A(new_n459), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n464), .A2(new_n465), .A3(new_n466), .A4(new_n433), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n460), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(G221), .ZN(new_n469));
  INV_X1    g283(.A(new_n424), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n469), .B1(new_n470), .B2(new_n187), .ZN(new_n471));
  XOR2_X1   g285(.A(KEYINPUT83), .B(G469), .Z(new_n472));
  XNOR2_X1  g286(.A(G110), .B(G140), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n473), .B(KEYINPUT80), .ZN(new_n474));
  AND2_X1   g288(.A1(new_n353), .A2(G227), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n474), .B(new_n475), .ZN(new_n476));
  AND2_X1   g290(.A1(KEYINPUT81), .A2(G104), .ZN(new_n477));
  NOR2_X1   g291(.A1(KEYINPUT81), .A2(G104), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(KEYINPUT3), .B1(new_n479), .B2(G107), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT3), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n481), .A2(new_n401), .A3(G104), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT82), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n481), .A2(new_n401), .A3(KEYINPUT82), .A4(G104), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(G101), .ZN(new_n487));
  INV_X1    g301(.A(new_n478), .ZN(new_n488));
  NAND2_X1  g302(.A1(KEYINPUT81), .A2(G104), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n488), .A2(G107), .A3(new_n489), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n480), .A2(new_n486), .A3(new_n487), .A4(new_n490), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n479), .A2(G107), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n401), .A2(G104), .ZN(new_n493));
  OAI21_X1  g307(.A(G101), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n237), .A2(new_n242), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(KEYINPUT10), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n389), .A2(KEYINPUT3), .ZN(new_n499));
  AOI21_X1  g313(.A(KEYINPUT82), .B1(new_n499), .B2(new_n401), .ZN(new_n500));
  INV_X1    g314(.A(new_n485), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n490), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n488), .A2(new_n489), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n481), .B1(new_n503), .B2(new_n401), .ZN(new_n504));
  OAI21_X1  g318(.A(G101), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n505), .A2(KEYINPUT4), .A3(new_n491), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT4), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n507), .B(G101), .C1(new_n502), .C2(new_n504), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n506), .A2(new_n229), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT10), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n510), .B1(new_n495), .B2(new_n496), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n498), .A2(new_n509), .A3(new_n264), .A4(new_n511), .ZN(new_n512));
  AOI22_X1  g326(.A1(new_n491), .A2(new_n494), .B1(new_n242), .B2(new_n237), .ZN(new_n513));
  OR2_X1    g327(.A1(new_n497), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(KEYINPUT12), .B1(new_n514), .B2(new_n224), .ZN(new_n515));
  OAI211_X1 g329(.A(KEYINPUT12), .B(new_n224), .C1(new_n497), .C2(new_n513), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n476), .B(new_n512), .C1(new_n515), .C2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n498), .A2(new_n509), .A3(new_n511), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(new_n224), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n476), .B1(new_n520), .B2(new_n512), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT84), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n518), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AOI211_X1 g337(.A(KEYINPUT84), .B(new_n476), .C1(new_n520), .C2(new_n512), .ZN(new_n524));
  OAI211_X1 g338(.A(new_n187), .B(new_n472), .C1(new_n523), .C2(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n512), .B1(new_n515), .B2(new_n517), .ZN(new_n526));
  INV_X1    g340(.A(new_n476), .ZN(new_n527));
  AND2_X1   g341(.A1(new_n512), .A2(new_n476), .ZN(new_n528));
  AOI22_X1  g342(.A1(new_n526), .A2(new_n527), .B1(new_n528), .B2(new_n520), .ZN(new_n529));
  OAI21_X1  g343(.A(G469), .B1(new_n529), .B2(G902), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n471), .B1(new_n525), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(G214), .B1(G237), .B2(G902), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  AND3_X1   g347(.A1(new_n505), .A2(KEYINPUT4), .A3(new_n491), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n258), .A2(new_n508), .ZN(new_n535));
  OAI21_X1  g349(.A(KEYINPUT85), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT85), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n506), .A2(new_n537), .A3(new_n258), .A4(new_n508), .ZN(new_n538));
  AND3_X1   g352(.A1(new_n195), .A2(new_n197), .A3(KEYINPUT69), .ZN(new_n539));
  AOI21_X1  g353(.A(KEYINPUT69), .B1(new_n195), .B2(new_n197), .ZN(new_n540));
  OAI21_X1  g354(.A(KEYINPUT5), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n195), .A2(KEYINPUT5), .ZN(new_n542));
  INV_X1    g356(.A(G113), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n199), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n545), .A2(new_n491), .A3(new_n494), .ZN(new_n546));
  XNOR2_X1  g360(.A(G110), .B(G122), .ZN(new_n547));
  AND4_X1   g361(.A1(new_n536), .A2(new_n538), .A3(new_n546), .A4(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n229), .A2(G125), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n549), .B1(G125), .B2(new_n496), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n353), .A2(G224), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(KEYINPUT7), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n550), .B(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT88), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n495), .A2(new_n545), .ZN(new_n555));
  AOI211_X1 g369(.A(new_n543), .B(new_n542), .C1(KEYINPUT5), .C2(new_n204), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n491), .B(new_n494), .C1(new_n556), .C2(new_n199), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n547), .B(KEYINPUT8), .ZN(new_n558));
  AND4_X1   g372(.A1(new_n554), .A2(new_n555), .A3(new_n557), .A4(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n558), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n560), .B1(new_n495), .B2(new_n545), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n554), .B1(new_n561), .B2(new_n557), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n553), .B1(new_n559), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n187), .B1(new_n548), .B2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT89), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n547), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n538), .A2(new_n546), .ZN(new_n568));
  AND2_X1   g382(.A1(new_n258), .A2(new_n508), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n537), .B1(new_n569), .B2(new_n506), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n567), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n536), .A2(new_n538), .A3(new_n546), .A4(new_n547), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT6), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n573), .A2(KEYINPUT86), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n571), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT87), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n550), .B(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(new_n551), .ZN(new_n578));
  OAI221_X1 g392(.A(new_n567), .B1(KEYINPUT86), .B2(new_n573), .C1(new_n568), .C2(new_n570), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n575), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  OAI211_X1 g394(.A(KEYINPUT89), .B(new_n187), .C1(new_n548), .C2(new_n563), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n566), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  OAI21_X1  g396(.A(G210), .B1(G237), .B2(G902), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n566), .A2(new_n580), .A3(new_n583), .A4(new_n581), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n533), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n468), .A2(new_n531), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n241), .A2(G119), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT23), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n241), .A2(KEYINPUT23), .A3(G119), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n194), .A2(G128), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(G110), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n589), .A2(new_n593), .ZN(new_n596));
  XNOR2_X1  g410(.A(KEYINPUT24), .B(G110), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n386), .B(new_n595), .C1(new_n596), .C2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n596), .A2(new_n597), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n599), .B1(new_n594), .B2(G110), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n385), .A2(new_n340), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(KEYINPUT22), .B(G137), .ZN(new_n603));
  AND3_X1   g417(.A1(new_n353), .A2(G221), .A3(G234), .ZN(new_n604));
  XOR2_X1   g418(.A(new_n603), .B(new_n604), .Z(new_n605));
  NAND2_X1  g419(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n605), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n598), .A2(new_n601), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(G902), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT25), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n423), .B1(G234), .B2(new_n187), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n614), .B1(new_n609), .B2(new_n610), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n606), .A2(new_n608), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n613), .A2(G902), .ZN(new_n617));
  AOI22_X1  g431(.A1(new_n612), .A2(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT75), .ZN(new_n619));
  OAI211_X1 g433(.A(new_n307), .B(new_n619), .C1(new_n327), .C2(new_n329), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n331), .A2(new_n588), .A3(new_n618), .A4(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(G101), .ZN(G3));
  NAND2_X1  g436(.A1(new_n585), .A2(new_n586), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n532), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n624), .A2(new_n459), .ZN(new_n625));
  AOI211_X1 g439(.A(G478), .B(G902), .C1(new_n426), .C2(new_n428), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n429), .A2(KEYINPUT33), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT33), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n628), .B1(new_n426), .B2(new_n428), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n187), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n626), .B1(new_n630), .B2(G478), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n463), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n625), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n325), .A2(new_n326), .ZN(new_n635));
  OAI21_X1  g449(.A(G472), .B1(new_n328), .B2(G902), .ZN(new_n636));
  AND4_X1   g450(.A1(new_n618), .A2(new_n531), .A3(new_n635), .A4(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(KEYINPUT96), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT34), .B(G104), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G6));
  OR2_X1    g456(.A1(new_n430), .A2(new_n432), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n464), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n625), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n646), .A2(new_n638), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT35), .B(G107), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G9));
  AND2_X1   g463(.A1(new_n635), .A2(new_n636), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n607), .A2(KEYINPUT36), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n602), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n617), .ZN(new_n653));
  INV_X1    g467(.A(new_n615), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n653), .B1(new_n654), .B2(new_n611), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n588), .A2(new_n650), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT37), .B(G110), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G12));
  AND2_X1   g472(.A1(new_n331), .A2(new_n620), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n531), .A2(new_n655), .ZN(new_n660));
  INV_X1    g474(.A(G900), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n457), .A2(KEYINPUT97), .A3(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n454), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT97), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n664), .B1(new_n456), .B2(G900), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n662), .A2(new_n663), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n645), .A2(new_n666), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n624), .A2(new_n660), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n659), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G128), .ZN(G30));
  XNOR2_X1  g484(.A(new_n666), .B(KEYINPUT39), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n531), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(new_n672), .B(KEYINPUT40), .Z(new_n673));
  XOR2_X1   g487(.A(new_n623), .B(KEYINPUT38), .Z(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  OR2_X1    g489(.A1(new_n327), .A2(new_n329), .ZN(new_n676));
  OR2_X1    g490(.A1(new_n246), .A2(new_n260), .ZN(new_n677));
  AOI22_X1  g491(.A1(new_n315), .A2(new_n313), .B1(new_n323), .B2(new_n677), .ZN(new_n678));
  OAI21_X1  g492(.A(G472), .B1(new_n678), .B2(G902), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n463), .A2(new_n643), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n655), .A2(new_n681), .A3(new_n533), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n673), .A2(new_n675), .A3(new_n680), .A4(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(new_n683), .B(KEYINPUT98), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G143), .ZN(G45));
  NAND2_X1  g499(.A1(new_n633), .A2(new_n666), .ZN(new_n686));
  NOR3_X1   g500(.A1(new_n624), .A2(new_n660), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n659), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G146), .ZN(G48));
  AND3_X1   g503(.A1(new_n331), .A2(new_n618), .A3(new_n620), .ZN(new_n690));
  INV_X1    g504(.A(new_n634), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n187), .B1(new_n523), .B2(new_n524), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(G469), .ZN(new_n693));
  INV_X1    g507(.A(new_n471), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n693), .A2(new_n694), .A3(new_n525), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n690), .A2(KEYINPUT99), .A3(new_n691), .A4(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT99), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n331), .A2(new_n618), .A3(new_n620), .A4(new_n696), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n698), .B1(new_n699), .B2(new_n634), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(KEYINPUT41), .B(G113), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G15));
  NOR2_X1   g517(.A1(new_n699), .A2(new_n646), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(new_n196), .ZN(G18));
  NOR2_X1   g519(.A1(new_n624), .A2(new_n695), .ZN(new_n706));
  INV_X1    g520(.A(new_n655), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n707), .B1(new_n460), .B2(new_n467), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n331), .A2(new_n620), .A3(new_n706), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G119), .ZN(G21));
  NOR2_X1   g524(.A1(new_n624), .A2(new_n681), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n263), .A2(new_n270), .A3(new_n286), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(KEYINPUT100), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT100), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n263), .A2(new_n270), .A3(new_n714), .A4(new_n286), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n302), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n322), .ZN(new_n717));
  OAI211_X1 g531(.A(new_n326), .B(new_n187), .C1(new_n716), .C2(new_n717), .ZN(new_n718));
  AND3_X1   g532(.A1(new_n718), .A2(new_n618), .A3(new_n636), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n711), .A2(new_n719), .A3(new_n466), .A4(new_n696), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G122), .ZN(G24));
  INV_X1    g535(.A(new_n666), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n632), .A2(new_n722), .ZN(new_n723));
  AND4_X1   g537(.A1(new_n636), .A2(new_n718), .A3(new_n723), .A4(new_n655), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n724), .A2(KEYINPUT101), .A3(new_n706), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT101), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n696), .A2(new_n587), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n718), .A2(new_n723), .A3(new_n636), .A4(new_n655), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n726), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n725), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G125), .ZN(G27));
  NAND4_X1  g545(.A1(new_n585), .A2(new_n694), .A3(new_n532), .A4(new_n586), .ZN(new_n732));
  NAND2_X1  g546(.A1(G469), .A2(G902), .ZN(new_n733));
  XOR2_X1   g547(.A(new_n733), .B(KEYINPUT102), .Z(new_n734));
  AOI21_X1  g548(.A(new_n734), .B1(new_n529), .B2(G469), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n525), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n732), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n723), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n330), .A2(new_n618), .ZN(new_n739));
  OAI21_X1  g553(.A(KEYINPUT42), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n331), .A2(new_n618), .A3(new_n620), .A4(new_n737), .ZN(new_n741));
  OR2_X1    g555(.A1(new_n686), .A2(KEYINPUT42), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n740), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(new_n220), .ZN(G33));
  OR2_X1    g558(.A1(new_n741), .A2(new_n667), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G134), .ZN(G36));
  INV_X1    g560(.A(KEYINPUT103), .ZN(new_n747));
  INV_X1    g561(.A(G469), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT45), .ZN(new_n749));
  OR2_X1    g563(.A1(new_n529), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n529), .A2(new_n749), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n748), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  OR2_X1    g566(.A1(new_n752), .A2(new_n734), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT46), .ZN(new_n754));
  OAI211_X1 g568(.A(new_n747), .B(new_n525), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n752), .A2(new_n754), .A3(new_n734), .ZN(new_n756));
  INV_X1    g570(.A(new_n525), .ZN(new_n757));
  OAI21_X1  g571(.A(KEYINPUT103), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n753), .A2(new_n754), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n755), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n760), .A2(new_n694), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n761), .A2(new_n671), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n585), .A2(new_n532), .A3(new_n586), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n464), .A2(new_n631), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(KEYINPUT43), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n765), .A2(new_n650), .A3(new_n707), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n763), .B1(new_n766), .B2(KEYINPUT44), .ZN(new_n767));
  OAI211_X1 g581(.A(new_n762), .B(new_n767), .C1(KEYINPUT44), .C2(new_n766), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G137), .ZN(G39));
  NOR4_X1   g583(.A1(new_n659), .A2(new_n618), .A3(new_n686), .A4(new_n763), .ZN(new_n770));
  AND3_X1   g584(.A1(new_n760), .A2(KEYINPUT47), .A3(new_n694), .ZN(new_n771));
  AOI21_X1  g585(.A(KEYINPUT47), .B1(new_n760), .B2(new_n694), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n770), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G140), .ZN(G42));
  NOR2_X1   g588(.A1(new_n771), .A2(new_n772), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n693), .A2(new_n471), .A3(new_n525), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(KEYINPUT110), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n765), .A2(new_n663), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n779), .A2(new_n719), .ZN(new_n780));
  INV_X1    g594(.A(new_n763), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(KEYINPUT51), .B1(new_n778), .B2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT112), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT50), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n696), .A2(new_n533), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT111), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n674), .A2(new_n779), .A3(new_n719), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n785), .B(new_n786), .C1(new_n789), .C2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n787), .B(KEYINPUT111), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n785), .A2(new_n786), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n792), .A2(new_n780), .A3(new_n674), .A4(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n718), .A2(new_n636), .A3(new_n655), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n693), .A2(new_n525), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n732), .A2(new_n797), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n779), .A2(new_n796), .A3(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n680), .ZN(new_n800));
  AND4_X1   g614(.A1(new_n618), .A2(new_n800), .A3(new_n454), .A4(new_n798), .ZN(new_n801));
  OR2_X1    g615(.A1(new_n631), .A2(new_n463), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n799), .B1(new_n801), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n795), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n805), .A2(KEYINPUT113), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT113), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n807), .B1(new_n795), .B2(new_n804), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n784), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n782), .B1(new_n775), .B2(new_n776), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT114), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n805), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n795), .A2(KEYINPUT114), .A3(new_n804), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n810), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT51), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n809), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n739), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n817), .A2(new_n779), .A3(new_n798), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(KEYINPUT48), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n801), .A2(new_n633), .ZN(new_n820));
  XOR2_X1   g634(.A(new_n453), .B(KEYINPUT115), .Z(new_n821));
  AOI21_X1  g635(.A(new_n821), .B1(new_n780), .B2(new_n706), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n819), .A2(new_n820), .A3(new_n822), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n816), .A2(KEYINPUT116), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(KEYINPUT116), .B1(new_n816), .B2(new_n823), .ZN(new_n825));
  OR2_X1    g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n463), .A2(new_n643), .A3(new_n722), .ZN(new_n827));
  AND4_X1   g641(.A1(new_n532), .A2(new_n827), .A3(new_n585), .A4(new_n586), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n660), .B1(new_n828), .B2(KEYINPUT104), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT104), .ZN(new_n830));
  INV_X1    g644(.A(new_n827), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n830), .B1(new_n763), .B2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n829), .A2(new_n331), .A3(new_n620), .A4(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n724), .A2(new_n737), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n833), .B(new_n834), .C1(new_n741), .C2(new_n667), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n625), .B(new_n637), .C1(new_n633), .C2(new_n645), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n621), .A2(new_n656), .A3(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n743), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n709), .B(new_n720), .C1(new_n699), .C2(new_n646), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n838), .A2(new_n701), .A3(new_n839), .A4(new_n841), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(KEYINPUT105), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n331), .B(new_n620), .C1(new_n668), .C2(new_n687), .ZN(new_n845));
  NOR4_X1   g659(.A1(new_n736), .A2(new_n655), .A3(new_n471), .A4(new_n722), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n680), .A2(new_n711), .A3(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n845), .A2(new_n730), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT52), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT52), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n845), .A2(new_n730), .A3(new_n850), .A4(new_n847), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT106), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n849), .A2(KEYINPUT106), .A3(new_n851), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n843), .A2(new_n844), .A3(new_n856), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n835), .A2(new_n743), .A3(new_n837), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n840), .B1(new_n700), .B2(new_n697), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n858), .A2(new_n859), .A3(new_n849), .A4(new_n851), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(KEYINPUT53), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n857), .A2(KEYINPUT54), .A3(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT107), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n857), .A2(KEYINPUT107), .A3(KEYINPUT54), .A4(new_n861), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n858), .A2(new_n859), .A3(KEYINPUT53), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n866), .B1(new_n854), .B2(new_n855), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n844), .B1(new_n842), .B2(new_n852), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT108), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n860), .A2(KEYINPUT108), .A3(new_n844), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n867), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  XOR2_X1   g686(.A(KEYINPUT109), .B(KEYINPUT54), .Z(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n864), .A2(new_n865), .A3(new_n874), .ZN(new_n875));
  OAI22_X1  g689(.A1(new_n826), .A2(new_n875), .B1(G952), .B2(G953), .ZN(new_n876));
  XOR2_X1   g690(.A(new_n797), .B(KEYINPUT49), .Z(new_n877));
  NAND3_X1  g691(.A1(new_n618), .A2(new_n694), .A3(new_n532), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n878), .A2(new_n764), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n800), .A2(new_n877), .A3(new_n674), .A4(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n876), .A2(new_n880), .ZN(G75));
  INV_X1    g695(.A(new_n866), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n856), .A2(new_n882), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n860), .A2(KEYINPUT108), .A3(new_n844), .ZN(new_n884));
  AOI21_X1  g698(.A(KEYINPUT108), .B1(new_n860), .B2(new_n844), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n886), .A2(G210), .A3(G902), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT117), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT56), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n575), .A2(new_n579), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(new_n578), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(KEYINPUT55), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n887), .A2(new_n888), .A3(new_n889), .A4(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n353), .A2(G952), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n887), .A2(new_n889), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n892), .B1(new_n897), .B2(new_n888), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n888), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n896), .B1(new_n898), .B2(new_n899), .ZN(G51));
  XNOR2_X1  g714(.A(new_n886), .B(new_n873), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n734), .B(KEYINPUT57), .Z(new_n902));
  OAI22_X1  g716(.A1(new_n901), .A2(new_n902), .B1(new_n524), .B2(new_n523), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n886), .A2(G902), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(new_n752), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n894), .B1(new_n903), .B2(new_n906), .ZN(G54));
  NAND4_X1  g721(.A1(new_n905), .A2(KEYINPUT58), .A3(G475), .A4(new_n447), .ZN(new_n908));
  NAND2_X1  g722(.A1(KEYINPUT58), .A2(G475), .ZN(new_n909));
  OAI211_X1 g723(.A(new_n393), .B(new_n446), .C1(new_n904), .C2(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n908), .A2(new_n910), .A3(new_n895), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT118), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n908), .A2(new_n910), .A3(KEYINPUT118), .A4(new_n895), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(G60));
  OR2_X1    g729(.A1(new_n627), .A2(new_n629), .ZN(new_n916));
  NAND2_X1  g730(.A1(G478), .A2(G902), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT59), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n916), .B1(new_n875), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n916), .A2(new_n918), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n895), .B1(new_n901), .B2(new_n920), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n919), .A2(new_n921), .ZN(G63));
  INV_X1    g736(.A(KEYINPUT119), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT61), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT120), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n894), .B1(new_n923), .B2(new_n924), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(G217), .A2(G902), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT60), .Z(new_n931));
  NAND2_X1  g745(.A1(new_n886), .A2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(new_n616), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n929), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n886), .A2(new_n652), .A3(new_n931), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n927), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(new_n931), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n933), .B1(new_n872), .B2(new_n937), .ZN(new_n938));
  AND4_X1   g752(.A1(new_n927), .A2(new_n938), .A3(new_n935), .A4(new_n928), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n926), .B1(new_n936), .B2(new_n939), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n938), .A2(new_n935), .A3(new_n928), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(KEYINPUT120), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n934), .A2(new_n927), .A3(new_n935), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n942), .A2(new_n943), .A3(new_n925), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n940), .A2(new_n944), .ZN(G66));
  NAND2_X1  g759(.A1(G224), .A2(G953), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n458), .A2(new_n946), .ZN(new_n947));
  AOI211_X1 g761(.A(new_n837), .B(new_n840), .C1(new_n700), .C2(new_n697), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n947), .B1(new_n948), .B2(new_n353), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n890), .B1(G898), .B2(new_n353), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n949), .B(new_n950), .ZN(G69));
  INV_X1    g765(.A(KEYINPUT124), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n762), .A2(KEYINPUT123), .A3(new_n711), .A4(new_n817), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT123), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n761), .A2(new_n671), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n817), .A2(new_n711), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n953), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n839), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n845), .A2(new_n730), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n773), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n961), .A2(new_n768), .A3(new_n745), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n952), .B1(new_n959), .B2(new_n962), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n768), .A2(new_n745), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n743), .B1(new_n953), .B2(new_n957), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n964), .A2(new_n965), .A3(KEYINPUT124), .A4(new_n961), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n963), .A2(new_n353), .A3(new_n966), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n443), .B(KEYINPUT121), .Z(new_n968));
  XNOR2_X1  g782(.A(new_n314), .B(new_n968), .ZN(new_n969));
  OAI211_X1 g783(.A(new_n967), .B(new_n969), .C1(new_n661), .C2(new_n353), .ZN(new_n970));
  AOI211_X1 g784(.A(new_n763), .B(new_n672), .C1(new_n632), .C2(new_n644), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n690), .A2(new_n971), .ZN(new_n972));
  AND3_X1   g786(.A1(new_n768), .A2(new_n773), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(KEYINPUT62), .B1(new_n684), .B2(new_n960), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n684), .A2(KEYINPUT62), .A3(new_n960), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n973), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT122), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n973), .B(KEYINPUT122), .C1(new_n974), .C2(new_n975), .ZN(new_n979));
  AOI21_X1  g793(.A(G953), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n970), .B1(new_n980), .B2(new_n969), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n353), .B1(G227), .B2(G900), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(new_n982), .ZN(new_n984));
  OAI211_X1 g798(.A(new_n970), .B(new_n984), .C1(new_n980), .C2(new_n969), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n983), .A2(new_n985), .ZN(G72));
  NAND3_X1  g800(.A1(new_n978), .A2(new_n948), .A3(new_n979), .ZN(new_n987));
  XNOR2_X1  g801(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n326), .A2(new_n187), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n988), .B(new_n989), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(KEYINPUT126), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n987), .A2(new_n991), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n295), .A2(new_n260), .ZN(new_n993));
  INV_X1    g807(.A(new_n993), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n992), .A2(new_n285), .A3(new_n994), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n296), .B(KEYINPUT127), .Z(new_n996));
  NAND2_X1  g810(.A1(new_n313), .A2(new_n315), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n990), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n857), .A2(new_n861), .A3(new_n998), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n963), .A2(new_n948), .A3(new_n966), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n1000), .A2(new_n991), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n994), .A2(new_n285), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n894), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  AND3_X1   g817(.A1(new_n995), .A2(new_n999), .A3(new_n1003), .ZN(G57));
endmodule


