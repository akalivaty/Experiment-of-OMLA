//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 1 0 0 0 0 0 1 1 0 0 0 0 1 0 1 0 1 0 1 0 0 0 1 0 0 0 1 1 0 0 0 1 0 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n768, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n984, new_n985, new_n986, new_n987, new_n988;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT0), .ZN(new_n203));
  XNOR2_X1  g002(.A(G57gat), .B(G85gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT6), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n205), .A2(KEYINPUT6), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT79), .ZN(new_n212));
  XNOR2_X1  g011(.A(G155gat), .B(G162gat), .ZN(new_n213));
  XOR2_X1   g012(.A(G141gat), .B(G148gat), .Z(new_n214));
  INV_X1    g013(.A(KEYINPUT2), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT74), .ZN(new_n218));
  INV_X1    g017(.A(G141gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(KEYINPUT74), .A2(G141gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n220), .A2(G148gat), .A3(new_n221), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n219), .A2(G148gat), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(KEYINPUT75), .A2(G162gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT2), .ZN(new_n227));
  INV_X1    g026(.A(G162gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(G155gat), .ZN(new_n229));
  INV_X1    g028(.A(G155gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(G162gat), .ZN(new_n231));
  AND3_X1   g030(.A1(new_n227), .A2(new_n229), .A3(new_n231), .ZN(new_n232));
  AND3_X1   g031(.A1(new_n225), .A2(KEYINPUT76), .A3(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT76), .B1(new_n225), .B2(new_n232), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n217), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(G120gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(G113gat), .ZN(new_n237));
  INV_X1    g036(.A(G113gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(G120gat), .ZN(new_n239));
  AOI21_X1  g038(.A(KEYINPUT1), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(G127gat), .ZN(new_n241));
  INV_X1    g040(.A(G134gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(G127gat), .A2(G134gat), .ZN(new_n244));
  AND2_X1   g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT1), .ZN(new_n246));
  AND2_X1   g045(.A1(new_n246), .A2(KEYINPUT71), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n240), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  AOI22_X1  g047(.A1(new_n243), .A2(new_n244), .B1(KEYINPUT71), .B2(new_n246), .ZN(new_n249));
  AND2_X1   g048(.A1(new_n237), .A2(new_n239), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n249), .B1(new_n250), .B2(KEYINPUT1), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n235), .A2(new_n253), .ZN(new_n254));
  OAI211_X1 g053(.A(new_n252), .B(new_n217), .C1(new_n233), .C2(new_n234), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(G225gat), .A2(G233gat), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n212), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  AOI211_X1 g058(.A(KEYINPUT79), .B(new_n257), .C1(new_n254), .C2(new_n255), .ZN(new_n260));
  OAI21_X1  g059(.A(KEYINPUT5), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT78), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n255), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT76), .ZN(new_n265));
  AND2_X1   g064(.A1(KEYINPUT74), .A2(G141gat), .ZN(new_n266));
  NOR2_X1   g065(.A1(KEYINPUT74), .A2(G141gat), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n223), .B1(new_n268), .B2(G148gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n213), .A2(new_n227), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n265), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n225), .A2(new_n232), .A3(KEYINPUT76), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n216), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n273), .A2(KEYINPUT4), .A3(new_n252), .ZN(new_n274));
  AND3_X1   g073(.A1(new_n264), .A2(new_n274), .A3(new_n257), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT77), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT3), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n276), .B1(new_n273), .B2(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n252), .B1(new_n273), .B2(new_n277), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n235), .A2(KEYINPUT77), .A3(KEYINPUT3), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n262), .B1(new_n275), .B2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n275), .A2(new_n262), .A3(new_n281), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n261), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n264), .A2(new_n274), .A3(new_n286), .A4(new_n257), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n288), .A2(KEYINPUT80), .A3(new_n281), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT80), .ZN(new_n290));
  AND3_X1   g089(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n290), .B1(new_n291), .B2(new_n287), .ZN(new_n292));
  AND2_X1   g091(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  OAI211_X1 g092(.A(new_n209), .B(new_n211), .C1(new_n285), .C2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n255), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n271), .A2(new_n272), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n252), .B1(new_n296), .B2(new_n217), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n258), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT79), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n256), .A2(new_n212), .A3(new_n258), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n286), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  AND3_X1   g100(.A1(new_n275), .A2(new_n262), .A3(new_n281), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n301), .B1(new_n302), .B2(new_n282), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n289), .A2(new_n292), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n303), .A2(new_n207), .A3(new_n304), .A4(new_n206), .ZN(new_n305));
  OR2_X1    g104(.A1(KEYINPUT66), .A2(G176gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(KEYINPUT66), .A2(G176gat), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n306), .A2(KEYINPUT23), .A3(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(G169gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT65), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT65), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(G169gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(KEYINPUT67), .B1(new_n308), .B2(new_n313), .ZN(new_n314));
  AND2_X1   g113(.A1(KEYINPUT66), .A2(G176gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(KEYINPUT66), .A2(G176gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(KEYINPUT65), .B(G169gat), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT67), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n317), .A2(new_n318), .A3(new_n319), .A4(KEYINPUT23), .ZN(new_n320));
  NAND2_X1  g119(.A1(G169gat), .A2(G176gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(G183gat), .A2(G190gat), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n321), .B1(new_n322), .B2(KEYINPUT24), .ZN(new_n323));
  INV_X1    g122(.A(G183gat), .ZN(new_n324));
  INV_X1    g123(.A(G190gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  AND2_X1   g125(.A1(new_n322), .A2(KEYINPUT24), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n323), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G176gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n309), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT23), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n330), .A2(KEYINPUT68), .A3(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT68), .ZN(new_n333));
  NOR2_X1   g132(.A1(G169gat), .A2(G176gat), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n333), .B1(new_n334), .B2(KEYINPUT23), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n314), .A2(new_n320), .A3(new_n328), .A4(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  AND2_X1   g138(.A1(new_n328), .A2(new_n336), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT25), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n341), .B1(new_n334), .B2(KEYINPUT23), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  AND2_X1   g143(.A1(G226gat), .A2(G233gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(KEYINPUT27), .B(G183gat), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT28), .B1(new_n346), .B2(new_n325), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n324), .A2(KEYINPUT27), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT27), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(G183gat), .ZN(new_n350));
  AND4_X1   g149(.A1(KEYINPUT28), .A2(new_n348), .A3(new_n350), .A4(new_n325), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n322), .B1(new_n347), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n354), .A2(KEYINPUT69), .A3(new_n330), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT69), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n356), .B1(new_n353), .B2(new_n334), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT26), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n334), .A2(new_n358), .ZN(new_n359));
  AND3_X1   g158(.A1(new_n355), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(KEYINPUT70), .B1(new_n352), .B2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n348), .A2(new_n350), .A3(new_n325), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT28), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n346), .A2(KEYINPUT28), .A3(new_n325), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n355), .A2(new_n357), .A3(new_n359), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT70), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n366), .A2(new_n367), .A3(new_n368), .A4(new_n322), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n344), .A2(new_n345), .A3(new_n361), .A4(new_n369), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n345), .A2(KEYINPUT29), .ZN(new_n371));
  AOI22_X1  g170(.A1(new_n337), .A2(new_n338), .B1(new_n340), .B2(new_n342), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n352), .A2(new_n360), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n371), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n370), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n376));
  OR2_X1    g175(.A1(G197gat), .A2(G204gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(G197gat), .A2(G204gat), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n379), .B(KEYINPUT73), .ZN(new_n380));
  XOR2_X1   g179(.A(G211gat), .B(G218gat), .Z(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n379), .A2(KEYINPUT73), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(new_n381), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n375), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n361), .A2(new_n369), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n371), .B1(new_n388), .B2(new_n372), .ZN(new_n389));
  INV_X1    g188(.A(new_n386), .ZN(new_n390));
  INV_X1    g189(.A(new_n373), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n344), .A2(new_n391), .A3(new_n345), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n389), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT30), .ZN(new_n394));
  XNOR2_X1  g193(.A(G8gat), .B(G36gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(G64gat), .B(G92gat), .ZN(new_n396));
  XOR2_X1   g195(.A(new_n395), .B(new_n396), .Z(new_n397));
  NAND4_X1  g196(.A1(new_n387), .A2(new_n393), .A3(new_n394), .A4(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n397), .ZN(new_n399));
  AND3_X1   g198(.A1(new_n389), .A2(new_n390), .A3(new_n392), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n390), .B1(new_n370), .B2(new_n374), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n399), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n387), .A2(new_n393), .A3(new_n397), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n402), .A2(new_n403), .A3(KEYINPUT30), .ZN(new_n404));
  AOI22_X1  g203(.A1(new_n294), .A2(new_n305), .B1(new_n398), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n252), .B1(new_n388), .B2(new_n372), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n344), .A2(new_n253), .A3(new_n361), .A4(new_n369), .ZN(new_n407));
  NAND2_X1  g206(.A1(G227gat), .A2(G233gat), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n406), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(KEYINPUT32), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT33), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  XOR2_X1   g212(.A(G15gat), .B(G43gat), .Z(new_n414));
  XNOR2_X1  g213(.A(G71gat), .B(G99gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n411), .A2(new_n413), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n416), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n410), .B(KEYINPUT32), .C1(new_n412), .C2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n409), .B1(new_n406), .B2(new_n407), .ZN(new_n421));
  AND2_X1   g220(.A1(KEYINPUT72), .A2(KEYINPUT34), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n423), .B1(new_n421), .B2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n420), .A2(new_n426), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n235), .A2(KEYINPUT3), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n390), .B1(new_n428), .B2(KEYINPUT29), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT29), .B1(new_n383), .B2(new_n385), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n235), .B1(new_n430), .B2(KEYINPUT3), .ZN(new_n431));
  XNOR2_X1  g230(.A(G78gat), .B(G106gat), .ZN(new_n432));
  INV_X1    g231(.A(G50gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n432), .B(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n429), .A2(new_n431), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n435), .B1(new_n429), .B2(new_n431), .ZN(new_n438));
  NAND2_X1  g237(.A1(G228gat), .A2(G233gat), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n439), .B(G22gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n441));
  XOR2_X1   g240(.A(new_n440), .B(new_n441), .Z(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  OR3_X1    g242(.A1(new_n437), .A2(new_n438), .A3(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n443), .B1(new_n437), .B2(new_n438), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n425), .A2(new_n417), .A3(new_n419), .ZN(new_n447));
  AND3_X1   g246(.A1(new_n427), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n405), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(KEYINPUT35), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT84), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n404), .A2(new_n398), .ZN(new_n452));
  AOI211_X1 g251(.A(new_n208), .B(new_n210), .C1(new_n303), .C2(new_n304), .ZN(new_n453));
  AND4_X1   g252(.A1(new_n207), .A2(new_n303), .A3(new_n304), .A4(new_n206), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  XOR2_X1   g254(.A(KEYINPUT83), .B(KEYINPUT35), .Z(new_n456));
  NAND4_X1  g255(.A1(new_n427), .A2(new_n446), .A3(new_n447), .A4(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n451), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  AND4_X1   g257(.A1(new_n446), .A2(new_n427), .A3(new_n447), .A4(new_n456), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n459), .A2(new_n405), .A3(KEYINPUT84), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n446), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n303), .A2(new_n304), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n452), .B1(new_n463), .B2(new_n206), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n254), .A2(new_n255), .A3(new_n257), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(KEYINPUT39), .ZN(new_n466));
  OR2_X1    g265(.A1(new_n466), .A2(KEYINPUT82), .ZN(new_n467));
  AND2_X1   g266(.A1(new_n264), .A2(new_n274), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(new_n281), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n258), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n466), .A2(KEYINPUT82), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n467), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n257), .B1(new_n468), .B2(new_n281), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT39), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n206), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  AND3_X1   g274(.A1(new_n472), .A2(new_n475), .A3(KEYINPUT40), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT40), .B1(new_n472), .B2(new_n475), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n462), .B1(new_n464), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n403), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT37), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n402), .B1(new_n481), .B2(new_n397), .ZN(new_n482));
  AND2_X1   g281(.A1(new_n389), .A2(new_n392), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n481), .B1(new_n483), .B2(new_n386), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n375), .A2(new_n390), .ZN(new_n485));
  AOI21_X1  g284(.A(KEYINPUT38), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n480), .B1(new_n482), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n387), .A2(new_n393), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n399), .B1(new_n488), .B2(KEYINPUT37), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n481), .B1(new_n387), .B2(new_n393), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT38), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n294), .A2(new_n487), .A3(new_n491), .A4(new_n305), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n427), .A2(KEYINPUT36), .A3(new_n447), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT36), .ZN(new_n494));
  INV_X1    g293(.A(new_n447), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n425), .B1(new_n417), .B2(new_n419), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  AOI22_X1  g296(.A1(new_n479), .A2(new_n492), .B1(new_n493), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n455), .A2(new_n462), .ZN(new_n499));
  AOI22_X1  g298(.A1(new_n450), .A2(new_n461), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G15gat), .B(G22gat), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT16), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n501), .B1(new_n502), .B2(G1gat), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n503), .B1(G1gat), .B2(new_n501), .ZN(new_n504));
  XOR2_X1   g303(.A(new_n504), .B(G8gat), .Z(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(G43gat), .B(G50gat), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT15), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n512));
  NOR3_X1   g311(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n513));
  AND2_X1   g312(.A1(new_n513), .A2(KEYINPUT88), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n513), .A2(KEYINPUT88), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n512), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n508), .A2(new_n509), .ZN(new_n517));
  NAND2_X1  g316(.A1(G29gat), .A2(G36gat), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n511), .A2(new_n516), .A3(new_n517), .A4(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n513), .B(KEYINPUT85), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT86), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n521), .A2(new_n522), .A3(new_n512), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(new_n518), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n522), .B1(new_n521), .B2(new_n512), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n510), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT87), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT87), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n528), .B(new_n510), .C1(new_n524), .C2(new_n525), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n520), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n506), .B1(new_n530), .B2(KEYINPUT17), .ZN(new_n531));
  INV_X1    g330(.A(new_n529), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n521), .A2(new_n512), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT86), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n534), .A2(new_n518), .A3(new_n523), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n528), .B1(new_n535), .B2(new_n510), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n519), .B1(new_n532), .B2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT17), .ZN(new_n538));
  AOI21_X1  g337(.A(KEYINPUT89), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT89), .ZN(new_n540));
  NOR3_X1   g339(.A1(new_n530), .A2(new_n540), .A3(KEYINPUT17), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n531), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(G229gat), .A2(G233gat), .ZN(new_n543));
  XOR2_X1   g342(.A(new_n543), .B(KEYINPUT90), .Z(new_n544));
  NAND2_X1  g343(.A1(new_n537), .A2(new_n506), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n542), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT18), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n542), .A2(KEYINPUT18), .A3(new_n544), .A4(new_n545), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n530), .A2(new_n505), .ZN(new_n550));
  OR2_X1    g349(.A1(new_n550), .A2(KEYINPUT91), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(KEYINPUT91), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n551), .A2(new_n545), .A3(new_n552), .ZN(new_n553));
  XOR2_X1   g352(.A(new_n544), .B(KEYINPUT13), .Z(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n548), .A2(new_n549), .A3(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(G113gat), .B(G141gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(G197gat), .ZN(new_n558));
  XOR2_X1   g357(.A(KEYINPUT11), .B(G169gat), .Z(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  XOR2_X1   g359(.A(new_n560), .B(KEYINPUT12), .Z(new_n561));
  NAND2_X1  g360(.A1(new_n556), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n561), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n548), .A2(new_n563), .A3(new_n549), .A4(new_n555), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(G57gat), .ZN(new_n567));
  OAI21_X1  g366(.A(KEYINPUT92), .B1(new_n567), .B2(G64gat), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT92), .ZN(new_n569));
  INV_X1    g368(.A(G64gat), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n569), .A2(new_n570), .A3(G57gat), .ZN(new_n571));
  OAI211_X1 g370(.A(new_n568), .B(new_n571), .C1(G57gat), .C2(new_n570), .ZN(new_n572));
  NAND2_X1  g371(.A1(G71gat), .A2(G78gat), .ZN(new_n573));
  OR2_X1    g372(.A1(G71gat), .A2(G78gat), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT9), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(G57gat), .B(G64gat), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n573), .B(new_n574), .C1(new_n578), .C2(new_n575), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(KEYINPUT93), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT21), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(G231gat), .A2(G233gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(G127gat), .ZN(new_n586));
  XOR2_X1   g385(.A(G183gat), .B(G211gat), .Z(new_n587));
  XOR2_X1   g386(.A(new_n586), .B(new_n587), .Z(new_n588));
  OAI21_X1  g387(.A(new_n505), .B1(new_n581), .B2(new_n582), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT94), .ZN(new_n590));
  XNOR2_X1  g389(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(new_n230), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n590), .B(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n588), .B(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(G134gat), .B(G162gat), .Z(new_n595));
  AND2_X1   g394(.A1(G232gat), .A2(G233gat), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n596), .A2(KEYINPUT41), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n595), .B(new_n597), .ZN(new_n598));
  XOR2_X1   g397(.A(new_n598), .B(KEYINPUT97), .Z(new_n599));
  OAI211_X1 g398(.A(KEYINPUT17), .B(new_n519), .C1(new_n532), .C2(new_n536), .ZN(new_n600));
  NAND2_X1  g399(.A1(G85gat), .A2(G92gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT7), .ZN(new_n602));
  INV_X1    g401(.A(G99gat), .ZN(new_n603));
  INV_X1    g402(.A(G106gat), .ZN(new_n604));
  OAI21_X1  g403(.A(KEYINPUT8), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  XOR2_X1   g404(.A(KEYINPUT95), .B(G92gat), .Z(new_n606));
  OAI211_X1 g405(.A(new_n602), .B(new_n605), .C1(G85gat), .C2(new_n606), .ZN(new_n607));
  XOR2_X1   g406(.A(G99gat), .B(G106gat), .Z(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n600), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n540), .B1(new_n530), .B2(KEYINPUT17), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n537), .A2(KEYINPUT89), .A3(new_n538), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n609), .ZN(new_n614));
  AOI22_X1  g413(.A1(new_n537), .A2(new_n614), .B1(KEYINPUT41), .B2(new_n596), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(KEYINPUT96), .B1(new_n613), .B2(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n614), .B1(new_n530), .B2(KEYINPUT17), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n618), .B1(new_n539), .B2(new_n541), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT96), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n619), .A2(new_n620), .A3(new_n615), .ZN(new_n621));
  XNOR2_X1  g420(.A(G190gat), .B(G218gat), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  AND3_X1   g422(.A1(new_n617), .A2(new_n621), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n623), .B1(new_n617), .B2(new_n621), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n599), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NOR3_X1   g425(.A1(new_n613), .A2(KEYINPUT96), .A3(new_n616), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n620), .B1(new_n619), .B2(new_n615), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n622), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n598), .A2(KEYINPUT97), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n617), .A2(new_n621), .A3(new_n623), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n626), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n594), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(G230gat), .ZN(new_n635));
  INV_X1    g434(.A(G233gat), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n614), .A2(new_n580), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT93), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n580), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(new_n609), .ZN(new_n642));
  AOI21_X1  g441(.A(KEYINPUT10), .B1(new_n639), .B2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT10), .ZN(new_n644));
  NOR3_X1   g443(.A1(new_n581), .A2(new_n609), .A3(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n638), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n639), .A2(new_n642), .A3(new_n637), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g447(.A(G176gat), .B(G204gat), .Z(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT100), .ZN(new_n650));
  XNOR2_X1  g449(.A(G120gat), .B(G148gat), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n650), .B(new_n651), .Z(new_n652));
  XNOR2_X1  g451(.A(KEYINPUT98), .B(KEYINPUT99), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n648), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n654), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n646), .A2(new_n647), .A3(new_n656), .ZN(new_n657));
  AND3_X1   g456(.A1(new_n655), .A2(KEYINPUT101), .A3(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(KEYINPUT101), .B1(new_n655), .B2(new_n657), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR4_X1   g459(.A1(new_n500), .A2(new_n566), .A3(new_n634), .A4(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n453), .A2(new_n454), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(G1gat), .ZN(G1324gat));
  INV_X1    g463(.A(new_n452), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n666), .A2(KEYINPUT102), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(KEYINPUT102), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n667), .A2(G8gat), .A3(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT42), .ZN(new_n670));
  XNOR2_X1  g469(.A(KEYINPUT16), .B(G8gat), .ZN(new_n671));
  OR3_X1    g470(.A1(new_n666), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n671), .B1(new_n667), .B2(new_n668), .ZN(new_n673));
  OAI211_X1 g472(.A(new_n669), .B(new_n672), .C1(new_n673), .C2(KEYINPUT42), .ZN(G1325gat));
  NOR2_X1   g473(.A1(new_n495), .A2(new_n496), .ZN(new_n675));
  AOI21_X1  g474(.A(G15gat), .B1(new_n661), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n497), .A2(new_n493), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(G15gat), .ZN(new_n679));
  XOR2_X1   g478(.A(new_n679), .B(KEYINPUT103), .Z(new_n680));
  AOI21_X1  g479(.A(new_n676), .B1(new_n661), .B2(new_n680), .ZN(G1326gat));
  NAND2_X1  g480(.A1(new_n661), .A2(new_n462), .ZN(new_n682));
  XNOR2_X1  g481(.A(KEYINPUT43), .B(G22gat), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n682), .B(new_n683), .ZN(G1327gat));
  NOR3_X1   g483(.A1(new_n566), .A2(new_n594), .A3(new_n660), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n498), .A2(new_n499), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n455), .A2(new_n451), .A3(new_n457), .ZN(new_n687));
  AOI21_X1  g486(.A(KEYINPUT84), .B1(new_n459), .B2(new_n405), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n450), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n626), .A2(new_n632), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n685), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n662), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n692), .A2(G29gat), .A3(new_n693), .ZN(new_n694));
  XOR2_X1   g493(.A(new_n694), .B(KEYINPUT45), .Z(new_n695));
  OAI21_X1  g494(.A(KEYINPUT44), .B1(new_n500), .B2(new_n633), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT105), .ZN(new_n697));
  OAI21_X1  g496(.A(KEYINPUT104), .B1(new_n405), .B2(new_n446), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT104), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n455), .A2(new_n699), .A3(new_n462), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n463), .A2(new_n206), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n472), .A2(new_n475), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT40), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n472), .A2(KEYINPUT40), .A3(new_n475), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n665), .A2(new_n701), .A3(new_n704), .A4(new_n705), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n492), .A2(new_n706), .A3(new_n446), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n698), .A2(new_n700), .A3(new_n707), .A4(new_n677), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n689), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT44), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n626), .A2(new_n632), .A3(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n697), .B1(new_n709), .B2(new_n712), .ZN(new_n713));
  AOI211_X1 g512(.A(KEYINPUT105), .B(new_n711), .C1(new_n689), .C2(new_n708), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n696), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n715), .A2(KEYINPUT106), .A3(new_n685), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  AOI21_X1  g516(.A(KEYINPUT106), .B1(new_n715), .B2(new_n685), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n717), .A2(new_n693), .A3(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(G29gat), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n695), .B1(new_n719), .B2(new_n720), .ZN(G1328gat));
  NOR3_X1   g520(.A1(new_n692), .A2(G36gat), .A3(new_n452), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(KEYINPUT46), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n717), .A2(new_n452), .A3(new_n718), .ZN(new_n724));
  INV_X1    g523(.A(G36gat), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n723), .B1(new_n724), .B2(new_n725), .ZN(G1329gat));
  INV_X1    g525(.A(new_n675), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n692), .A2(G43gat), .A3(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT47), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n710), .B1(new_n690), .B2(new_n691), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n709), .A2(new_n712), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(KEYINPUT105), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n709), .A2(new_n697), .A3(new_n712), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n731), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n685), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n735), .A2(new_n677), .A3(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(G43gat), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n730), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT106), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n740), .B1(new_n735), .B2(new_n736), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n741), .A2(new_n678), .A3(new_n716), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n728), .B1(new_n742), .B2(G43gat), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n739), .B1(new_n743), .B2(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g543(.A1(new_n692), .A2(G50gat), .A3(new_n446), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT48), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n735), .A2(new_n446), .A3(new_n736), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n747), .B1(new_n748), .B2(new_n433), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n741), .A2(new_n462), .A3(new_n716), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n745), .B1(new_n750), .B2(G50gat), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n749), .B1(new_n751), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g551(.A(new_n634), .ZN(new_n753));
  AND4_X1   g552(.A1(new_n566), .A2(new_n753), .A3(new_n709), .A4(new_n660), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(new_n662), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g555(.A(new_n452), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(KEYINPUT107), .ZN(new_n759));
  NOR2_X1   g558(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n759), .B(new_n760), .ZN(G1333gat));
  XOR2_X1   g560(.A(new_n675), .B(KEYINPUT108), .Z(new_n762));
  AOI21_X1  g561(.A(G71gat), .B1(new_n754), .B2(new_n762), .ZN(new_n763));
  AND2_X1   g562(.A1(new_n678), .A2(G71gat), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n763), .B1(new_n754), .B2(new_n764), .ZN(new_n765));
  XOR2_X1   g564(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n766));
  XNOR2_X1  g565(.A(new_n765), .B(new_n766), .ZN(G1334gat));
  NAND2_X1  g566(.A1(new_n754), .A2(new_n462), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g568(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n770));
  XOR2_X1   g569(.A(KEYINPUT110), .B(KEYINPUT51), .Z(new_n771));
  NOR3_X1   g570(.A1(new_n594), .A2(new_n633), .A3(new_n565), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n709), .ZN(new_n773));
  MUX2_X1   g572(.A(new_n770), .B(new_n771), .S(new_n773), .Z(new_n774));
  INV_X1    g573(.A(new_n660), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(G85gat), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n776), .A2(new_n777), .A3(new_n662), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n594), .A2(new_n565), .A3(new_n775), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n735), .A2(new_n693), .A3(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n778), .B1(new_n777), .B2(new_n781), .ZN(G1336gat));
  NAND3_X1  g581(.A1(new_n715), .A2(new_n665), .A3(new_n779), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n606), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT52), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n775), .A2(G92gat), .A3(new_n452), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n784), .B(new_n785), .C1(new_n774), .C2(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n789), .ZN(new_n790));
  OAI211_X1 g589(.A(new_n772), .B(new_n709), .C1(KEYINPUT111), .C2(KEYINPUT51), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n787), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n784), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(KEYINPUT112), .B1(new_n794), .B2(KEYINPUT52), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n792), .B1(new_n783), .B2(new_n606), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT112), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n796), .A2(new_n797), .A3(new_n785), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n788), .B1(new_n795), .B2(new_n798), .ZN(G1337gat));
  NAND3_X1  g598(.A1(new_n776), .A2(new_n603), .A3(new_n675), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n735), .A2(new_n677), .A3(new_n780), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n800), .B1(new_n603), .B2(new_n801), .ZN(G1338gat));
  NOR2_X1   g601(.A1(new_n735), .A2(new_n780), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n604), .B1(new_n803), .B2(new_n462), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n775), .A2(G106gat), .A3(new_n446), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n806), .B1(new_n790), .B2(new_n791), .ZN(new_n807));
  OAI21_X1  g606(.A(KEYINPUT53), .B1(new_n804), .B2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n809), .B1(new_n774), .B2(new_n806), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n808), .B1(new_n804), .B2(new_n810), .ZN(G1339gat));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n812), .B(new_n638), .C1(new_n643), .C2(new_n645), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n813), .A2(new_n654), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n639), .A2(new_n642), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n645), .B1(new_n815), .B2(new_n644), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n637), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n817), .A2(KEYINPUT54), .A3(new_n646), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n814), .A2(new_n818), .A3(KEYINPUT55), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n819), .A2(new_n657), .ZN(new_n820));
  AOI21_X1  g619(.A(KEYINPUT55), .B1(new_n814), .B2(new_n818), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT113), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  AOI211_X1 g622(.A(KEYINPUT113), .B(KEYINPUT55), .C1(new_n814), .C2(new_n818), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n820), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n825), .B1(new_n562), .B2(new_n564), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n553), .A2(new_n554), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n544), .B1(new_n542), .B2(new_n545), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n560), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n564), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n830), .A2(new_n775), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n633), .B1(new_n826), .B2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(new_n825), .ZN(new_n833));
  INV_X1    g632(.A(new_n830), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n691), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(new_n594), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n634), .A2(new_n565), .A3(new_n660), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n841), .A2(new_n662), .A3(new_n448), .ZN(new_n842));
  OAI21_X1  g641(.A(KEYINPUT115), .B1(new_n842), .B2(new_n665), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n594), .B1(new_n832), .B2(new_n835), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n844), .A2(new_n839), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n845), .A2(new_n693), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT115), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n846), .A2(new_n847), .A3(new_n452), .A4(new_n448), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n843), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n849), .A2(new_n238), .A3(new_n565), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n693), .A2(new_n665), .A3(new_n727), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n841), .A2(new_n446), .A3(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(G113gat), .B1(new_n852), .B2(new_n566), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(KEYINPUT114), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT114), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n855), .B(G113gat), .C1(new_n852), .C2(new_n566), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n850), .A2(new_n857), .ZN(G1340gat));
  NAND3_X1  g657(.A1(new_n849), .A2(new_n236), .A3(new_n660), .ZN(new_n859));
  OAI21_X1  g658(.A(G120gat), .B1(new_n852), .B2(new_n775), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(G1341gat));
  NOR2_X1   g660(.A1(new_n845), .A2(new_n462), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n862), .A2(G127gat), .A3(new_n594), .A4(new_n851), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n863), .B(KEYINPUT116), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n842), .A2(new_n665), .ZN(new_n865));
  AOI21_X1  g664(.A(G127gat), .B1(new_n865), .B2(new_n594), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n864), .A2(new_n866), .ZN(G1342gat));
  NAND3_X1  g666(.A1(new_n691), .A2(new_n242), .A3(new_n452), .ZN(new_n868));
  OAI22_X1  g667(.A1(new_n842), .A2(new_n868), .B1(KEYINPUT118), .B2(KEYINPUT56), .ZN(new_n869));
  NAND2_X1  g668(.A1(KEYINPUT118), .A2(KEYINPUT56), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OAI211_X1 g670(.A(KEYINPUT118), .B(KEYINPUT56), .C1(new_n842), .C2(new_n868), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n862), .A2(new_n691), .A3(new_n851), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n873), .A2(KEYINPUT117), .A3(G134gat), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(KEYINPUT117), .B1(new_n873), .B2(G134gat), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n871), .B(new_n872), .C1(new_n875), .C2(new_n876), .ZN(G1343gat));
  XNOR2_X1  g676(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n819), .A2(new_n657), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n879), .A2(new_n821), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n881), .B1(new_n562), .B2(new_n564), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n633), .B1(new_n882), .B2(new_n831), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n594), .B1(new_n883), .B2(new_n835), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n462), .B1(new_n884), .B2(new_n839), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(KEYINPUT57), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT57), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n887), .B(new_n462), .C1(new_n844), .C2(new_n839), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n678), .A2(new_n693), .A3(new_n665), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n886), .A2(new_n565), .A3(new_n888), .A4(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(new_n268), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n677), .A2(new_n462), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n893), .A2(new_n665), .ZN(new_n894));
  OAI211_X1 g693(.A(new_n662), .B(new_n894), .C1(new_n844), .C2(new_n839), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n565), .A2(new_n219), .ZN(new_n896));
  XOR2_X1   g695(.A(new_n896), .B(KEYINPUT119), .Z(new_n897));
  NOR2_X1   g696(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n878), .B1(new_n892), .B2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(new_n878), .ZN(new_n901));
  AOI211_X1 g700(.A(new_n898), .B(new_n901), .C1(new_n890), .C2(new_n891), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n900), .A2(new_n902), .ZN(G1344gat));
  OR3_X1    g702(.A1(new_n895), .A2(G148gat), .A3(new_n775), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT59), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(G148gat), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n886), .A2(new_n888), .A3(new_n889), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n906), .B1(new_n908), .B2(new_n660), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n887), .B(new_n462), .C1(new_n884), .C2(new_n839), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n889), .A2(new_n660), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n446), .B1(new_n838), .B2(new_n840), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n910), .B(new_n911), .C1(new_n912), .C2(new_n887), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n905), .B1(new_n913), .B2(G148gat), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n904), .B1(new_n909), .B2(new_n914), .ZN(G1345gat));
  OAI21_X1  g714(.A(G155gat), .B1(new_n907), .B2(new_n837), .ZN(new_n916));
  INV_X1    g715(.A(new_n895), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n917), .A2(new_n230), .A3(new_n594), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n916), .A2(new_n918), .ZN(G1346gat));
  XOR2_X1   g718(.A(KEYINPUT75), .B(G162gat), .Z(new_n920));
  NAND3_X1  g719(.A1(new_n917), .A2(new_n691), .A3(new_n920), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n907), .A2(new_n633), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n921), .B1(new_n922), .B2(new_n920), .ZN(G1347gat));
  NOR2_X1   g722(.A1(new_n662), .A2(new_n452), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n762), .A2(new_n924), .ZN(new_n925));
  OAI211_X1 g724(.A(new_n446), .B(new_n925), .C1(new_n844), .C2(new_n839), .ZN(new_n926));
  OAI21_X1  g725(.A(G169gat), .B1(new_n926), .B2(new_n566), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n448), .A2(new_n665), .ZN(new_n928));
  OAI211_X1 g727(.A(new_n693), .B(new_n928), .C1(new_n844), .C2(new_n839), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n565), .A2(new_n318), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n927), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n931), .B(KEYINPUT121), .ZN(G1348gat));
  NOR3_X1   g731(.A1(new_n926), .A2(new_n317), .A3(new_n775), .ZN(new_n933));
  INV_X1    g732(.A(new_n929), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(new_n660), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n933), .B1(new_n935), .B2(new_n329), .ZN(G1349gat));
  NAND2_X1  g735(.A1(new_n594), .A2(new_n346), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n934), .A2(KEYINPUT122), .A3(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT122), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n940), .B1(new_n929), .B2(new_n937), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g741(.A(G183gat), .B1(new_n926), .B2(new_n837), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(KEYINPUT60), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT60), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n942), .A2(new_n946), .A3(new_n943), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n945), .A2(new_n947), .ZN(G1350gat));
  NAND3_X1  g747(.A1(new_n934), .A2(new_n325), .A3(new_n691), .ZN(new_n949));
  OAI21_X1  g748(.A(G190gat), .B1(new_n926), .B2(new_n633), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(KEYINPUT123), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT61), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT123), .ZN(new_n953));
  OAI211_X1 g752(.A(new_n953), .B(G190gat), .C1(new_n926), .C2(new_n633), .ZN(new_n954));
  AND3_X1   g753(.A1(new_n951), .A2(new_n952), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n952), .B1(new_n951), .B2(new_n954), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n949), .B1(new_n955), .B2(new_n956), .ZN(G1351gat));
  NOR2_X1   g756(.A1(new_n893), .A2(new_n452), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n841), .A2(new_n693), .A3(new_n958), .ZN(new_n959));
  OR3_X1    g758(.A1(new_n959), .A2(G197gat), .A3(new_n566), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n924), .A2(new_n677), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n961), .B(KEYINPUT124), .ZN(new_n962));
  OAI211_X1 g761(.A(new_n910), .B(new_n962), .C1(new_n912), .C2(new_n887), .ZN(new_n963));
  OAI21_X1  g762(.A(KEYINPUT125), .B1(new_n963), .B2(new_n566), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(G197gat), .ZN(new_n965));
  NOR3_X1   g764(.A1(new_n963), .A2(KEYINPUT125), .A3(new_n566), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n960), .B1(new_n965), .B2(new_n966), .ZN(G1352gat));
  OAI21_X1  g766(.A(G204gat), .B1(new_n963), .B2(new_n775), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n775), .A2(G204gat), .ZN(new_n969));
  INV_X1    g768(.A(new_n969), .ZN(new_n970));
  OR3_X1    g769(.A1(new_n959), .A2(KEYINPUT62), .A3(new_n970), .ZN(new_n971));
  OAI21_X1  g770(.A(KEYINPUT62), .B1(new_n959), .B2(new_n970), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n968), .A2(new_n971), .A3(new_n972), .ZN(G1353gat));
  INV_X1    g772(.A(KEYINPUT126), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n837), .A2(new_n961), .ZN(new_n975));
  OAI211_X1 g774(.A(new_n910), .B(new_n975), .C1(new_n912), .C2(new_n887), .ZN(new_n976));
  AND4_X1   g775(.A1(new_n974), .A2(new_n976), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n977));
  INV_X1    g776(.A(G211gat), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT63), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n978), .B1(KEYINPUT126), .B2(new_n979), .ZN(new_n980));
  AOI22_X1  g779(.A1(new_n976), .A2(new_n980), .B1(new_n974), .B2(KEYINPUT63), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n594), .A2(new_n978), .ZN(new_n982));
  OAI22_X1  g781(.A1(new_n977), .A2(new_n981), .B1(new_n959), .B2(new_n982), .ZN(G1354gat));
  NOR2_X1   g782(.A1(new_n959), .A2(new_n633), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n984), .A2(G218gat), .ZN(new_n985));
  INV_X1    g784(.A(new_n963), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n691), .A2(G218gat), .ZN(new_n987));
  XOR2_X1   g786(.A(new_n987), .B(KEYINPUT127), .Z(new_n988));
  AOI21_X1  g787(.A(new_n985), .B1(new_n986), .B2(new_n988), .ZN(G1355gat));
endmodule


