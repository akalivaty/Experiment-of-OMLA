

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U552 ( .A(n660), .ZN(n633) );
  XOR2_X1 U553 ( .A(KEYINPUT72), .B(n619), .Z(n519) );
  OR2_X1 U554 ( .A1(n707), .A2(n706), .ZN(n520) );
  AND2_X1 U555 ( .A1(n703), .A2(n702), .ZN(n521) );
  XNOR2_X1 U556 ( .A(KEYINPUT32), .B(KEYINPUT100), .ZN(n670) );
  XNOR2_X1 U557 ( .A(n671), .B(n670), .ZN(n696) );
  XNOR2_X1 U558 ( .A(n623), .B(KEYINPUT15), .ZN(n841) );
  NOR2_X1 U559 ( .A1(G651), .A2(n575), .ZN(n793) );
  NOR2_X1 U560 ( .A1(n537), .A2(n536), .ZN(G160) );
  NOR2_X1 U561 ( .A1(G2105), .A2(G2104), .ZN(n522) );
  XOR2_X1 U562 ( .A(KEYINPUT17), .B(n522), .Z(n890) );
  NAND2_X1 U563 ( .A1(G138), .A2(n890), .ZN(n525) );
  INV_X1 U564 ( .A(G2105), .ZN(n526) );
  NAND2_X1 U565 ( .A1(n526), .A2(G2104), .ZN(n523) );
  XNOR2_X2 U566 ( .A(n523), .B(KEYINPUT65), .ZN(n891) );
  NAND2_X1 U567 ( .A1(G102), .A2(n891), .ZN(n524) );
  NAND2_X1 U568 ( .A1(n525), .A2(n524), .ZN(n530) );
  NOR2_X1 U569 ( .A1(G2104), .A2(n526), .ZN(n894) );
  NAND2_X1 U570 ( .A1(G126), .A2(n894), .ZN(n528) );
  AND2_X1 U571 ( .A1(G2105), .A2(G2104), .ZN(n895) );
  NAND2_X1 U572 ( .A1(G114), .A2(n895), .ZN(n527) );
  NAND2_X1 U573 ( .A1(n528), .A2(n527), .ZN(n529) );
  NOR2_X1 U574 ( .A1(n530), .A2(n529), .ZN(G164) );
  NAND2_X1 U575 ( .A1(G125), .A2(n894), .ZN(n532) );
  NAND2_X1 U576 ( .A1(G113), .A2(n895), .ZN(n531) );
  NAND2_X1 U577 ( .A1(n532), .A2(n531), .ZN(n537) );
  NAND2_X1 U578 ( .A1(G101), .A2(n891), .ZN(n533) );
  XOR2_X1 U579 ( .A(KEYINPUT23), .B(n533), .Z(n535) );
  NAND2_X1 U580 ( .A1(n890), .A2(G137), .ZN(n534) );
  NAND2_X1 U581 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U582 ( .A(G651), .B(KEYINPUT66), .Z(n541) );
  NOR2_X1 U583 ( .A1(G543), .A2(n541), .ZN(n538) );
  XOR2_X2 U584 ( .A(KEYINPUT1), .B(n538), .Z(n796) );
  NAND2_X1 U585 ( .A1(G64), .A2(n796), .ZN(n540) );
  XOR2_X1 U586 ( .A(KEYINPUT0), .B(G543), .Z(n575) );
  NAND2_X1 U587 ( .A1(G52), .A2(n793), .ZN(n539) );
  NAND2_X1 U588 ( .A1(n540), .A2(n539), .ZN(n548) );
  OR2_X1 U589 ( .A1(n575), .A2(n541), .ZN(n542) );
  XNOR2_X1 U590 ( .A(n542), .B(KEYINPUT67), .ZN(n792) );
  NAND2_X1 U591 ( .A1(n792), .A2(G77), .ZN(n545) );
  NOR2_X1 U592 ( .A1(G543), .A2(G651), .ZN(n543) );
  XNOR2_X1 U593 ( .A(n543), .B(KEYINPUT64), .ZN(n797) );
  NAND2_X1 U594 ( .A1(G90), .A2(n797), .ZN(n544) );
  NAND2_X1 U595 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U596 ( .A(KEYINPUT9), .B(n546), .Z(n547) );
  NOR2_X1 U597 ( .A1(n548), .A2(n547), .ZN(G171) );
  NAND2_X1 U598 ( .A1(G78), .A2(n792), .ZN(n550) );
  NAND2_X1 U599 ( .A1(G53), .A2(n793), .ZN(n549) );
  NAND2_X1 U600 ( .A1(n550), .A2(n549), .ZN(n554) );
  NAND2_X1 U601 ( .A1(n796), .A2(G65), .ZN(n552) );
  NAND2_X1 U602 ( .A1(G91), .A2(n797), .ZN(n551) );
  NAND2_X1 U603 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X1 U604 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U605 ( .A(n555), .B(KEYINPUT69), .ZN(G299) );
  NAND2_X1 U606 ( .A1(G89), .A2(n797), .ZN(n556) );
  XNOR2_X1 U607 ( .A(n556), .B(KEYINPUT4), .ZN(n558) );
  NAND2_X1 U608 ( .A1(G76), .A2(n792), .ZN(n557) );
  NAND2_X1 U609 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U610 ( .A(KEYINPUT5), .B(n559), .ZN(n565) );
  NAND2_X1 U611 ( .A1(n793), .A2(G51), .ZN(n560) );
  XOR2_X1 U612 ( .A(KEYINPUT73), .B(n560), .Z(n562) );
  NAND2_X1 U613 ( .A1(n796), .A2(G63), .ZN(n561) );
  NAND2_X1 U614 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U615 ( .A(KEYINPUT6), .B(n563), .Z(n564) );
  NAND2_X1 U616 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U617 ( .A(KEYINPUT7), .B(n566), .ZN(G168) );
  NAND2_X1 U618 ( .A1(n796), .A2(G62), .ZN(n567) );
  XNOR2_X1 U619 ( .A(n567), .B(KEYINPUT80), .ZN(n569) );
  NAND2_X1 U620 ( .A1(G50), .A2(n793), .ZN(n568) );
  NAND2_X1 U621 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U622 ( .A(KEYINPUT81), .B(n570), .ZN(n574) );
  NAND2_X1 U623 ( .A1(n797), .A2(G88), .ZN(n572) );
  NAND2_X1 U624 ( .A1(n792), .A2(G75), .ZN(n571) );
  AND2_X1 U625 ( .A1(n572), .A2(n571), .ZN(n573) );
  NAND2_X1 U626 ( .A1(n574), .A2(n573), .ZN(G303) );
  XOR2_X1 U627 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U628 ( .A1(G87), .A2(n575), .ZN(n577) );
  NAND2_X1 U629 ( .A1(G74), .A2(G651), .ZN(n576) );
  NAND2_X1 U630 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U631 ( .A1(n796), .A2(n578), .ZN(n580) );
  NAND2_X1 U632 ( .A1(n793), .A2(G49), .ZN(n579) );
  NAND2_X1 U633 ( .A1(n580), .A2(n579), .ZN(G288) );
  NAND2_X1 U634 ( .A1(G73), .A2(n792), .ZN(n581) );
  XNOR2_X1 U635 ( .A(n581), .B(KEYINPUT2), .ZN(n582) );
  XNOR2_X1 U636 ( .A(n582), .B(KEYINPUT78), .ZN(n584) );
  NAND2_X1 U637 ( .A1(G86), .A2(n797), .ZN(n583) );
  NAND2_X1 U638 ( .A1(n584), .A2(n583), .ZN(n587) );
  NAND2_X1 U639 ( .A1(G48), .A2(n793), .ZN(n585) );
  XNOR2_X1 U640 ( .A(KEYINPUT79), .B(n585), .ZN(n586) );
  NOR2_X1 U641 ( .A1(n587), .A2(n586), .ZN(n590) );
  NAND2_X1 U642 ( .A1(G61), .A2(n796), .ZN(n588) );
  XOR2_X1 U643 ( .A(KEYINPUT77), .B(n588), .Z(n589) );
  NAND2_X1 U644 ( .A1(n590), .A2(n589), .ZN(G305) );
  NAND2_X1 U645 ( .A1(n792), .A2(G72), .ZN(n592) );
  NAND2_X1 U646 ( .A1(G85), .A2(n797), .ZN(n591) );
  NAND2_X1 U647 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U648 ( .A(KEYINPUT68), .B(n593), .Z(n597) );
  NAND2_X1 U649 ( .A1(G60), .A2(n796), .ZN(n595) );
  NAND2_X1 U650 ( .A1(G47), .A2(n793), .ZN(n594) );
  AND2_X1 U651 ( .A1(n595), .A2(n594), .ZN(n596) );
  NAND2_X1 U652 ( .A1(n597), .A2(n596), .ZN(G290) );
  NOR2_X1 U653 ( .A1(G164), .A2(G1384), .ZN(n720) );
  NAND2_X1 U654 ( .A1(G160), .A2(G40), .ZN(n719) );
  INV_X1 U655 ( .A(n719), .ZN(n598) );
  NAND2_X1 U656 ( .A1(n720), .A2(n598), .ZN(n660) );
  OR2_X1 U657 ( .A1(n633), .A2(G1961), .ZN(n600) );
  XNOR2_X1 U658 ( .A(KEYINPUT25), .B(G2078), .ZN(n923) );
  NAND2_X1 U659 ( .A1(n633), .A2(n923), .ZN(n599) );
  NAND2_X1 U660 ( .A1(n600), .A2(n599), .ZN(n654) );
  NAND2_X1 U661 ( .A1(n654), .A2(G171), .ZN(n647) );
  NOR2_X1 U662 ( .A1(n633), .A2(G1348), .ZN(n602) );
  NOR2_X1 U663 ( .A1(G2067), .A2(n660), .ZN(n601) );
  NOR2_X1 U664 ( .A1(n602), .A2(n601), .ZN(n626) );
  AND2_X1 U665 ( .A1(n633), .A2(G1996), .ZN(n603) );
  XOR2_X1 U666 ( .A(n603), .B(KEYINPUT26), .Z(n605) );
  NAND2_X1 U667 ( .A1(n660), .A2(G1341), .ZN(n604) );
  AND2_X1 U668 ( .A1(n605), .A2(n604), .ZN(n628) );
  NAND2_X1 U669 ( .A1(G56), .A2(n796), .ZN(n606) );
  XOR2_X1 U670 ( .A(KEYINPUT14), .B(n606), .Z(n614) );
  XOR2_X1 U671 ( .A(KEYINPUT12), .B(KEYINPUT71), .Z(n608) );
  NAND2_X1 U672 ( .A1(G81), .A2(n797), .ZN(n607) );
  XNOR2_X1 U673 ( .A(n608), .B(n607), .ZN(n609) );
  XNOR2_X1 U674 ( .A(KEYINPUT70), .B(n609), .ZN(n611) );
  NAND2_X1 U675 ( .A1(n792), .A2(G68), .ZN(n610) );
  NAND2_X1 U676 ( .A1(n611), .A2(n610), .ZN(n612) );
  XOR2_X1 U677 ( .A(KEYINPUT13), .B(n612), .Z(n613) );
  NOR2_X1 U678 ( .A1(n614), .A2(n613), .ZN(n616) );
  NAND2_X1 U679 ( .A1(n793), .A2(G43), .ZN(n615) );
  NAND2_X1 U680 ( .A1(n616), .A2(n615), .ZN(n936) );
  INV_X1 U681 ( .A(n936), .ZN(n629) );
  NAND2_X1 U682 ( .A1(G54), .A2(n793), .ZN(n622) );
  NAND2_X1 U683 ( .A1(n792), .A2(G79), .ZN(n618) );
  NAND2_X1 U684 ( .A1(G92), .A2(n797), .ZN(n617) );
  NAND2_X1 U685 ( .A1(n618), .A2(n617), .ZN(n620) );
  NAND2_X1 U686 ( .A1(n796), .A2(G66), .ZN(n619) );
  NOR2_X1 U687 ( .A1(n620), .A2(n519), .ZN(n621) );
  NAND2_X1 U688 ( .A1(n622), .A2(n621), .ZN(n623) );
  AND2_X1 U689 ( .A1(n629), .A2(n841), .ZN(n624) );
  NAND2_X1 U690 ( .A1(n628), .A2(n624), .ZN(n625) );
  NAND2_X1 U691 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X1 U692 ( .A(n627), .B(KEYINPUT96), .ZN(n632) );
  AND2_X1 U693 ( .A1(n629), .A2(n628), .ZN(n630) );
  OR2_X1 U694 ( .A1(n841), .A2(n630), .ZN(n631) );
  NAND2_X1 U695 ( .A1(n632), .A2(n631), .ZN(n639) );
  INV_X1 U696 ( .A(G299), .ZN(n953) );
  NAND2_X1 U697 ( .A1(n633), .A2(G2072), .ZN(n634) );
  XNOR2_X1 U698 ( .A(KEYINPUT27), .B(n634), .ZN(n637) );
  NAND2_X1 U699 ( .A1(G1956), .A2(n660), .ZN(n635) );
  XOR2_X1 U700 ( .A(KEYINPUT94), .B(n635), .Z(n636) );
  NOR2_X1 U701 ( .A1(n637), .A2(n636), .ZN(n640) );
  NAND2_X1 U702 ( .A1(n953), .A2(n640), .ZN(n638) );
  NAND2_X1 U703 ( .A1(n639), .A2(n638), .ZN(n644) );
  NOR2_X1 U704 ( .A1(n953), .A2(n640), .ZN(n642) );
  XNOR2_X1 U705 ( .A(KEYINPUT95), .B(KEYINPUT28), .ZN(n641) );
  XNOR2_X1 U706 ( .A(n642), .B(n641), .ZN(n643) );
  NAND2_X1 U707 ( .A1(n644), .A2(n643), .ZN(n645) );
  XOR2_X1 U708 ( .A(KEYINPUT29), .B(n645), .Z(n646) );
  NAND2_X1 U709 ( .A1(n647), .A2(n646), .ZN(n673) );
  NOR2_X1 U710 ( .A1(G2084), .A2(n660), .ZN(n674) );
  INV_X1 U711 ( .A(G8), .ZN(n648) );
  NOR2_X1 U712 ( .A1(n648), .A2(G1966), .ZN(n649) );
  AND2_X1 U713 ( .A1(n649), .A2(n660), .ZN(n650) );
  XNOR2_X1 U714 ( .A(n650), .B(KEYINPUT93), .ZN(n676) );
  NAND2_X1 U715 ( .A1(G8), .A2(n676), .ZN(n651) );
  NOR2_X1 U716 ( .A1(n674), .A2(n651), .ZN(n652) );
  XOR2_X1 U717 ( .A(KEYINPUT30), .B(n652), .Z(n653) );
  NOR2_X1 U718 ( .A1(G168), .A2(n653), .ZN(n656) );
  NOR2_X1 U719 ( .A1(G171), .A2(n654), .ZN(n655) );
  NOR2_X1 U720 ( .A1(n656), .A2(n655), .ZN(n657) );
  XOR2_X1 U721 ( .A(n657), .B(KEYINPUT31), .Z(n672) );
  NOR2_X1 U722 ( .A1(G2090), .A2(n660), .ZN(n658) );
  XOR2_X1 U723 ( .A(KEYINPUT98), .B(n658), .Z(n659) );
  NAND2_X1 U724 ( .A1(n659), .A2(G303), .ZN(n662) );
  NAND2_X1 U725 ( .A1(G8), .A2(n660), .ZN(n707) );
  NOR2_X1 U726 ( .A1(G1971), .A2(n707), .ZN(n661) );
  NOR2_X1 U727 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U728 ( .A(n663), .B(KEYINPUT99), .ZN(n665) );
  AND2_X1 U729 ( .A1(n672), .A2(n665), .ZN(n664) );
  NAND2_X1 U730 ( .A1(n673), .A2(n664), .ZN(n668) );
  INV_X1 U731 ( .A(n665), .ZN(n666) );
  OR2_X1 U732 ( .A1(n666), .A2(G286), .ZN(n667) );
  AND2_X1 U733 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U734 ( .A1(n669), .A2(G8), .ZN(n671) );
  AND2_X1 U735 ( .A1(n673), .A2(n672), .ZN(n678) );
  NAND2_X1 U736 ( .A1(G8), .A2(n674), .ZN(n675) );
  NAND2_X1 U737 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U738 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U739 ( .A(KEYINPUT97), .B(n679), .ZN(n697) );
  NOR2_X1 U740 ( .A1(G1976), .A2(G288), .ZN(n688) );
  INV_X1 U741 ( .A(n707), .ZN(n680) );
  NAND2_X1 U742 ( .A1(n688), .A2(n680), .ZN(n681) );
  NAND2_X1 U743 ( .A1(n681), .A2(KEYINPUT33), .ZN(n689) );
  INV_X1 U744 ( .A(n689), .ZN(n684) );
  NOR2_X1 U745 ( .A1(n707), .A2(KEYINPUT33), .ZN(n682) );
  NAND2_X1 U746 ( .A1(G1976), .A2(G288), .ZN(n940) );
  AND2_X1 U747 ( .A1(n682), .A2(n940), .ZN(n683) );
  OR2_X1 U748 ( .A1(n684), .A2(n683), .ZN(n686) );
  AND2_X1 U749 ( .A1(n697), .A2(n686), .ZN(n685) );
  NAND2_X1 U750 ( .A1(n696), .A2(n685), .ZN(n693) );
  INV_X1 U751 ( .A(n686), .ZN(n691) );
  NOR2_X1 U752 ( .A1(G1971), .A2(G303), .ZN(n687) );
  NOR2_X1 U753 ( .A1(n688), .A2(n687), .ZN(n941) );
  AND2_X1 U754 ( .A1(n941), .A2(n689), .ZN(n690) );
  OR2_X1 U755 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U756 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U757 ( .A(KEYINPUT101), .B(n694), .Z(n695) );
  XOR2_X1 U758 ( .A(G1981), .B(G305), .Z(n937) );
  NAND2_X1 U759 ( .A1(n695), .A2(n937), .ZN(n703) );
  NAND2_X1 U760 ( .A1(n697), .A2(n696), .ZN(n700) );
  NOR2_X1 U761 ( .A1(G2090), .A2(G303), .ZN(n698) );
  NAND2_X1 U762 ( .A1(G8), .A2(n698), .ZN(n699) );
  NAND2_X1 U763 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U764 ( .A1(n701), .A2(n707), .ZN(n702) );
  NOR2_X1 U765 ( .A1(G1981), .A2(G305), .ZN(n704) );
  XOR2_X1 U766 ( .A(n704), .B(KEYINPUT24), .Z(n705) );
  XNOR2_X1 U767 ( .A(KEYINPUT92), .B(n705), .ZN(n706) );
  NAND2_X1 U768 ( .A1(n521), .A2(n520), .ZN(n743) );
  XNOR2_X1 U769 ( .A(G2067), .B(KEYINPUT37), .ZN(n744) );
  NAND2_X1 U770 ( .A1(n891), .A2(G104), .ZN(n708) );
  XOR2_X1 U771 ( .A(KEYINPUT87), .B(n708), .Z(n710) );
  NAND2_X1 U772 ( .A1(n890), .A2(G140), .ZN(n709) );
  NAND2_X1 U773 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U774 ( .A(KEYINPUT34), .B(n711), .ZN(n717) );
  NAND2_X1 U775 ( .A1(n894), .A2(G128), .ZN(n712) );
  XNOR2_X1 U776 ( .A(n712), .B(KEYINPUT88), .ZN(n714) );
  NAND2_X1 U777 ( .A1(G116), .A2(n895), .ZN(n713) );
  NAND2_X1 U778 ( .A1(n714), .A2(n713), .ZN(n715) );
  XOR2_X1 U779 ( .A(KEYINPUT35), .B(n715), .Z(n716) );
  NOR2_X1 U780 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U781 ( .A(KEYINPUT36), .B(n718), .ZN(n904) );
  NOR2_X1 U782 ( .A1(n744), .A2(n904), .ZN(n1017) );
  NOR2_X1 U783 ( .A1(n720), .A2(n719), .ZN(n753) );
  NAND2_X1 U784 ( .A1(n1017), .A2(n753), .ZN(n721) );
  XOR2_X1 U785 ( .A(KEYINPUT89), .B(n721), .Z(n750) );
  NAND2_X1 U786 ( .A1(G129), .A2(n894), .ZN(n723) );
  NAND2_X1 U787 ( .A1(G117), .A2(n895), .ZN(n722) );
  NAND2_X1 U788 ( .A1(n723), .A2(n722), .ZN(n726) );
  NAND2_X1 U789 ( .A1(n891), .A2(G105), .ZN(n724) );
  XOR2_X1 U790 ( .A(KEYINPUT38), .B(n724), .Z(n725) );
  NOR2_X1 U791 ( .A1(n726), .A2(n725), .ZN(n728) );
  NAND2_X1 U792 ( .A1(n890), .A2(G141), .ZN(n727) );
  NAND2_X1 U793 ( .A1(n728), .A2(n727), .ZN(n875) );
  NAND2_X1 U794 ( .A1(G1996), .A2(n875), .ZN(n729) );
  XNOR2_X1 U795 ( .A(n729), .B(KEYINPUT90), .ZN(n737) );
  NAND2_X1 U796 ( .A1(G131), .A2(n890), .ZN(n731) );
  NAND2_X1 U797 ( .A1(G95), .A2(n891), .ZN(n730) );
  NAND2_X1 U798 ( .A1(n731), .A2(n730), .ZN(n735) );
  NAND2_X1 U799 ( .A1(G119), .A2(n894), .ZN(n733) );
  NAND2_X1 U800 ( .A1(G107), .A2(n895), .ZN(n732) );
  NAND2_X1 U801 ( .A1(n733), .A2(n732), .ZN(n734) );
  OR2_X1 U802 ( .A1(n735), .A2(n734), .ZN(n876) );
  NAND2_X1 U803 ( .A1(G1991), .A2(n876), .ZN(n736) );
  NAND2_X1 U804 ( .A1(n737), .A2(n736), .ZN(n1006) );
  NAND2_X1 U805 ( .A1(n753), .A2(n1006), .ZN(n738) );
  NAND2_X1 U806 ( .A1(n750), .A2(n738), .ZN(n739) );
  XOR2_X1 U807 ( .A(KEYINPUT91), .B(n739), .Z(n741) );
  XNOR2_X1 U808 ( .A(G1986), .B(G290), .ZN(n955) );
  AND2_X1 U809 ( .A1(n955), .A2(n753), .ZN(n740) );
  NOR2_X1 U810 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U811 ( .A1(n743), .A2(n742), .ZN(n756) );
  NAND2_X1 U812 ( .A1(n744), .A2(n904), .ZN(n1014) );
  NOR2_X1 U813 ( .A1(G1996), .A2(n875), .ZN(n1010) );
  NOR2_X1 U814 ( .A1(G1986), .A2(G290), .ZN(n745) );
  NOR2_X1 U815 ( .A1(G1991), .A2(n876), .ZN(n997) );
  NOR2_X1 U816 ( .A1(n745), .A2(n997), .ZN(n746) );
  NOR2_X1 U817 ( .A1(n1006), .A2(n746), .ZN(n747) );
  NOR2_X1 U818 ( .A1(n1010), .A2(n747), .ZN(n748) );
  XNOR2_X1 U819 ( .A(KEYINPUT102), .B(n748), .ZN(n749) );
  XNOR2_X1 U820 ( .A(n749), .B(KEYINPUT39), .ZN(n751) );
  NAND2_X1 U821 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U822 ( .A1(n1014), .A2(n752), .ZN(n754) );
  NAND2_X1 U823 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U824 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U825 ( .A(n757), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U826 ( .A(KEYINPUT103), .B(G2435), .Z(n759) );
  XNOR2_X1 U827 ( .A(G2430), .B(G2438), .ZN(n758) );
  XNOR2_X1 U828 ( .A(n759), .B(n758), .ZN(n766) );
  XOR2_X1 U829 ( .A(G2446), .B(G2454), .Z(n761) );
  XNOR2_X1 U830 ( .A(G2451), .B(G2443), .ZN(n760) );
  XNOR2_X1 U831 ( .A(n761), .B(n760), .ZN(n762) );
  XOR2_X1 U832 ( .A(n762), .B(G2427), .Z(n764) );
  XNOR2_X1 U833 ( .A(G1341), .B(G1348), .ZN(n763) );
  XNOR2_X1 U834 ( .A(n764), .B(n763), .ZN(n765) );
  XNOR2_X1 U835 ( .A(n766), .B(n765), .ZN(n767) );
  AND2_X1 U836 ( .A1(n767), .A2(G14), .ZN(G401) );
  AND2_X1 U837 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U838 ( .A(G108), .ZN(G238) );
  INV_X1 U839 ( .A(G120), .ZN(G236) );
  INV_X1 U840 ( .A(G69), .ZN(G235) );
  INV_X1 U841 ( .A(G132), .ZN(G219) );
  INV_X1 U842 ( .A(G82), .ZN(G220) );
  NAND2_X1 U843 ( .A1(G7), .A2(G661), .ZN(n768) );
  XNOR2_X1 U844 ( .A(n768), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U845 ( .A(G223), .ZN(n828) );
  NAND2_X1 U846 ( .A1(n828), .A2(G567), .ZN(n769) );
  XOR2_X1 U847 ( .A(KEYINPUT11), .B(n769), .Z(G234) );
  INV_X1 U848 ( .A(G860), .ZN(n834) );
  OR2_X1 U849 ( .A1(n936), .A2(n834), .ZN(G153) );
  INV_X1 U850 ( .A(G171), .ZN(G301) );
  NAND2_X1 U851 ( .A1(G868), .A2(G301), .ZN(n771) );
  INV_X1 U852 ( .A(n841), .ZN(n947) );
  INV_X1 U853 ( .A(G868), .ZN(n808) );
  NAND2_X1 U854 ( .A1(n947), .A2(n808), .ZN(n770) );
  NAND2_X1 U855 ( .A1(n771), .A2(n770), .ZN(G284) );
  NAND2_X1 U856 ( .A1(G286), .A2(G868), .ZN(n773) );
  NAND2_X1 U857 ( .A1(G299), .A2(n808), .ZN(n772) );
  NAND2_X1 U858 ( .A1(n773), .A2(n772), .ZN(G297) );
  NAND2_X1 U859 ( .A1(n834), .A2(G559), .ZN(n774) );
  NAND2_X1 U860 ( .A1(n774), .A2(n841), .ZN(n775) );
  XNOR2_X1 U861 ( .A(n775), .B(KEYINPUT74), .ZN(n776) );
  XNOR2_X1 U862 ( .A(KEYINPUT16), .B(n776), .ZN(G148) );
  NOR2_X1 U863 ( .A1(n947), .A2(n808), .ZN(n777) );
  XNOR2_X1 U864 ( .A(n777), .B(KEYINPUT75), .ZN(n778) );
  NOR2_X1 U865 ( .A1(G559), .A2(n778), .ZN(n780) );
  NOR2_X1 U866 ( .A1(G868), .A2(n936), .ZN(n779) );
  NOR2_X1 U867 ( .A1(n780), .A2(n779), .ZN(G282) );
  NAND2_X1 U868 ( .A1(n894), .A2(G123), .ZN(n781) );
  XNOR2_X1 U869 ( .A(n781), .B(KEYINPUT18), .ZN(n783) );
  NAND2_X1 U870 ( .A1(G111), .A2(n895), .ZN(n782) );
  NAND2_X1 U871 ( .A1(n783), .A2(n782), .ZN(n787) );
  NAND2_X1 U872 ( .A1(G135), .A2(n890), .ZN(n785) );
  NAND2_X1 U873 ( .A1(G99), .A2(n891), .ZN(n784) );
  NAND2_X1 U874 ( .A1(n785), .A2(n784), .ZN(n786) );
  NOR2_X1 U875 ( .A1(n787), .A2(n786), .ZN(n996) );
  XNOR2_X1 U876 ( .A(G2096), .B(n996), .ZN(n789) );
  INV_X1 U877 ( .A(G2100), .ZN(n788) );
  NAND2_X1 U878 ( .A1(n789), .A2(n788), .ZN(G156) );
  INV_X1 U879 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U880 ( .A(G288), .B(KEYINPUT19), .ZN(n791) );
  XNOR2_X1 U881 ( .A(n953), .B(G166), .ZN(n790) );
  XNOR2_X1 U882 ( .A(n791), .B(n790), .ZN(n805) );
  XNOR2_X1 U883 ( .A(G290), .B(G305), .ZN(n803) );
  NAND2_X1 U884 ( .A1(G80), .A2(n792), .ZN(n795) );
  NAND2_X1 U885 ( .A1(G55), .A2(n793), .ZN(n794) );
  NAND2_X1 U886 ( .A1(n795), .A2(n794), .ZN(n801) );
  NAND2_X1 U887 ( .A1(n796), .A2(G67), .ZN(n799) );
  NAND2_X1 U888 ( .A1(G93), .A2(n797), .ZN(n798) );
  NAND2_X1 U889 ( .A1(n799), .A2(n798), .ZN(n800) );
  NOR2_X1 U890 ( .A1(n801), .A2(n800), .ZN(n802) );
  XOR2_X1 U891 ( .A(n802), .B(KEYINPUT76), .Z(n835) );
  XOR2_X1 U892 ( .A(n803), .B(n835), .Z(n804) );
  XNOR2_X1 U893 ( .A(n805), .B(n804), .ZN(n840) );
  NAND2_X1 U894 ( .A1(G559), .A2(n841), .ZN(n806) );
  XOR2_X1 U895 ( .A(n936), .B(n806), .Z(n833) );
  XOR2_X1 U896 ( .A(n840), .B(n833), .Z(n807) );
  NOR2_X1 U897 ( .A1(n808), .A2(n807), .ZN(n810) );
  NOR2_X1 U898 ( .A1(n835), .A2(G868), .ZN(n809) );
  NOR2_X1 U899 ( .A1(n810), .A2(n809), .ZN(G295) );
  NAND2_X1 U900 ( .A1(G2078), .A2(G2084), .ZN(n812) );
  XOR2_X1 U901 ( .A(KEYINPUT20), .B(KEYINPUT82), .Z(n811) );
  XNOR2_X1 U902 ( .A(n812), .B(n811), .ZN(n813) );
  NAND2_X1 U903 ( .A1(G2090), .A2(n813), .ZN(n814) );
  XNOR2_X1 U904 ( .A(KEYINPUT21), .B(n814), .ZN(n815) );
  NAND2_X1 U905 ( .A1(n815), .A2(G2072), .ZN(n816) );
  XOR2_X1 U906 ( .A(KEYINPUT83), .B(n816), .Z(G158) );
  XNOR2_X1 U907 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U908 ( .A1(G220), .A2(G219), .ZN(n817) );
  XOR2_X1 U909 ( .A(KEYINPUT22), .B(n817), .Z(n818) );
  NOR2_X1 U910 ( .A1(G218), .A2(n818), .ZN(n819) );
  NAND2_X1 U911 ( .A1(G96), .A2(n819), .ZN(n838) );
  NAND2_X1 U912 ( .A1(n838), .A2(G2106), .ZN(n825) );
  NOR2_X1 U913 ( .A1(G235), .A2(G236), .ZN(n820) );
  XNOR2_X1 U914 ( .A(KEYINPUT84), .B(n820), .ZN(n821) );
  NAND2_X1 U915 ( .A1(n821), .A2(G57), .ZN(n822) );
  NOR2_X1 U916 ( .A1(n822), .A2(G238), .ZN(n823) );
  XNOR2_X1 U917 ( .A(n823), .B(KEYINPUT85), .ZN(n837) );
  NAND2_X1 U918 ( .A1(n837), .A2(G567), .ZN(n824) );
  NAND2_X1 U919 ( .A1(n825), .A2(n824), .ZN(n915) );
  NAND2_X1 U920 ( .A1(G661), .A2(G483), .ZN(n826) );
  NOR2_X1 U921 ( .A1(n915), .A2(n826), .ZN(n832) );
  NAND2_X1 U922 ( .A1(G36), .A2(n832), .ZN(n827) );
  XNOR2_X1 U923 ( .A(n827), .B(KEYINPUT86), .ZN(G176) );
  NAND2_X1 U924 ( .A1(n828), .A2(G2106), .ZN(n829) );
  XNOR2_X1 U925 ( .A(n829), .B(KEYINPUT104), .ZN(G217) );
  AND2_X1 U926 ( .A1(G15), .A2(G2), .ZN(n830) );
  NAND2_X1 U927 ( .A1(G661), .A2(n830), .ZN(G259) );
  NAND2_X1 U928 ( .A1(G3), .A2(G1), .ZN(n831) );
  NAND2_X1 U929 ( .A1(n832), .A2(n831), .ZN(G188) );
  NAND2_X1 U931 ( .A1(n834), .A2(n833), .ZN(n836) );
  XNOR2_X1 U932 ( .A(n836), .B(n835), .ZN(G145) );
  INV_X1 U933 ( .A(G96), .ZN(G221) );
  INV_X1 U934 ( .A(G57), .ZN(G237) );
  NOR2_X1 U935 ( .A1(n838), .A2(n837), .ZN(n839) );
  XNOR2_X1 U936 ( .A(n839), .B(KEYINPUT105), .ZN(G261) );
  INV_X1 U937 ( .A(G261), .ZN(G325) );
  XNOR2_X1 U938 ( .A(n936), .B(n840), .ZN(n843) );
  XNOR2_X1 U939 ( .A(G171), .B(n841), .ZN(n842) );
  XNOR2_X1 U940 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U941 ( .A(G286), .B(n844), .Z(n845) );
  NOR2_X1 U942 ( .A1(G37), .A2(n845), .ZN(G397) );
  XOR2_X1 U943 ( .A(G2096), .B(KEYINPUT106), .Z(n847) );
  XNOR2_X1 U944 ( .A(G2090), .B(KEYINPUT43), .ZN(n846) );
  XNOR2_X1 U945 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U946 ( .A(n848), .B(KEYINPUT42), .Z(n850) );
  XNOR2_X1 U947 ( .A(G2067), .B(G2072), .ZN(n849) );
  XNOR2_X1 U948 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U949 ( .A(G2678), .B(G2100), .Z(n852) );
  XNOR2_X1 U950 ( .A(G2078), .B(G2084), .ZN(n851) );
  XNOR2_X1 U951 ( .A(n852), .B(n851), .ZN(n853) );
  XNOR2_X1 U952 ( .A(n854), .B(n853), .ZN(G227) );
  XOR2_X1 U953 ( .A(G1971), .B(G1956), .Z(n856) );
  XNOR2_X1 U954 ( .A(G1986), .B(G1961), .ZN(n855) );
  XNOR2_X1 U955 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U956 ( .A(G1981), .B(G1966), .Z(n858) );
  XNOR2_X1 U957 ( .A(G1996), .B(G1991), .ZN(n857) );
  XNOR2_X1 U958 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U959 ( .A(n860), .B(n859), .Z(n862) );
  XNOR2_X1 U960 ( .A(KEYINPUT107), .B(G2474), .ZN(n861) );
  XNOR2_X1 U961 ( .A(n862), .B(n861), .ZN(n864) );
  XOR2_X1 U962 ( .A(G1976), .B(KEYINPUT41), .Z(n863) );
  XNOR2_X1 U963 ( .A(n864), .B(n863), .ZN(G229) );
  NAND2_X1 U964 ( .A1(G100), .A2(n891), .ZN(n865) );
  XNOR2_X1 U965 ( .A(n865), .B(KEYINPUT108), .ZN(n872) );
  NAND2_X1 U966 ( .A1(G136), .A2(n890), .ZN(n867) );
  NAND2_X1 U967 ( .A1(G112), .A2(n895), .ZN(n866) );
  NAND2_X1 U968 ( .A1(n867), .A2(n866), .ZN(n870) );
  NAND2_X1 U969 ( .A1(n894), .A2(G124), .ZN(n868) );
  XOR2_X1 U970 ( .A(KEYINPUT44), .B(n868), .Z(n869) );
  NOR2_X1 U971 ( .A1(n870), .A2(n869), .ZN(n871) );
  NAND2_X1 U972 ( .A1(n872), .A2(n871), .ZN(n873) );
  XNOR2_X1 U973 ( .A(KEYINPUT109), .B(n873), .ZN(G162) );
  XOR2_X1 U974 ( .A(G160), .B(G162), .Z(n874) );
  XNOR2_X1 U975 ( .A(n875), .B(n874), .ZN(n880) );
  XNOR2_X1 U976 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n878) );
  XNOR2_X1 U977 ( .A(n876), .B(KEYINPUT110), .ZN(n877) );
  XNOR2_X1 U978 ( .A(n878), .B(n877), .ZN(n879) );
  XOR2_X1 U979 ( .A(n880), .B(n879), .Z(n882) );
  XNOR2_X1 U980 ( .A(G164), .B(n996), .ZN(n881) );
  XNOR2_X1 U981 ( .A(n882), .B(n881), .ZN(n906) );
  NAND2_X1 U982 ( .A1(G130), .A2(n894), .ZN(n884) );
  NAND2_X1 U983 ( .A1(G118), .A2(n895), .ZN(n883) );
  NAND2_X1 U984 ( .A1(n884), .A2(n883), .ZN(n889) );
  NAND2_X1 U985 ( .A1(G142), .A2(n890), .ZN(n886) );
  NAND2_X1 U986 ( .A1(G106), .A2(n891), .ZN(n885) );
  NAND2_X1 U987 ( .A1(n886), .A2(n885), .ZN(n887) );
  XOR2_X1 U988 ( .A(n887), .B(KEYINPUT45), .Z(n888) );
  NOR2_X1 U989 ( .A1(n889), .A2(n888), .ZN(n902) );
  NAND2_X1 U990 ( .A1(G139), .A2(n890), .ZN(n893) );
  NAND2_X1 U991 ( .A1(G103), .A2(n891), .ZN(n892) );
  NAND2_X1 U992 ( .A1(n893), .A2(n892), .ZN(n900) );
  NAND2_X1 U993 ( .A1(G127), .A2(n894), .ZN(n897) );
  NAND2_X1 U994 ( .A1(G115), .A2(n895), .ZN(n896) );
  NAND2_X1 U995 ( .A1(n897), .A2(n896), .ZN(n898) );
  XOR2_X1 U996 ( .A(KEYINPUT47), .B(n898), .Z(n899) );
  NOR2_X1 U997 ( .A1(n900), .A2(n899), .ZN(n901) );
  XNOR2_X1 U998 ( .A(KEYINPUT111), .B(n901), .ZN(n998) );
  XNOR2_X1 U999 ( .A(n902), .B(n998), .ZN(n903) );
  XOR2_X1 U1000 ( .A(n904), .B(n903), .Z(n905) );
  XNOR2_X1 U1001 ( .A(n906), .B(n905), .ZN(n907) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n907), .ZN(n908) );
  XNOR2_X1 U1003 ( .A(KEYINPUT112), .B(n908), .ZN(G395) );
  NOR2_X1 U1004 ( .A1(G227), .A2(G229), .ZN(n909) );
  XNOR2_X1 U1005 ( .A(KEYINPUT49), .B(n909), .ZN(n910) );
  NOR2_X1 U1006 ( .A1(G397), .A2(n910), .ZN(n914) );
  NOR2_X1 U1007 ( .A1(G401), .A2(n915), .ZN(n911) );
  XNOR2_X1 U1008 ( .A(KEYINPUT113), .B(n911), .ZN(n912) );
  NOR2_X1 U1009 ( .A1(G395), .A2(n912), .ZN(n913) );
  NAND2_X1 U1010 ( .A1(n914), .A2(n913), .ZN(G225) );
  INV_X1 U1011 ( .A(G225), .ZN(G308) );
  INV_X1 U1012 ( .A(n915), .ZN(G319) );
  XNOR2_X1 U1013 ( .A(G1996), .B(G32), .ZN(n917) );
  XNOR2_X1 U1014 ( .A(G33), .B(G2072), .ZN(n916) );
  NOR2_X1 U1015 ( .A1(n917), .A2(n916), .ZN(n922) );
  XOR2_X1 U1016 ( .A(G1991), .B(G25), .Z(n918) );
  NAND2_X1 U1017 ( .A1(n918), .A2(G28), .ZN(n920) );
  XNOR2_X1 U1018 ( .A(G26), .B(G2067), .ZN(n919) );
  NOR2_X1 U1019 ( .A1(n920), .A2(n919), .ZN(n921) );
  NAND2_X1 U1020 ( .A1(n922), .A2(n921), .ZN(n925) );
  XOR2_X1 U1021 ( .A(G27), .B(n923), .Z(n924) );
  NOR2_X1 U1022 ( .A1(n925), .A2(n924), .ZN(n926) );
  XOR2_X1 U1023 ( .A(KEYINPUT53), .B(n926), .Z(n930) );
  XNOR2_X1 U1024 ( .A(KEYINPUT54), .B(G34), .ZN(n927) );
  XNOR2_X1 U1025 ( .A(n927), .B(KEYINPUT115), .ZN(n928) );
  XNOR2_X1 U1026 ( .A(G2084), .B(n928), .ZN(n929) );
  NAND2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(n932) );
  XNOR2_X1 U1028 ( .A(G35), .B(G2090), .ZN(n931) );
  NOR2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1030 ( .A(KEYINPUT55), .B(n933), .Z(n934) );
  NOR2_X1 U1031 ( .A1(G29), .A2(n934), .ZN(n994) );
  XOR2_X1 U1032 ( .A(G16), .B(KEYINPUT56), .Z(n962) );
  XOR2_X1 U1033 ( .A(G1341), .B(KEYINPUT119), .Z(n935) );
  XNOR2_X1 U1034 ( .A(n936), .B(n935), .ZN(n960) );
  XNOR2_X1 U1035 ( .A(G168), .B(G1966), .ZN(n938) );
  NAND2_X1 U1036 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1037 ( .A(n939), .B(KEYINPUT57), .ZN(n946) );
  AND2_X1 U1038 ( .A1(G303), .A2(G1971), .ZN(n943) );
  NAND2_X1 U1039 ( .A1(n941), .A2(n940), .ZN(n942) );
  NOR2_X1 U1040 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1041 ( .A(n944), .B(KEYINPUT118), .ZN(n945) );
  NAND2_X1 U1042 ( .A1(n946), .A2(n945), .ZN(n952) );
  XNOR2_X1 U1043 ( .A(G301), .B(G1961), .ZN(n949) );
  XNOR2_X1 U1044 ( .A(n947), .B(G1348), .ZN(n948) );
  NOR2_X1 U1045 ( .A1(n949), .A2(n948), .ZN(n950) );
  XOR2_X1 U1046 ( .A(KEYINPUT116), .B(n950), .Z(n951) );
  NOR2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n958) );
  XNOR2_X1 U1048 ( .A(n953), .B(G1956), .ZN(n954) );
  XNOR2_X1 U1049 ( .A(n954), .B(KEYINPUT117), .ZN(n956) );
  NOR2_X1 U1050 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1051 ( .A1(n958), .A2(n957), .ZN(n959) );
  NOR2_X1 U1052 ( .A1(n960), .A2(n959), .ZN(n961) );
  NOR2_X1 U1053 ( .A1(n962), .A2(n961), .ZN(n991) );
  XOR2_X1 U1054 ( .A(G16), .B(KEYINPUT120), .Z(n988) );
  XOR2_X1 U1055 ( .A(KEYINPUT60), .B(KEYINPUT123), .Z(n973) );
  XOR2_X1 U1056 ( .A(KEYINPUT122), .B(G4), .Z(n964) );
  XNOR2_X1 U1057 ( .A(G1348), .B(KEYINPUT59), .ZN(n963) );
  XNOR2_X1 U1058 ( .A(n964), .B(n963), .ZN(n967) );
  XOR2_X1 U1059 ( .A(KEYINPUT121), .B(G1981), .Z(n965) );
  XNOR2_X1 U1060 ( .A(G6), .B(n965), .ZN(n966) );
  NOR2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(n971) );
  XNOR2_X1 U1062 ( .A(G1956), .B(G20), .ZN(n969) );
  XNOR2_X1 U1063 ( .A(G19), .B(G1341), .ZN(n968) );
  NOR2_X1 U1064 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1065 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1066 ( .A(n973), .B(n972), .ZN(n985) );
  XNOR2_X1 U1067 ( .A(G1971), .B(G22), .ZN(n975) );
  XNOR2_X1 U1068 ( .A(G23), .B(G1976), .ZN(n974) );
  NOR2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n977) );
  XOR2_X1 U1070 ( .A(G1986), .B(G24), .Z(n976) );
  NAND2_X1 U1071 ( .A1(n977), .A2(n976), .ZN(n979) );
  XOR2_X1 U1072 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n978) );
  XNOR2_X1 U1073 ( .A(n979), .B(n978), .ZN(n983) );
  XNOR2_X1 U1074 ( .A(G1961), .B(G5), .ZN(n981) );
  XNOR2_X1 U1075 ( .A(G21), .B(G1966), .ZN(n980) );
  NOR2_X1 U1076 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1077 ( .A1(n983), .A2(n982), .ZN(n984) );
  NOR2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1079 ( .A(KEYINPUT61), .B(n986), .ZN(n987) );
  NAND2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1081 ( .A(KEYINPUT125), .B(n989), .ZN(n990) );
  NOR2_X1 U1082 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1083 ( .A1(G11), .A2(n992), .ZN(n993) );
  NOR2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1085 ( .A(KEYINPUT126), .B(n995), .ZN(n1023) );
  NOR2_X1 U1086 ( .A1(n997), .A2(n996), .ZN(n1008) );
  XNOR2_X1 U1087 ( .A(G2072), .B(KEYINPUT114), .ZN(n999) );
  XNOR2_X1 U1088 ( .A(n999), .B(n998), .ZN(n1001) );
  XOR2_X1 U1089 ( .A(G164), .B(G2078), .Z(n1000) );
  NOR2_X1 U1090 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1091 ( .A(KEYINPUT50), .B(n1002), .ZN(n1004) );
  XNOR2_X1 U1092 ( .A(G160), .B(G2084), .ZN(n1003) );
  NAND2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1095 ( .A1(n1008), .A2(n1007), .ZN(n1013) );
  XOR2_X1 U1096 ( .A(G2090), .B(G162), .Z(n1009) );
  NOR2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1098 ( .A(KEYINPUT51), .B(n1011), .ZN(n1012) );
  NOR2_X1 U1099 ( .A1(n1013), .A2(n1012), .ZN(n1015) );
  NAND2_X1 U1100 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1101 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1102 ( .A(KEYINPUT52), .B(n1018), .ZN(n1020) );
  INV_X1 U1103 ( .A(KEYINPUT55), .ZN(n1019) );
  NAND2_X1 U1104 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1105 ( .A1(n1021), .A2(G29), .ZN(n1022) );
  NAND2_X1 U1106 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1107 ( .A(n1024), .B(KEYINPUT62), .ZN(n1025) );
  XNOR2_X1 U1108 ( .A(KEYINPUT127), .B(n1025), .ZN(G311) );
  INV_X1 U1109 ( .A(G311), .ZN(G150) );
endmodule

