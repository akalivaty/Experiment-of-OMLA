

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777;

  XNOR2_X1 U378 ( .A(n561), .B(n532), .ZN(n701) );
  INV_X1 U379 ( .A(n553), .ZN(n691) );
  XOR2_X1 U380 ( .A(n447), .B(n467), .Z(n357) );
  NOR2_X2 U381 ( .A1(n580), .A2(n717), .ZN(n582) );
  XNOR2_X2 U382 ( .A(n539), .B(n368), .ZN(n594) );
  XNOR2_X2 U383 ( .A(KEYINPUT18), .B(KEYINPUT78), .ZN(n455) );
  OR2_X2 U384 ( .A1(n372), .A2(n514), .ZN(n605) );
  OR2_X1 U385 ( .A1(n748), .A2(n749), .ZN(n385) );
  XNOR2_X1 U386 ( .A(n391), .B(KEYINPUT89), .ZN(n648) );
  NAND2_X1 U387 ( .A1(n742), .A2(n648), .ZN(n737) );
  XNOR2_X1 U388 ( .A(n575), .B(n574), .ZN(n393) );
  XNOR2_X1 U389 ( .A(n501), .B(KEYINPUT4), .ZN(n463) );
  NOR2_X1 U390 ( .A1(n453), .A2(n452), .ZN(n533) );
  XNOR2_X1 U391 ( .A(n535), .B(KEYINPUT40), .ZN(n545) );
  XNOR2_X1 U392 ( .A(n427), .B(n362), .ZN(n358) );
  XNOR2_X1 U393 ( .A(n427), .B(n362), .ZN(n713) );
  BUF_X1 U394 ( .A(n397), .Z(n359) );
  XNOR2_X1 U395 ( .A(n378), .B(KEYINPUT0), .ZN(n360) );
  XNOR2_X1 U396 ( .A(n621), .B(n620), .ZN(n361) );
  XNOR2_X1 U397 ( .A(n378), .B(KEYINPUT0), .ZN(n585) );
  XNOR2_X1 U398 ( .A(n621), .B(n620), .ZN(n742) );
  XNOR2_X1 U399 ( .A(n650), .B(G146), .ZN(n441) );
  NOR2_X1 U400 ( .A1(n558), .A2(n401), .ZN(n400) );
  NAND2_X1 U401 ( .A1(n539), .A2(n538), .ZN(n401) );
  XNOR2_X1 U402 ( .A(n463), .B(n363), .ZN(n650) );
  NAND2_X1 U403 ( .A1(n640), .A2(n486), .ZN(n448) );
  INV_X1 U404 ( .A(KEYINPUT44), .ZN(n373) );
  NAND2_X1 U405 ( .A1(n573), .A2(n572), .ZN(n575) );
  XNOR2_X1 U406 ( .A(G122), .B(G104), .ZN(n481) );
  INV_X1 U407 ( .A(G137), .ZN(n404) );
  XNOR2_X1 U408 ( .A(n403), .B(n420), .ZN(n375) );
  XOR2_X1 U409 ( .A(G107), .B(G101), .Z(n403) );
  NOR2_X1 U410 ( .A1(n580), .A2(n366), .ZN(n525) );
  XNOR2_X1 U411 ( .A(n410), .B(n409), .ZN(n540) );
  NOR2_X1 U412 ( .A1(n672), .A2(G902), .ZN(n410) );
  XNOR2_X1 U413 ( .A(n540), .B(KEYINPUT1), .ZN(n718) );
  XNOR2_X1 U414 ( .A(n357), .B(n441), .ZN(n640) );
  NAND2_X1 U415 ( .A1(n512), .A2(n519), .ZN(n558) );
  BUF_X1 U416 ( .A(n718), .Z(n374) );
  NOR2_X1 U417 ( .A1(n396), .A2(n395), .ZN(n394) );
  INV_X1 U418 ( .A(G210), .ZN(n395) );
  INV_X1 U419 ( .A(n638), .ZN(n396) );
  XNOR2_X1 U420 ( .A(G902), .B(KEYINPUT15), .ZN(n627) );
  XNOR2_X1 U421 ( .A(n386), .B(KEYINPUT19), .ZN(n548) );
  XOR2_X1 U422 ( .A(KEYINPUT5), .B(G116), .Z(n443) );
  AND2_X1 U423 ( .A1(n775), .A2(n577), .ZN(n392) );
  INV_X1 U424 ( .A(G116), .ZN(n466) );
  XNOR2_X1 U425 ( .A(G143), .B(G131), .ZN(n478) );
  XNOR2_X1 U426 ( .A(KEYINPUT93), .B(KEYINPUT94), .ZN(n460) );
  XNOR2_X1 U427 ( .A(KEYINPUT66), .B(KEYINPUT45), .ZN(n620) );
  XNOR2_X1 U428 ( .A(n377), .B(n376), .ZN(n707) );
  INV_X1 U429 ( .A(KEYINPUT106), .ZN(n376) );
  INV_X1 U430 ( .A(G902), .ZN(n486) );
  BUF_X1 U431 ( .A(n648), .Z(n741) );
  BUF_X1 U432 ( .A(n361), .Z(n761) );
  XNOR2_X1 U433 ( .A(G119), .B(G128), .ZN(n412) );
  XNOR2_X1 U434 ( .A(KEYINPUT24), .B(G110), .ZN(n411) );
  XNOR2_X1 U435 ( .A(KEYINPUT96), .B(KEYINPUT97), .ZN(n414) );
  XNOR2_X1 U436 ( .A(KEYINPUT23), .B(KEYINPUT95), .ZN(n413) );
  XNOR2_X1 U437 ( .A(n490), .B(n489), .ZN(n494) );
  XNOR2_X1 U438 ( .A(G134), .B(G122), .ZN(n489) );
  XOR2_X1 U439 ( .A(KEYINPUT7), .B(KEYINPUT104), .Z(n492) );
  XNOR2_X1 U440 ( .A(n375), .B(n364), .ZN(n406) );
  NOR2_X1 U441 ( .A1(n542), .A2(n541), .ZN(n550) );
  XNOR2_X1 U442 ( .A(n400), .B(n399), .ZN(n542) );
  INV_X1 U443 ( .A(KEYINPUT28), .ZN(n399) );
  BUF_X1 U444 ( .A(n360), .Z(n583) );
  OR2_X1 U445 ( .A1(n552), .A2(n551), .ZN(n553) );
  INV_X1 U446 ( .A(KEYINPUT6), .ZN(n368) );
  XNOR2_X1 U447 ( .A(n640), .B(n639), .ZN(n641) );
  XOR2_X1 U448 ( .A(n664), .B(KEYINPUT59), .Z(n665) );
  AND2_X1 U449 ( .A1(n560), .A2(n380), .ZN(n562) );
  AND2_X1 U450 ( .A1(n559), .A2(n381), .ZN(n380) );
  AND2_X1 U451 ( .A1(n552), .A2(n551), .ZN(n694) );
  AND2_X2 U452 ( .A1(n589), .A2(n717), .ZN(n681) );
  XNOR2_X1 U453 ( .A(n398), .B(n755), .ZN(n757) );
  INV_X1 U454 ( .A(KEYINPUT53), .ZN(n382) );
  NAND2_X1 U455 ( .A1(n550), .A2(n549), .ZN(n389) );
  XOR2_X1 U456 ( .A(n426), .B(KEYINPUT25), .Z(n362) );
  BUF_X1 U457 ( .A(n505), .Z(n561) );
  XOR2_X1 U458 ( .A(G134), .B(G131), .Z(n363) );
  AND2_X1 U459 ( .A1(n393), .A2(n577), .ZN(n633) );
  AND2_X1 U460 ( .A1(n434), .A2(G227), .ZN(n364) );
  AND2_X1 U461 ( .A1(n538), .A2(n702), .ZN(n365) );
  INV_X1 U462 ( .A(n389), .ZN(n565) );
  INV_X1 U463 ( .A(n702), .ZN(n387) );
  INV_X1 U464 ( .A(G953), .ZN(n760) );
  AND2_X1 U465 ( .A1(n594), .A2(n365), .ZN(n517) );
  INV_X1 U466 ( .A(n594), .ZN(n366) );
  XNOR2_X1 U467 ( .A(n594), .B(n367), .ZN(n600) );
  INV_X1 U468 ( .A(KEYINPUT82), .ZN(n367) );
  NAND2_X1 U469 ( .A1(n701), .A2(n702), .ZN(n377) );
  XNOR2_X1 U470 ( .A(n588), .B(KEYINPUT98), .ZN(n589) );
  BUF_X1 U471 ( .A(n659), .Z(n369) );
  BUF_X1 U472 ( .A(n774), .Z(n370) );
  BUF_X1 U473 ( .A(n548), .Z(n371) );
  XNOR2_X1 U474 ( .A(n511), .B(KEYINPUT22), .ZN(n372) );
  XNOR2_X1 U475 ( .A(n511), .B(KEYINPUT22), .ZN(n603) );
  XNOR2_X1 U476 ( .A(n456), .B(n457), .ZN(n459) );
  AND2_X1 U477 ( .A1(n706), .A2(n549), .ZN(n390) );
  XNOR2_X1 U478 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U479 ( .A(n499), .B(n500), .ZN(n502) );
  AND2_X1 U480 ( .A1(n613), .A2(n373), .ZN(n615) );
  NAND2_X1 U481 ( .A1(n733), .A2(n550), .ZN(n544) );
  XNOR2_X2 U482 ( .A(n537), .B(KEYINPUT41), .ZN(n733) );
  NOR2_X2 U483 ( .A1(n548), .A2(n509), .ZN(n378) );
  XNOR2_X1 U484 ( .A(n379), .B(n419), .ZN(n422) );
  NAND2_X1 U485 ( .A1(n418), .A2(G221), .ZN(n379) );
  INV_X1 U486 ( .A(n358), .ZN(n512) );
  NAND2_X1 U487 ( .A1(n713), .A2(n714), .ZN(n433) );
  NOR2_X1 U488 ( .A1(n569), .A2(n568), .ZN(n571) );
  INV_X1 U489 ( .A(n561), .ZN(n381) );
  XNOR2_X2 U490 ( .A(n534), .B(KEYINPUT39), .ZN(n578) );
  XNOR2_X1 U491 ( .A(n383), .B(n382), .ZN(G75) );
  NAND2_X1 U492 ( .A1(n384), .A2(n760), .ZN(n383) );
  XNOR2_X1 U493 ( .A(n385), .B(n750), .ZN(n384) );
  NOR2_X2 U494 ( .A1(n505), .A2(n387), .ZN(n386) );
  XNOR2_X2 U495 ( .A(n473), .B(n472), .ZN(n505) );
  NAND2_X1 U496 ( .A1(n388), .A2(KEYINPUT47), .ZN(n556) );
  NAND2_X1 U497 ( .A1(n390), .A2(n550), .ZN(n388) );
  NAND2_X1 U498 ( .A1(n393), .A2(n392), .ZN(n391) );
  AND2_X2 U499 ( .A1(n397), .A2(n638), .ZN(n751) );
  XNOR2_X2 U500 ( .A(n632), .B(KEYINPUT67), .ZN(n397) );
  NAND2_X1 U501 ( .A1(n359), .A2(n394), .ZN(n398) );
  INV_X1 U502 ( .A(KEYINPUT48), .ZN(n574) );
  XNOR2_X1 U503 ( .A(n442), .B(G137), .ZN(n444) );
  INV_X1 U504 ( .A(n576), .ZN(n577) );
  INV_X1 U505 ( .A(KEYINPUT70), .ZN(n432) );
  XNOR2_X1 U506 ( .A(n444), .B(n443), .ZN(n447) );
  XNOR2_X1 U507 ( .A(n417), .B(KEYINPUT8), .ZN(n496) );
  INV_X1 U508 ( .A(KEYINPUT103), .ZN(n497) );
  INV_X1 U509 ( .A(n746), .ZN(n638) );
  INV_X1 U510 ( .A(KEYINPUT99), .ZN(n581) );
  BUF_X1 U511 ( .A(n545), .Z(n536) );
  XNOR2_X2 U512 ( .A(G143), .B(G128), .ZN(n501) );
  INV_X2 U513 ( .A(KEYINPUT64), .ZN(n402) );
  XNOR2_X2 U514 ( .A(n402), .B(G953), .ZN(n454) );
  XNOR2_X1 U515 ( .A(n404), .B(G140), .ZN(n420) );
  XNOR2_X1 U516 ( .A(G110), .B(KEYINPUT76), .ZN(n768) );
  XNOR2_X1 U517 ( .A(n768), .B(KEYINPUT73), .ZN(n458) );
  XNOR2_X1 U518 ( .A(G104), .B(n458), .ZN(n405) );
  XNOR2_X1 U519 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U520 ( .A(n441), .B(n407), .ZN(n672) );
  INV_X1 U521 ( .A(KEYINPUT72), .ZN(n408) );
  XNOR2_X1 U522 ( .A(n408), .B(G469), .ZN(n409) );
  XNOR2_X1 U523 ( .A(n412), .B(n411), .ZN(n416) );
  XNOR2_X1 U524 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U525 ( .A(n416), .B(n415), .ZN(n419) );
  NAND2_X1 U526 ( .A1(n454), .A2(G234), .ZN(n417) );
  INV_X1 U527 ( .A(n496), .ZN(n418) );
  XNOR2_X1 U528 ( .A(G146), .B(G125), .ZN(n461) );
  XNOR2_X1 U529 ( .A(n461), .B(KEYINPUT10), .ZN(n483) );
  INV_X1 U530 ( .A(n420), .ZN(n421) );
  XNOR2_X1 U531 ( .A(n483), .B(n421), .ZN(n649) );
  XNOR2_X1 U532 ( .A(n422), .B(n649), .ZN(n659) );
  OR2_X2 U533 ( .A1(n659), .A2(G902), .ZN(n427) );
  NAND2_X1 U534 ( .A1(n627), .A2(G234), .ZN(n424) );
  INV_X1 U535 ( .A(KEYINPUT20), .ZN(n423) );
  XNOR2_X1 U536 ( .A(n424), .B(n423), .ZN(n429) );
  INV_X1 U537 ( .A(n429), .ZN(n425) );
  NAND2_X1 U538 ( .A1(n425), .A2(G217), .ZN(n426) );
  INV_X1 U539 ( .A(G221), .ZN(n428) );
  OR2_X1 U540 ( .A1(n429), .A2(n428), .ZN(n431) );
  INV_X1 U541 ( .A(KEYINPUT21), .ZN(n430) );
  XNOR2_X1 U542 ( .A(n431), .B(n430), .ZN(n714) );
  XNOR2_X2 U543 ( .A(n433), .B(n432), .ZN(n719) );
  NAND2_X1 U544 ( .A1(n540), .A2(n719), .ZN(n586) );
  BUF_X1 U545 ( .A(n454), .Z(n434) );
  INV_X1 U546 ( .A(n434), .ZN(n644) );
  NOR2_X1 U547 ( .A1(n486), .A2(G900), .ZN(n435) );
  NAND2_X1 U548 ( .A1(n644), .A2(n435), .ZN(n436) );
  NAND2_X1 U549 ( .A1(n760), .A2(G952), .ZN(n506) );
  NAND2_X1 U550 ( .A1(n436), .A2(n506), .ZN(n538) );
  NAND2_X1 U551 ( .A1(G237), .A2(G234), .ZN(n438) );
  INV_X1 U552 ( .A(KEYINPUT14), .ZN(n437) );
  XNOR2_X1 U553 ( .A(n438), .B(n437), .ZN(n731) );
  INV_X1 U554 ( .A(n731), .ZN(n518) );
  NAND2_X1 U555 ( .A1(n538), .A2(n518), .ZN(n439) );
  NOR2_X2 U556 ( .A1(n586), .A2(n439), .ZN(n440) );
  XNOR2_X1 U557 ( .A(n440), .B(KEYINPUT77), .ZN(n453) );
  NOR2_X1 U558 ( .A1(G953), .A2(G237), .ZN(n474) );
  NAND2_X1 U559 ( .A1(n474), .A2(G210), .ZN(n442) );
  XNOR2_X1 U560 ( .A(G113), .B(G101), .ZN(n446) );
  XNOR2_X1 U561 ( .A(KEYINPUT3), .B(G119), .ZN(n445) );
  XNOR2_X1 U562 ( .A(n446), .B(n445), .ZN(n467) );
  XNOR2_X2 U563 ( .A(n448), .B(G472), .ZN(n539) );
  INV_X1 U564 ( .A(G237), .ZN(n449) );
  NAND2_X1 U565 ( .A1(n486), .A2(n449), .ZN(n471) );
  NAND2_X1 U566 ( .A1(n471), .A2(G214), .ZN(n702) );
  NAND2_X1 U567 ( .A1(n539), .A2(n702), .ZN(n451) );
  XOR2_X1 U568 ( .A(KEYINPUT105), .B(KEYINPUT30), .Z(n450) );
  XNOR2_X1 U569 ( .A(n451), .B(n450), .ZN(n452) );
  NAND2_X1 U570 ( .A1(n454), .A2(G224), .ZN(n457) );
  XNOR2_X1 U571 ( .A(n455), .B(KEYINPUT17), .ZN(n456) );
  XNOR2_X1 U572 ( .A(n459), .B(n458), .ZN(n465) );
  XNOR2_X1 U573 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U574 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U575 ( .A(n465), .B(n464), .ZN(n470) );
  XNOR2_X1 U576 ( .A(n466), .B(G107), .ZN(n490) );
  XNOR2_X1 U577 ( .A(n467), .B(n490), .ZN(n469) );
  XNOR2_X1 U578 ( .A(n481), .B(KEYINPUT16), .ZN(n468) );
  XNOR2_X1 U579 ( .A(n469), .B(n468), .ZN(n767) );
  XNOR2_X1 U580 ( .A(n470), .B(n767), .ZN(n752) );
  NAND2_X1 U581 ( .A1(n752), .A2(n627), .ZN(n473) );
  NAND2_X1 U582 ( .A1(n471), .A2(G210), .ZN(n472) );
  XOR2_X1 U583 ( .A(KEYINPUT101), .B(KEYINPUT11), .Z(n476) );
  NAND2_X1 U584 ( .A1(G214), .A2(n474), .ZN(n475) );
  XNOR2_X1 U585 ( .A(n476), .B(n475), .ZN(n477) );
  XOR2_X1 U586 ( .A(n477), .B(KEYINPUT12), .Z(n485) );
  XOR2_X1 U587 ( .A(G140), .B(G113), .Z(n479) );
  XNOR2_X1 U588 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U589 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U590 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U591 ( .A(n485), .B(n484), .ZN(n664) );
  NAND2_X1 U592 ( .A1(n664), .A2(n486), .ZN(n488) );
  XNOR2_X1 U593 ( .A(KEYINPUT13), .B(G475), .ZN(n487) );
  XNOR2_X1 U594 ( .A(n488), .B(n487), .ZN(n552) );
  XNOR2_X1 U595 ( .A(KEYINPUT102), .B(KEYINPUT9), .ZN(n491) );
  XNOR2_X1 U596 ( .A(n492), .B(n491), .ZN(n493) );
  XOR2_X1 U597 ( .A(n494), .B(n493), .Z(n500) );
  INV_X1 U598 ( .A(G217), .ZN(n495) );
  NOR2_X1 U599 ( .A1(n496), .A2(n495), .ZN(n498) );
  XNOR2_X1 U600 ( .A(n502), .B(n501), .ZN(n661) );
  NOR2_X1 U601 ( .A1(G902), .A2(n661), .ZN(n503) );
  XNOR2_X1 U602 ( .A(n503), .B(G478), .ZN(n516) );
  NOR2_X1 U603 ( .A1(n552), .A2(n516), .ZN(n528) );
  AND2_X1 U604 ( .A1(n381), .A2(n528), .ZN(n504) );
  NAND2_X1 U605 ( .A1(n533), .A2(n504), .ZN(n555) );
  XNOR2_X1 U606 ( .A(n555), .B(G143), .ZN(G45) );
  NOR2_X1 U607 ( .A1(G898), .A2(n760), .ZN(n769) );
  NAND2_X1 U608 ( .A1(n769), .A2(G902), .ZN(n507) );
  NAND2_X1 U609 ( .A1(n507), .A2(n506), .ZN(n508) );
  NAND2_X1 U610 ( .A1(n508), .A2(n518), .ZN(n509) );
  AND2_X1 U611 ( .A1(n516), .A2(n552), .ZN(n705) );
  AND2_X1 U612 ( .A1(n705), .A2(n714), .ZN(n510) );
  NAND2_X1 U613 ( .A1(n585), .A2(n510), .ZN(n511) );
  INV_X1 U614 ( .A(n539), .ZN(n717) );
  NAND2_X1 U615 ( .A1(n512), .A2(n717), .ZN(n513) );
  OR2_X1 U616 ( .A1(n374), .A2(n513), .ZN(n514) );
  XOR2_X1 U617 ( .A(G110), .B(KEYINPUT113), .Z(n515) );
  XNOR2_X1 U618 ( .A(n605), .B(n515), .ZN(G12) );
  XOR2_X1 U619 ( .A(G140), .B(KEYINPUT119), .Z(n523) );
  INV_X1 U620 ( .A(n516), .ZN(n551) );
  AND2_X1 U621 ( .A1(n517), .A2(n691), .ZN(n560) );
  AND2_X1 U622 ( .A1(n714), .A2(n518), .ZN(n519) );
  NOR2_X1 U623 ( .A1(n374), .A2(n558), .ZN(n520) );
  NAND2_X1 U624 ( .A1(n560), .A2(n520), .ZN(n521) );
  XOR2_X1 U625 ( .A(KEYINPUT43), .B(n521), .Z(n522) );
  NOR2_X1 U626 ( .A1(n522), .A2(n381), .ZN(n576) );
  XOR2_X1 U627 ( .A(n523), .B(n576), .Z(G42) );
  NAND2_X1 U628 ( .A1(n719), .A2(n718), .ZN(n580) );
  XOR2_X1 U629 ( .A(KEYINPUT74), .B(KEYINPUT33), .Z(n524) );
  XNOR2_X1 U630 ( .A(n525), .B(n524), .ZN(n710) );
  NAND2_X1 U631 ( .A1(n710), .A2(n583), .ZN(n527) );
  XOR2_X1 U632 ( .A(KEYINPUT80), .B(KEYINPUT34), .Z(n526) );
  XNOR2_X1 U633 ( .A(n527), .B(n526), .ZN(n529) );
  NAND2_X1 U634 ( .A1(n529), .A2(n528), .ZN(n531) );
  XNOR2_X1 U635 ( .A(KEYINPUT79), .B(KEYINPUT35), .ZN(n530) );
  XNOR2_X1 U636 ( .A(n531), .B(n530), .ZN(n613) );
  XNOR2_X1 U637 ( .A(n613), .B(G122), .ZN(G24) );
  XOR2_X1 U638 ( .A(KEYINPUT75), .B(KEYINPUT38), .Z(n532) );
  NAND2_X1 U639 ( .A1(n533), .A2(n701), .ZN(n534) );
  NAND2_X1 U640 ( .A1(n578), .A2(n691), .ZN(n535) );
  XNOR2_X1 U641 ( .A(n536), .B(G131), .ZN(G33) );
  NAND2_X1 U642 ( .A1(n705), .A2(n707), .ZN(n537) );
  INV_X1 U643 ( .A(n540), .ZN(n541) );
  XOR2_X1 U644 ( .A(KEYINPUT107), .B(KEYINPUT42), .Z(n543) );
  XNOR2_X1 U645 ( .A(n544), .B(n543), .ZN(n776) );
  NAND2_X1 U646 ( .A1(n545), .A2(n776), .ZN(n547) );
  XNOR2_X1 U647 ( .A(KEYINPUT65), .B(KEYINPUT46), .ZN(n546) );
  XNOR2_X1 U648 ( .A(n547), .B(n546), .ZN(n573) );
  INV_X1 U649 ( .A(n371), .ZN(n549) );
  INV_X1 U650 ( .A(n694), .ZN(n554) );
  NAND2_X1 U651 ( .A1(n554), .A2(n553), .ZN(n706) );
  NAND2_X1 U652 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U653 ( .A(n557), .B(KEYINPUT85), .ZN(n564) );
  INV_X1 U654 ( .A(n558), .ZN(n559) );
  XNOR2_X1 U655 ( .A(n562), .B(KEYINPUT36), .ZN(n563) );
  NAND2_X1 U656 ( .A1(n563), .A2(n374), .ZN(n699) );
  NAND2_X1 U657 ( .A1(n564), .A2(n699), .ZN(n569) );
  XNOR2_X1 U658 ( .A(n706), .B(KEYINPUT86), .ZN(n591) );
  INV_X1 U659 ( .A(KEYINPUT47), .ZN(n566) );
  NAND2_X1 U660 ( .A1(n591), .A2(n566), .ZN(n567) );
  NOR2_X1 U661 ( .A1(n389), .A2(n567), .ZN(n568) );
  INV_X1 U662 ( .A(KEYINPUT71), .ZN(n570) );
  XNOR2_X1 U663 ( .A(n571), .B(n570), .ZN(n572) );
  NAND2_X1 U664 ( .A1(n578), .A2(n694), .ZN(n579) );
  XNOR2_X1 U665 ( .A(n579), .B(KEYINPUT108), .ZN(n775) );
  XNOR2_X1 U666 ( .A(n582), .B(n581), .ZN(n724) );
  NAND2_X1 U667 ( .A1(n724), .A2(n583), .ZN(n584) );
  XNOR2_X1 U668 ( .A(n584), .B(KEYINPUT31), .ZN(n695) );
  INV_X1 U669 ( .A(n360), .ZN(n587) );
  NOR2_X1 U670 ( .A1(n587), .A2(n586), .ZN(n588) );
  NOR2_X1 U671 ( .A1(n695), .A2(n681), .ZN(n590) );
  XNOR2_X1 U672 ( .A(n590), .B(KEYINPUT100), .ZN(n593) );
  INV_X1 U673 ( .A(n591), .ZN(n592) );
  NOR2_X1 U674 ( .A1(n593), .A2(n592), .ZN(n598) );
  INV_X1 U675 ( .A(n374), .ZN(n596) );
  NOR2_X1 U676 ( .A1(n594), .A2(n512), .ZN(n595) );
  NAND2_X1 U677 ( .A1(n596), .A2(n595), .ZN(n597) );
  NOR2_X1 U678 ( .A1(n372), .A2(n597), .ZN(n678) );
  NOR2_X1 U679 ( .A1(n598), .A2(n678), .ZN(n610) );
  AND2_X1 U680 ( .A1(n718), .A2(n512), .ZN(n599) );
  AND2_X1 U681 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U682 ( .A(n601), .B(KEYINPUT81), .ZN(n602) );
  NOR2_X1 U683 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U684 ( .A(n604), .B(KEYINPUT32), .ZN(n774) );
  INV_X1 U685 ( .A(n605), .ZN(n606) );
  NOR2_X1 U686 ( .A1(n774), .A2(n606), .ZN(n607) );
  XNOR2_X1 U687 ( .A(n607), .B(KEYINPUT92), .ZN(n612) );
  NAND2_X1 U688 ( .A1(n612), .A2(n613), .ZN(n608) );
  NAND2_X1 U689 ( .A1(n608), .A2(KEYINPUT44), .ZN(n609) );
  NAND2_X1 U690 ( .A1(n609), .A2(n610), .ZN(n611) );
  XNOR2_X1 U691 ( .A(n611), .B(KEYINPUT91), .ZN(n619) );
  BUF_X1 U692 ( .A(n612), .Z(n617) );
  INV_X1 U693 ( .A(KEYINPUT69), .ZN(n614) );
  XNOR2_X1 U694 ( .A(n615), .B(n614), .ZN(n616) );
  NAND2_X1 U695 ( .A1(n617), .A2(n616), .ZN(n618) );
  NAND2_X1 U696 ( .A1(n619), .A2(n618), .ZN(n621) );
  NAND2_X1 U697 ( .A1(KEYINPUT88), .A2(KEYINPUT2), .ZN(n624) );
  INV_X1 U698 ( .A(KEYINPUT2), .ZN(n622) );
  NOR2_X1 U699 ( .A1(n622), .A2(KEYINPUT88), .ZN(n623) );
  NAND2_X1 U700 ( .A1(n627), .A2(n623), .ZN(n626) );
  AND2_X1 U701 ( .A1(n624), .A2(n626), .ZN(n625) );
  NAND2_X1 U702 ( .A1(n737), .A2(n625), .ZN(n631) );
  INV_X1 U703 ( .A(n626), .ZN(n629) );
  INV_X1 U704 ( .A(n627), .ZN(n628) );
  OR2_X1 U705 ( .A1(n629), .A2(n628), .ZN(n630) );
  NAND2_X1 U706 ( .A1(n631), .A2(n630), .ZN(n632) );
  INV_X1 U707 ( .A(n361), .ZN(n637) );
  NAND2_X1 U708 ( .A1(n775), .A2(KEYINPUT2), .ZN(n634) );
  XNOR2_X1 U709 ( .A(n634), .B(KEYINPUT83), .ZN(n635) );
  NAND2_X1 U710 ( .A1(n633), .A2(n635), .ZN(n636) );
  NOR2_X1 U711 ( .A1(n637), .A2(n636), .ZN(n746) );
  NAND2_X1 U712 ( .A1(n751), .A2(G472), .ZN(n642) );
  XOR2_X1 U713 ( .A(KEYINPUT109), .B(KEYINPUT62), .Z(n639) );
  XNOR2_X1 U714 ( .A(n642), .B(n641), .ZN(n645) );
  INV_X1 U715 ( .A(G952), .ZN(n643) );
  NAND2_X1 U716 ( .A1(n644), .A2(n643), .ZN(n667) );
  NAND2_X1 U717 ( .A1(n645), .A2(n667), .ZN(n647) );
  XNOR2_X1 U718 ( .A(KEYINPUT110), .B(KEYINPUT63), .ZN(n646) );
  XNOR2_X1 U719 ( .A(n647), .B(n646), .ZN(G57) );
  XOR2_X1 U720 ( .A(n650), .B(n649), .Z(n653) );
  XNOR2_X1 U721 ( .A(n653), .B(KEYINPUT126), .ZN(n651) );
  XNOR2_X1 U722 ( .A(n741), .B(n651), .ZN(n652) );
  NAND2_X1 U723 ( .A1(n652), .A2(n434), .ZN(n657) );
  XOR2_X1 U724 ( .A(G227), .B(n653), .Z(n654) );
  NAND2_X1 U725 ( .A1(n654), .A2(G900), .ZN(n655) );
  NAND2_X1 U726 ( .A1(n655), .A2(G953), .ZN(n656) );
  NAND2_X1 U727 ( .A1(n657), .A2(n656), .ZN(G72) );
  BUF_X2 U728 ( .A(n751), .Z(n671) );
  NAND2_X1 U729 ( .A1(n671), .A2(G217), .ZN(n658) );
  XNOR2_X1 U730 ( .A(n369), .B(n658), .ZN(n660) );
  INV_X1 U731 ( .A(n667), .ZN(n756) );
  NOR2_X1 U732 ( .A1(n660), .A2(n756), .ZN(G66) );
  NAND2_X1 U733 ( .A1(n671), .A2(G478), .ZN(n662) );
  XNOR2_X1 U734 ( .A(n662), .B(n661), .ZN(n663) );
  NOR2_X1 U735 ( .A1(n663), .A2(n756), .ZN(G63) );
  NAND2_X1 U736 ( .A1(n751), .A2(G475), .ZN(n666) );
  XNOR2_X1 U737 ( .A(n666), .B(n665), .ZN(n668) );
  NAND2_X1 U738 ( .A1(n668), .A2(n667), .ZN(n670) );
  XOR2_X1 U739 ( .A(KEYINPUT68), .B(KEYINPUT60), .Z(n669) );
  XNOR2_X1 U740 ( .A(n670), .B(n669), .ZN(G60) );
  NAND2_X1 U741 ( .A1(n671), .A2(G469), .ZN(n676) );
  XNOR2_X1 U742 ( .A(KEYINPUT58), .B(KEYINPUT123), .ZN(n674) );
  XNOR2_X1 U743 ( .A(n672), .B(KEYINPUT57), .ZN(n673) );
  XNOR2_X1 U744 ( .A(n674), .B(n673), .ZN(n675) );
  XNOR2_X1 U745 ( .A(n676), .B(n675), .ZN(n677) );
  NOR2_X1 U746 ( .A1(n677), .A2(n756), .ZN(G54) );
  XNOR2_X1 U747 ( .A(n678), .B(G101), .ZN(n679) );
  XNOR2_X1 U748 ( .A(n679), .B(KEYINPUT111), .ZN(G3) );
  NAND2_X1 U749 ( .A1(n681), .A2(n691), .ZN(n680) );
  XNOR2_X1 U750 ( .A(n680), .B(G104), .ZN(G6) );
  XNOR2_X1 U751 ( .A(KEYINPUT27), .B(KEYINPUT112), .ZN(n685) );
  XOR2_X1 U752 ( .A(G107), .B(KEYINPUT26), .Z(n683) );
  NAND2_X1 U753 ( .A1(n681), .A2(n694), .ZN(n682) );
  XNOR2_X1 U754 ( .A(n683), .B(n682), .ZN(n684) );
  XNOR2_X1 U755 ( .A(n685), .B(n684), .ZN(G9) );
  XOR2_X1 U756 ( .A(KEYINPUT114), .B(KEYINPUT29), .Z(n687) );
  NAND2_X1 U757 ( .A1(n565), .A2(n694), .ZN(n686) );
  XNOR2_X1 U758 ( .A(n687), .B(n686), .ZN(n688) );
  XNOR2_X1 U759 ( .A(G128), .B(n688), .ZN(G30) );
  XOR2_X1 U760 ( .A(G146), .B(KEYINPUT115), .Z(n690) );
  NAND2_X1 U761 ( .A1(n565), .A2(n691), .ZN(n689) );
  XNOR2_X1 U762 ( .A(n690), .B(n689), .ZN(G48) );
  NAND2_X1 U763 ( .A1(n695), .A2(n691), .ZN(n692) );
  XNOR2_X1 U764 ( .A(n692), .B(KEYINPUT116), .ZN(n693) );
  XNOR2_X1 U765 ( .A(G113), .B(n693), .ZN(G15) );
  XOR2_X1 U766 ( .A(G116), .B(KEYINPUT117), .Z(n697) );
  NAND2_X1 U767 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U768 ( .A(n697), .B(n696), .ZN(G18) );
  XOR2_X1 U769 ( .A(KEYINPUT37), .B(KEYINPUT118), .Z(n698) );
  XNOR2_X1 U770 ( .A(n699), .B(n698), .ZN(n700) );
  XNOR2_X1 U771 ( .A(G125), .B(n700), .ZN(G27) );
  INV_X1 U772 ( .A(n701), .ZN(n703) );
  NAND2_X1 U773 ( .A1(n703), .A2(n387), .ZN(n704) );
  NAND2_X1 U774 ( .A1(n705), .A2(n704), .ZN(n709) );
  NAND2_X1 U775 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U776 ( .A1(n709), .A2(n708), .ZN(n711) );
  NAND2_X1 U777 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U778 ( .A(n712), .B(KEYINPUT120), .ZN(n728) );
  NOR2_X1 U779 ( .A1(n358), .A2(n714), .ZN(n715) );
  XNOR2_X1 U780 ( .A(n715), .B(KEYINPUT49), .ZN(n716) );
  NAND2_X1 U781 ( .A1(n717), .A2(n716), .ZN(n722) );
  NOR2_X1 U782 ( .A1(n719), .A2(n374), .ZN(n720) );
  XNOR2_X1 U783 ( .A(n720), .B(KEYINPUT50), .ZN(n721) );
  NOR2_X1 U784 ( .A1(n722), .A2(n721), .ZN(n723) );
  NOR2_X1 U785 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U786 ( .A(KEYINPUT51), .B(n725), .ZN(n726) );
  NAND2_X1 U787 ( .A1(n726), .A2(n733), .ZN(n727) );
  NAND2_X1 U788 ( .A1(n728), .A2(n727), .ZN(n729) );
  XOR2_X1 U789 ( .A(KEYINPUT52), .B(n729), .Z(n730) );
  NOR2_X1 U790 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U791 ( .A1(G952), .A2(n732), .ZN(n735) );
  NAND2_X1 U792 ( .A1(n733), .A2(n710), .ZN(n734) );
  NAND2_X1 U793 ( .A1(n735), .A2(n734), .ZN(n736) );
  XOR2_X1 U794 ( .A(KEYINPUT121), .B(n736), .Z(n749) );
  XOR2_X1 U795 ( .A(KEYINPUT2), .B(KEYINPUT84), .Z(n739) );
  AND2_X1 U796 ( .A1(n737), .A2(n739), .ZN(n738) );
  NOR2_X1 U797 ( .A1(n738), .A2(KEYINPUT87), .ZN(n745) );
  AND2_X1 U798 ( .A1(n739), .A2(KEYINPUT87), .ZN(n740) );
  NAND2_X1 U799 ( .A1(n741), .A2(n740), .ZN(n743) );
  NOR2_X1 U800 ( .A1(n743), .A2(n761), .ZN(n744) );
  NOR2_X1 U801 ( .A1(n745), .A2(n744), .ZN(n747) );
  NOR2_X1 U802 ( .A1(n747), .A2(n746), .ZN(n748) );
  INV_X1 U803 ( .A(KEYINPUT122), .ZN(n750) );
  XOR2_X1 U804 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n754) );
  BUF_X1 U805 ( .A(n752), .Z(n753) );
  XOR2_X1 U806 ( .A(n754), .B(n753), .Z(n755) );
  NOR2_X2 U807 ( .A1(n757), .A2(n756), .ZN(n759) );
  XNOR2_X1 U808 ( .A(KEYINPUT90), .B(KEYINPUT56), .ZN(n758) );
  XNOR2_X1 U809 ( .A(n759), .B(n758), .ZN(G51) );
  NAND2_X1 U810 ( .A1(n761), .A2(n760), .ZN(n766) );
  NAND2_X1 U811 ( .A1(G953), .A2(G224), .ZN(n762) );
  XNOR2_X1 U812 ( .A(KEYINPUT61), .B(n762), .ZN(n763) );
  NAND2_X1 U813 ( .A1(n763), .A2(G898), .ZN(n764) );
  XNOR2_X1 U814 ( .A(n764), .B(KEYINPUT124), .ZN(n765) );
  NAND2_X1 U815 ( .A1(n766), .A2(n765), .ZN(n773) );
  XOR2_X1 U816 ( .A(n768), .B(n767), .Z(n770) );
  NOR2_X1 U817 ( .A1(n770), .A2(n769), .ZN(n771) );
  XOR2_X1 U818 ( .A(KEYINPUT125), .B(n771), .Z(n772) );
  XNOR2_X1 U819 ( .A(n773), .B(n772), .ZN(G69) );
  XOR2_X1 U820 ( .A(n370), .B(G119), .Z(G21) );
  XNOR2_X1 U821 ( .A(G134), .B(n775), .ZN(G36) );
  XOR2_X1 U822 ( .A(G137), .B(n776), .Z(n777) );
  XNOR2_X1 U823 ( .A(KEYINPUT127), .B(n777), .ZN(G39) );
endmodule

