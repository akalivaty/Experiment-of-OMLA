//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 1 0 1 1 1 0 1 0 1 1 1 1 0 1 0 0 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 0 0 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:03 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  INV_X1    g0009(.A(G58), .ZN(new_n210));
  INV_X1    g0010(.A(G232), .ZN(new_n211));
  INV_X1    g0011(.A(G77), .ZN(new_n212));
  INV_X1    g0012(.A(G244), .ZN(new_n213));
  OAI22_X1  g0013(.A1(new_n210), .A2(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(G50), .ZN(new_n215));
  INV_X1    g0015(.A(G226), .ZN(new_n216));
  INV_X1    g0016(.A(G116), .ZN(new_n217));
  INV_X1    g0017(.A(G270), .ZN(new_n218));
  OAI22_X1  g0018(.A1(new_n215), .A2(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g0019(.A(KEYINPUT65), .B(G68), .ZN(new_n220));
  XNOR2_X1  g0020(.A(KEYINPUT66), .B(G238), .ZN(new_n221));
  AOI211_X1 g0021(.A(new_n214), .B(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G87), .ZN(new_n223));
  INV_X1    g0023(.A(G250), .ZN(new_n224));
  INV_X1    g0024(.A(G97), .ZN(new_n225));
  INV_X1    g0025(.A(G257), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  AND2_X1   g0027(.A1(G107), .A2(G264), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n206), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT1), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(G20), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT64), .ZN(new_n234));
  NOR2_X1   g0034(.A1(G58), .A2(G68), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g0036(.A1(new_n236), .A2(G50), .ZN(new_n237));
  INV_X1    g0037(.A(new_n237), .ZN(new_n238));
  AOI211_X1 g0038(.A(new_n209), .B(new_n230), .C1(new_n234), .C2(new_n238), .ZN(G361));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G226), .B(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G250), .B(G257), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G264), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(new_n218), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G358));
  XOR2_X1   g0048(.A(G68), .B(G77), .Z(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G58), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(G87), .B(G97), .Z(new_n252));
  XNOR2_X1  g0052(.A(G107), .B(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n251), .B(new_n254), .ZN(G351));
  INV_X1    g0055(.A(KEYINPUT71), .ZN(new_n256));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n231), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n204), .A2(G33), .ZN(new_n259));
  XNOR2_X1  g0059(.A(new_n259), .B(KEYINPUT70), .ZN(new_n260));
  NOR3_X1   g0060(.A1(new_n210), .A2(KEYINPUT69), .A3(KEYINPUT8), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT8), .B(G58), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n261), .B1(new_n262), .B2(KEYINPUT69), .ZN(new_n263));
  AND2_X1   g0063(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G150), .ZN(new_n265));
  NOR2_X1   g0065(.A1(G20), .A2(G33), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NOR3_X1   g0067(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n268));
  OAI22_X1  g0068(.A1(new_n265), .A2(new_n267), .B1(new_n268), .B2(new_n204), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n256), .B(new_n258), .C1(new_n264), .C2(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n269), .B1(new_n260), .B2(new_n263), .ZN(new_n271));
  INV_X1    g0071(.A(new_n258), .ZN(new_n272));
  OAI21_X1  g0072(.A(KEYINPUT71), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n275), .A2(G50), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n258), .B1(new_n203), .B2(G20), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G50), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n274), .A2(new_n277), .A3(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT3), .ZN(new_n282));
  INV_X1    g0082(.A(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(KEYINPUT3), .A2(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G1698), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G222), .ZN(new_n288));
  INV_X1    g0088(.A(G223), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n286), .B(new_n288), .C1(new_n289), .C2(new_n287), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n231), .B1(G33), .B2(G41), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n290), .B(new_n291), .C1(G77), .C2(new_n286), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(KEYINPUT68), .ZN(new_n294));
  NAND2_X1  g0094(.A1(G33), .A2(G41), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n295), .A2(G1), .A3(G13), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT68), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n297), .B(new_n203), .C1(G41), .C2(G45), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n294), .A2(G274), .A3(new_n296), .A4(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n296), .A2(new_n293), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n292), .B(new_n299), .C1(new_n216), .C2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G169), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n303), .B1(G179), .B2(new_n301), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n281), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n278), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n307), .A2(new_n212), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n275), .A2(G77), .ZN(new_n309));
  INV_X1    g0109(.A(new_n262), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n310), .A2(new_n266), .B1(G20), .B2(G77), .ZN(new_n311));
  XNOR2_X1  g0111(.A(KEYINPUT15), .B(G87), .ZN(new_n312));
  XNOR2_X1  g0112(.A(new_n312), .B(KEYINPUT72), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n311), .B1(new_n313), .B2(new_n259), .ZN(new_n314));
  AOI211_X1 g0114(.A(new_n308), .B(new_n309), .C1(new_n314), .C2(new_n258), .ZN(new_n315));
  INV_X1    g0115(.A(new_n299), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n221), .A2(G1698), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n317), .B(new_n286), .C1(new_n211), .C2(G1698), .ZN(new_n318));
  AND2_X1   g0118(.A1(KEYINPUT3), .A2(G33), .ZN(new_n319));
  NOR2_X1   g0119(.A1(KEYINPUT3), .A2(G33), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G107), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n296), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n316), .B1(new_n318), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n324), .B1(new_n213), .B2(new_n300), .ZN(new_n325));
  OR3_X1    g0125(.A1(new_n325), .A2(KEYINPUT73), .A3(G179), .ZN(new_n326));
  OAI21_X1  g0126(.A(KEYINPUT73), .B1(new_n325), .B2(G179), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n315), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n325), .A2(new_n302), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n280), .A2(KEYINPUT74), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT9), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT74), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n274), .A2(new_n333), .A3(new_n277), .A4(new_n279), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n331), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n301), .A2(G200), .ZN(new_n336));
  XOR2_X1   g0136(.A(new_n336), .B(KEYINPUT76), .Z(new_n337));
  INV_X1    g0137(.A(G190), .ZN(new_n338));
  OR2_X1    g0138(.A1(new_n301), .A2(new_n338), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n335), .A2(new_n337), .A3(KEYINPUT75), .A4(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n332), .B1(new_n331), .B2(new_n334), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT10), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NOR3_X1   g0144(.A1(new_n340), .A2(KEYINPUT10), .A3(new_n341), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n306), .B(new_n330), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n211), .A2(G1698), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n286), .B(new_n347), .C1(G226), .C2(G1698), .ZN(new_n348));
  NAND2_X1  g0148(.A1(G33), .A2(G97), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n296), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(G238), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n299), .B1(new_n351), .B2(new_n300), .ZN(new_n352));
  OR3_X1    g0152(.A1(new_n350), .A2(new_n352), .A3(KEYINPUT13), .ZN(new_n353));
  OAI21_X1  g0153(.A(KEYINPUT13), .B1(new_n350), .B2(new_n352), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(G169), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n356), .A2(KEYINPUT77), .A3(KEYINPUT14), .ZN(new_n357));
  OR2_X1    g0157(.A1(KEYINPUT77), .A2(KEYINPUT14), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n353), .A2(G179), .A3(new_n354), .ZN(new_n359));
  NAND2_X1  g0159(.A1(KEYINPUT77), .A2(KEYINPUT14), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n355), .A2(G169), .A3(new_n360), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n357), .A2(new_n358), .A3(new_n359), .A4(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n260), .A2(G77), .ZN(new_n363));
  INV_X1    g0163(.A(G68), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(KEYINPUT65), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT65), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(G68), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n368), .A2(G20), .B1(G50), .B2(new_n266), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n363), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n258), .ZN(new_n371));
  XOR2_X1   g0171(.A(new_n371), .B(KEYINPUT11), .Z(new_n372));
  INV_X1    g0172(.A(new_n275), .ZN(new_n373));
  AND3_X1   g0173(.A1(new_n368), .A2(new_n373), .A3(KEYINPUT12), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n307), .A2(KEYINPUT12), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n374), .B1(new_n375), .B2(G68), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n376), .B1(KEYINPUT12), .B2(new_n373), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n372), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n362), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n355), .A2(G200), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n378), .B(new_n381), .C1(new_n338), .C2(new_n355), .ZN(new_n382));
  AND2_X1   g0182(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT80), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n289), .A2(new_n287), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n216), .A2(G1698), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n385), .B(new_n386), .C1(new_n319), .C2(new_n320), .ZN(new_n387));
  NAND2_X1  g0187(.A1(G33), .A2(G87), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n291), .ZN(new_n390));
  INV_X1    g0190(.A(new_n300), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(G232), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n390), .A2(G179), .A3(new_n299), .A4(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n296), .B1(new_n387), .B2(new_n388), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n300), .A2(new_n211), .ZN(new_n395));
  NOR3_X1   g0195(.A1(new_n316), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n384), .B(new_n393), .C1(new_n396), .C2(new_n302), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n390), .A2(new_n299), .A3(new_n392), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(G169), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n384), .B1(new_n400), .B2(new_n393), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n263), .A2(new_n373), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n403), .B1(new_n307), .B2(new_n263), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n365), .A2(new_n367), .A3(G58), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n204), .B1(new_n405), .B2(new_n236), .ZN(new_n406));
  INV_X1    g0206(.A(G159), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n267), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(KEYINPUT78), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT78), .ZN(new_n410));
  INV_X1    g0210(.A(new_n408), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n235), .B1(new_n220), .B2(G58), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n410), .B(new_n411), .C1(new_n412), .C2(new_n204), .ZN(new_n413));
  AOI21_X1  g0213(.A(KEYINPUT7), .B1(new_n321), .B2(new_n204), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n284), .A2(KEYINPUT7), .A3(new_n204), .A4(new_n285), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(G68), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n409), .A2(new_n413), .A3(KEYINPUT16), .A4(new_n417), .ZN(new_n418));
  AND2_X1   g0218(.A1(new_n418), .A2(new_n258), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n220), .B1(new_n414), .B2(new_n416), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT79), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n406), .A2(new_n408), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n284), .A2(new_n204), .A3(new_n285), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT7), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n415), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n427), .A2(KEYINPUT79), .A3(new_n220), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n422), .A2(new_n423), .A3(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT16), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n404), .B1(new_n419), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(KEYINPUT81), .B1(new_n402), .B2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n404), .ZN(new_n434));
  AOI21_X1  g0234(.A(KEYINPUT79), .B1(new_n427), .B2(new_n220), .ZN(new_n435));
  AOI211_X1 g0235(.A(new_n421), .B(new_n368), .C1(new_n426), .C2(new_n415), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(KEYINPUT16), .B1(new_n437), .B2(new_n423), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n418), .A2(new_n258), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n434), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n400), .A2(new_n393), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(KEYINPUT80), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n397), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT81), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n440), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  AND3_X1   g0245(.A1(new_n433), .A2(KEYINPUT18), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(KEYINPUT18), .B1(new_n433), .B2(new_n445), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(G200), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n396), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  XNOR2_X1  g0251(.A(KEYINPUT82), .B(G190), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n396), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n432), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT83), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT17), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  AOI211_X1 g0257(.A(new_n404), .B(new_n450), .C1(new_n419), .C2(new_n431), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n455), .A2(new_n456), .ZN(new_n459));
  NAND2_X1  g0259(.A1(KEYINPUT83), .A2(KEYINPUT17), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n458), .A2(new_n459), .A3(new_n460), .A4(new_n453), .ZN(new_n461));
  AND2_X1   g0261(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n325), .A2(G200), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n463), .B(new_n315), .C1(new_n338), .C2(new_n325), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n383), .A2(new_n448), .A3(new_n462), .A4(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n346), .A2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n373), .A2(new_n322), .ZN(new_n468));
  XNOR2_X1  g0268(.A(new_n468), .B(KEYINPUT25), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n204), .B(G87), .C1(new_n319), .C2(new_n320), .ZN(new_n470));
  NAND2_X1  g0270(.A1(KEYINPUT94), .A2(KEYINPUT22), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n286), .A2(new_n204), .A3(G87), .A4(new_n471), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n204), .A2(G107), .ZN(new_n476));
  XNOR2_X1  g0276(.A(new_n476), .B(KEYINPUT23), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n283), .A2(new_n217), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n204), .ZN(new_n479));
  AND4_X1   g0279(.A1(KEYINPUT24), .A2(new_n475), .A3(new_n477), .A4(new_n479), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n473), .A2(new_n474), .B1(new_n204), .B2(new_n478), .ZN(new_n481));
  AOI21_X1  g0281(.A(KEYINPUT24), .B1(new_n481), .B2(new_n477), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n469), .B1(new_n483), .B2(new_n258), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n226), .A2(G1698), .ZN(new_n485));
  OAI221_X1 g0285(.A(new_n485), .B1(G250), .B2(G1698), .C1(new_n319), .C2(new_n320), .ZN(new_n486));
  NAND2_X1  g0286(.A1(G33), .A2(G294), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(KEYINPUT95), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT95), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n486), .A2(new_n490), .A3(new_n487), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n489), .A2(new_n291), .A3(new_n491), .ZN(new_n492));
  AND2_X1   g0292(.A1(KEYINPUT5), .A2(G41), .ZN(new_n493));
  NOR2_X1   g0293(.A1(KEYINPUT5), .A2(G41), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n203), .A2(G45), .A3(G274), .ZN(new_n496));
  OAI21_X1  g0296(.A(KEYINPUT85), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  XNOR2_X1  g0297(.A(KEYINPUT5), .B(G41), .ZN(new_n498));
  INV_X1    g0298(.A(new_n496), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT85), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n497), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n203), .A2(G45), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n498), .A2(new_n504), .B1(new_n232), .B2(new_n295), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(G264), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n492), .A2(new_n502), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(G200), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n492), .A2(G190), .A3(new_n502), .A4(new_n506), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n203), .A2(G33), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n275), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n511), .A2(new_n258), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(G107), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n484), .A2(new_n508), .A3(new_n509), .A4(new_n513), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n414), .A2(new_n416), .ZN(new_n515));
  OAI22_X1  g0315(.A1(new_n515), .A2(new_n322), .B1(new_n212), .B2(new_n267), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n225), .A2(new_n322), .A3(KEYINPUT6), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT84), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT6), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(G97), .ZN(new_n520));
  AND3_X1   g0320(.A1(new_n517), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n518), .B1(new_n517), .B2(new_n520), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n322), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NOR3_X1   g0323(.A1(new_n519), .A2(G97), .A3(G107), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n225), .A2(KEYINPUT6), .ZN(new_n525));
  OAI21_X1  g0325(.A(KEYINPUT84), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n517), .A2(new_n518), .A3(new_n520), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n526), .A2(new_n527), .A3(G107), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n204), .B1(new_n523), .B2(new_n528), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n258), .B1(new_n516), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n512), .A2(G97), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n373), .A2(new_n225), .ZN(new_n532));
  AND3_X1   g0332(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT4), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n534), .A2(G1698), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n535), .B(G244), .C1(new_n320), .C2(new_n319), .ZN(new_n536));
  NAND2_X1  g0336(.A1(G33), .A2(G283), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n213), .B1(new_n284), .B2(new_n285), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n536), .B(new_n537), .C1(new_n538), .C2(KEYINPUT4), .ZN(new_n539));
  OAI21_X1  g0339(.A(G250), .B1(new_n319), .B2(new_n320), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n287), .B1(new_n540), .B2(KEYINPUT4), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n291), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n505), .A2(G257), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n542), .A2(new_n543), .A3(new_n502), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(KEYINPUT86), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT86), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n542), .A2(new_n546), .A3(new_n543), .A4(new_n502), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n545), .A2(G200), .A3(new_n547), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n542), .A2(G190), .A3(new_n543), .A4(new_n502), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n533), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n551));
  INV_X1    g0351(.A(new_n544), .ZN(new_n552));
  INV_X1    g0352(.A(G179), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n544), .A2(new_n302), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n551), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT92), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n505), .A2(new_n557), .A3(G270), .ZN(new_n558));
  OAI211_X1 g0358(.A(G270), .B(new_n296), .C1(new_n495), .C2(new_n503), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(KEYINPUT92), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n287), .A2(G257), .ZN(new_n561));
  NAND2_X1  g0361(.A1(G264), .A2(G1698), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n561), .B(new_n562), .C1(new_n319), .C2(new_n320), .ZN(new_n563));
  INV_X1    g0363(.A(G303), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n284), .A2(new_n564), .A3(new_n285), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n563), .A2(new_n291), .A3(new_n565), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n558), .A2(new_n560), .A3(new_n502), .A4(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(KEYINPUT93), .ZN(new_n568));
  AND2_X1   g0368(.A1(new_n563), .A2(new_n565), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n569), .A2(new_n291), .B1(new_n501), .B2(new_n497), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT93), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n570), .A2(new_n571), .A3(new_n560), .A4(new_n558), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n452), .ZN(new_n574));
  NOR3_X1   g0374(.A1(new_n511), .A2(new_n217), .A3(new_n258), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n537), .B(new_n204), .C1(G33), .C2(new_n225), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n217), .A2(G20), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n576), .A2(new_n258), .A3(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT20), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n576), .A2(KEYINPUT20), .A3(new_n258), .A4(new_n577), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n575), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n373), .A2(new_n217), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n568), .A2(new_n572), .A3(G200), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n574), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n514), .A2(new_n550), .A3(new_n556), .A4(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n302), .B1(new_n582), .B2(new_n583), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n568), .A2(new_n572), .A3(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT21), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AND2_X1   g0392(.A1(new_n558), .A2(new_n560), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n584), .A2(new_n593), .A3(G179), .A4(new_n570), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n568), .A2(new_n572), .A3(new_n589), .A4(KEYINPUT21), .ZN(new_n595));
  AND3_X1   g0395(.A1(new_n592), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n204), .B(G68), .C1(new_n319), .C2(new_n320), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT89), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n286), .A2(KEYINPUT89), .A3(new_n204), .A4(G68), .ZN(new_n600));
  AND2_X1   g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n204), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT88), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n223), .A2(new_n225), .A3(new_n322), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n602), .A2(KEYINPUT88), .A3(new_n204), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT19), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n609), .B1(new_n259), .B2(new_n225), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n601), .A2(KEYINPUT90), .A3(new_n608), .A4(new_n610), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n608), .A2(new_n610), .A3(new_n599), .A4(new_n600), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT90), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n611), .A2(new_n258), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n313), .A2(new_n373), .ZN(new_n616));
  AND2_X1   g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n296), .A2(G250), .A3(new_n503), .ZN(new_n618));
  XNOR2_X1  g0418(.A(new_n496), .B(KEYINPUT87), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n284), .A2(new_n285), .B1(new_n351), .B2(new_n287), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n213), .A2(G1698), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n478), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n618), .B(new_n619), .C1(new_n622), .C2(new_n296), .ZN(new_n623));
  OR3_X1    g0423(.A1(new_n623), .A2(KEYINPUT91), .A3(new_n338), .ZN(new_n624));
  OAI21_X1  g0424(.A(KEYINPUT91), .B1(new_n623), .B2(new_n338), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n623), .A2(G200), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n512), .A2(G87), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n617), .A2(new_n626), .A3(new_n627), .A4(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n475), .A2(new_n477), .A3(new_n479), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT24), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n481), .A2(KEYINPUT24), .A3(new_n477), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n632), .A2(new_n258), .A3(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n469), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n634), .A2(new_n513), .A3(new_n635), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n492), .A2(new_n502), .A3(new_n506), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n553), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n507), .A2(new_n302), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n636), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n313), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n512), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n615), .A2(new_n616), .A3(new_n642), .ZN(new_n643));
  OAI221_X1 g0443(.A(new_n621), .B1(G238), .B2(G1698), .C1(new_n319), .C2(new_n320), .ZN(new_n644));
  INV_X1    g0444(.A(new_n478), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n296), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n619), .ZN(new_n647));
  INV_X1    g0447(.A(new_n618), .ZN(new_n648));
  NOR3_X1   g0448(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n553), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n623), .A2(new_n302), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n643), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n596), .A2(new_n629), .A3(new_n640), .A4(new_n652), .ZN(new_n653));
  NOR3_X1   g0453(.A1(new_n467), .A2(new_n588), .A3(new_n653), .ZN(G372));
  XNOR2_X1  g0454(.A(new_n342), .B(new_n343), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n380), .A2(new_n330), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n656), .A2(new_n382), .A3(new_n462), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT18), .ZN(new_n658));
  INV_X1    g0458(.A(new_n441), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n658), .B1(new_n432), .B2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n440), .A2(KEYINPUT18), .A3(new_n441), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n657), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n305), .B1(new_n655), .B2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n652), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n615), .A2(new_n627), .A3(new_n628), .A4(new_n616), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n666), .A2(KEYINPUT96), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(KEYINPUT96), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n626), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  AND4_X1   g0469(.A1(new_n509), .A2(new_n634), .A3(new_n513), .A4(new_n635), .ZN(new_n670));
  AND4_X1   g0470(.A1(new_n549), .A2(new_n530), .A3(new_n531), .A4(new_n532), .ZN(new_n671));
  AOI22_X1  g0471(.A1(new_n670), .A2(new_n508), .B1(new_n671), .B2(new_n548), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n640), .A2(new_n594), .A3(new_n595), .A4(new_n592), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n669), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT26), .ZN(new_n675));
  INV_X1    g0475(.A(new_n556), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n669), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n674), .A2(new_n675), .A3(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n676), .A2(new_n629), .A3(KEYINPUT26), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n665), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n664), .B1(new_n467), .B2(new_n680), .ZN(G369));
  NAND3_X1  g0481(.A1(new_n592), .A2(new_n594), .A3(new_n595), .ZN(new_n682));
  INV_X1    g0482(.A(G13), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n683), .A2(G20), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(new_n203), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n685), .A2(KEYINPUT27), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(KEYINPUT27), .ZN(new_n687));
  AND3_X1   g0487(.A1(new_n686), .A2(G213), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(G343), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n689), .B(KEYINPUT97), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(new_n585), .ZN(new_n691));
  XNOR2_X1  g0491(.A(new_n682), .B(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(new_n587), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(G330), .ZN(new_n695));
  INV_X1    g0495(.A(new_n690), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n640), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n636), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n514), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n697), .B1(new_n699), .B2(new_n640), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n596), .A2(new_n696), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n695), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n700), .A2(new_n701), .ZN(new_n704));
  INV_X1    g0504(.A(new_n697), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n703), .A2(new_n707), .ZN(G399));
  INV_X1    g0508(.A(new_n207), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(G41), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(G1), .ZN(new_n712));
  OR2_X1    g0512(.A1(new_n606), .A2(G116), .ZN(new_n713));
  OAI22_X1  g0513(.A1(new_n712), .A2(new_n713), .B1(new_n237), .B2(new_n711), .ZN(new_n714));
  XNOR2_X1  g0514(.A(new_n714), .B(KEYINPUT28), .ZN(new_n715));
  AND3_X1   g0515(.A1(new_n636), .A2(new_n639), .A3(new_n638), .ZN(new_n716));
  OAI211_X1 g0516(.A(new_n550), .B(new_n514), .C1(new_n716), .C2(new_n682), .ZN(new_n717));
  OR2_X1    g0517(.A1(new_n666), .A2(KEYINPUT96), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n666), .A2(KEYINPUT96), .ZN(new_n719));
  AOI22_X1  g0519(.A1(new_n718), .A2(new_n719), .B1(new_n624), .B2(new_n625), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n675), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(new_n556), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n556), .B1(new_n669), .B2(KEYINPUT26), .ZN(new_n723));
  OR2_X1    g0523(.A1(new_n629), .A2(KEYINPUT26), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n722), .A2(new_n652), .A3(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n726), .A2(KEYINPUT29), .A3(new_n690), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT29), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n728), .B1(new_n680), .B2(new_n696), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n653), .A2(new_n588), .A3(new_n696), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT30), .ZN(new_n732));
  AND2_X1   g0532(.A1(new_n497), .A2(new_n501), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n224), .B1(new_n284), .B2(new_n285), .ZN(new_n734));
  OAI21_X1  g0534(.A(G1698), .B1(new_n734), .B2(new_n534), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n534), .B1(new_n321), .B2(new_n213), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n735), .A2(new_n537), .A3(new_n736), .A4(new_n536), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n733), .B1(new_n737), .B2(new_n291), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n738), .A2(new_n543), .A3(new_n506), .A4(new_n492), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n649), .A2(new_n593), .A3(G179), .A4(new_n570), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n732), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NOR3_X1   g0541(.A1(new_n567), .A2(new_n623), .A3(new_n553), .ZN(new_n742));
  AND2_X1   g0542(.A1(new_n492), .A2(new_n506), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n742), .A2(new_n552), .A3(new_n743), .A4(KEYINPUT30), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n568), .A2(new_n572), .A3(new_n544), .A4(new_n623), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n746), .A2(new_n637), .A3(G179), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n696), .B1(new_n745), .B2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT31), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  XOR2_X1   g0550(.A(KEYINPUT98), .B(KEYINPUT31), .Z(new_n751));
  OAI211_X1 g0551(.A(new_n696), .B(new_n751), .C1(new_n745), .C2(new_n747), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(G330), .B1(new_n731), .B2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT99), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  OAI211_X1 g0556(.A(KEYINPUT99), .B(G330), .C1(new_n731), .C2(new_n753), .ZN(new_n757));
  AND2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n730), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g0559(.A(new_n759), .B(KEYINPUT100), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n715), .B1(new_n760), .B2(G1), .ZN(G364));
  OR2_X1    g0561(.A1(new_n694), .A2(G330), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n712), .B1(G45), .B2(new_n684), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n762), .A2(new_n695), .A3(new_n764), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT101), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n204), .B1(KEYINPUT102), .B2(new_n302), .ZN(new_n767));
  OR2_X1    g0567(.A1(new_n302), .A2(KEYINPUT102), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n231), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n204), .A2(new_n553), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n452), .A2(new_n449), .A3(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n452), .A2(G200), .A3(new_n771), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI22_X1  g0575(.A1(G322), .A2(new_n773), .B1(new_n775), .B2(G326), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n204), .A2(G190), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n777), .A2(G179), .A3(G200), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(G317), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(KEYINPUT33), .ZN(new_n781));
  OR2_X1    g0581(.A1(new_n780), .A2(KEYINPUT33), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n779), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(G294), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n338), .A2(G179), .A3(G200), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n204), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n776), .B(new_n783), .C1(new_n784), .C2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n777), .ZN(new_n788));
  NOR3_X1   g0588(.A1(new_n788), .A2(G179), .A3(G200), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n787), .B1(G329), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n449), .A2(G179), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n791), .A2(G20), .A3(G190), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n286), .B1(new_n793), .B2(G303), .ZN(new_n794));
  AND2_X1   g0594(.A1(new_n790), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(G283), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n791), .A2(new_n777), .ZN(new_n797));
  INV_X1    g0597(.A(G311), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n771), .A2(new_n338), .A3(new_n449), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n795), .B1(new_n796), .B2(new_n797), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n775), .A2(G50), .B1(G87), .B2(new_n793), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n801), .B1(new_n210), .B2(new_n772), .C1(new_n364), .C2(new_n778), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(new_n321), .ZN(new_n803));
  INV_X1    g0603(.A(new_n786), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(G97), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n789), .A2(G159), .ZN(new_n806));
  XOR2_X1   g0606(.A(new_n806), .B(KEYINPUT32), .Z(new_n807));
  INV_X1    g0607(.A(new_n799), .ZN(new_n808));
  INV_X1    g0608(.A(new_n797), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n808), .A2(G77), .B1(new_n809), .B2(G107), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n803), .A2(new_n805), .A3(new_n807), .A4(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n770), .B1(new_n800), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n709), .A2(new_n286), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(G45), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n814), .B1(new_n815), .B2(new_n238), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n816), .B1(new_n251), .B2(new_n815), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n207), .A2(G355), .A3(new_n286), .ZN(new_n818));
  OAI211_X1 g0618(.A(new_n817), .B(new_n818), .C1(G116), .C2(new_n207), .ZN(new_n819));
  NOR2_X1   g0619(.A1(G13), .A2(G33), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(G20), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n769), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n819), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n822), .ZN(new_n825));
  OAI211_X1 g0625(.A(new_n824), .B(new_n763), .C1(new_n694), .C2(new_n825), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n766), .B1(new_n812), .B2(new_n826), .ZN(G396));
  OAI21_X1  g0627(.A(new_n464), .B1(new_n315), .B2(new_n690), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n330), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n328), .A2(new_n329), .A3(new_n690), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n758), .B(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n680), .A2(new_n696), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n832), .B(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n834), .A2(new_n764), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n805), .B1(new_n217), .B2(new_n799), .C1(new_n564), .C2(new_n774), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(G294), .B2(new_n773), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n809), .A2(G87), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n789), .A2(G311), .B1(new_n793), .B2(G107), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n286), .B1(new_n779), .B2(G283), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n837), .A2(new_n838), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n773), .A2(G143), .B1(G150), .B2(new_n779), .ZN(new_n842));
  INV_X1    g0642(.A(G137), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n842), .B1(new_n843), .B2(new_n774), .C1(new_n407), .C2(new_n799), .ZN(new_n844));
  XOR2_X1   g0644(.A(new_n844), .B(KEYINPUT34), .Z(new_n845));
  AOI21_X1  g0645(.A(new_n845), .B1(G50), .B2(new_n793), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n809), .A2(G68), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n846), .B(new_n847), .C1(new_n210), .C2(new_n786), .ZN(new_n848));
  INV_X1    g0648(.A(new_n789), .ZN(new_n849));
  INV_X1    g0649(.A(G132), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n286), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n841), .B1(new_n848), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n769), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n769), .A2(new_n820), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(new_n212), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n831), .A2(new_n820), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n853), .A2(new_n763), .A3(new_n855), .A4(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n835), .A2(new_n857), .ZN(G384));
  NAND2_X1  g0658(.A1(new_n440), .A2(new_n688), .ZN(new_n859));
  AND2_X1   g0659(.A1(new_n454), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(KEYINPUT37), .B1(new_n440), .B2(new_n443), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n409), .A2(new_n413), .A3(new_n417), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n862), .A2(new_n430), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n434), .B1(new_n863), .B2(new_n439), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n688), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n441), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n454), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  AOI22_X1  g0667(.A1(new_n860), .A2(new_n861), .B1(new_n867), .B2(KEYINPUT37), .ZN(new_n868));
  AND3_X1   g0668(.A1(new_n440), .A2(new_n443), .A3(new_n444), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n444), .B1(new_n440), .B2(new_n443), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n658), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n433), .A2(KEYINPUT18), .A3(new_n445), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n871), .A2(new_n457), .A3(new_n461), .A4(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n865), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n868), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(KEYINPUT38), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n662), .A2(new_n457), .A3(new_n461), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n877), .A2(new_n440), .A3(new_n688), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n860), .A2(new_n861), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n454), .A2(new_n859), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n432), .A2(new_n659), .ZN(new_n881));
  OAI21_X1  g0681(.A(KEYINPUT37), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n878), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT38), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n876), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n588), .ZN(new_n888));
  NOR3_X1   g0688(.A1(new_n716), .A2(new_n665), .A3(new_n682), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n888), .A2(new_n889), .A3(new_n629), .A4(new_n690), .ZN(new_n890));
  INV_X1    g0690(.A(new_n751), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n748), .A2(new_n891), .ZN(new_n892));
  OR2_X1    g0692(.A1(new_n748), .A2(new_n749), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n890), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n379), .A2(new_n696), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n380), .A2(new_n382), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n362), .A2(new_n379), .A3(new_n696), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n831), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n894), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n887), .A2(KEYINPUT40), .A3(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n894), .A2(new_n898), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n865), .B1(new_n448), .B2(new_n462), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n885), .B1(new_n903), .B2(new_n868), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n902), .B1(new_n904), .B2(new_n876), .ZN(new_n905));
  OAI21_X1  g0705(.A(KEYINPUT104), .B1(new_n905), .B2(KEYINPUT40), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n875), .A2(KEYINPUT38), .ZN(new_n907));
  AOI211_X1 g0707(.A(new_n885), .B(new_n868), .C1(new_n873), .C2(new_n874), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n899), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT104), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT40), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n901), .B1(new_n906), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n913), .A2(new_n466), .A3(new_n894), .ZN(new_n914));
  NOR3_X1   g0714(.A1(new_n905), .A2(KEYINPUT104), .A3(KEYINPUT40), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n910), .B1(new_n909), .B2(new_n911), .ZN(new_n916));
  OAI211_X1 g0716(.A(G330), .B(new_n900), .C1(new_n915), .C2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n894), .A2(G330), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n466), .A2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n914), .B1(new_n918), .B2(new_n921), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n922), .B(KEYINPUT103), .Z(new_n923));
  NAND3_X1  g0723(.A1(new_n466), .A2(new_n727), .A3(new_n729), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n664), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n923), .B(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n904), .A2(KEYINPUT39), .A3(new_n876), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT39), .ZN(new_n928));
  AOI21_X1  g0728(.A(KEYINPUT38), .B1(new_n878), .B2(new_n883), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n928), .B1(new_n908), .B2(new_n929), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n380), .A2(new_n696), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AND2_X1   g0733(.A1(new_n678), .A2(new_n679), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n690), .B(new_n829), .C1(new_n934), .C2(new_n665), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n830), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n896), .A2(new_n897), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n936), .B(new_n937), .C1(new_n907), .C2(new_n908), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n662), .A2(new_n688), .ZN(new_n939));
  AND3_X1   g0739(.A1(new_n933), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n926), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n926), .A2(new_n940), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n941), .B(new_n942), .C1(new_n203), .C2(new_n684), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n523), .A2(new_n528), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n217), .B1(new_n944), .B2(KEYINPUT35), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n945), .B(new_n234), .C1(KEYINPUT35), .C2(new_n944), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT36), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n238), .A2(G77), .A3(new_n405), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(G50), .B2(new_n364), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n949), .A2(G1), .A3(new_n683), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n943), .A2(new_n947), .A3(new_n950), .ZN(G367));
  OAI211_X1 g0751(.A(new_n550), .B(new_n556), .C1(new_n533), .C2(new_n690), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n676), .A2(new_n696), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT106), .ZN(new_n955));
  OR3_X1    g0755(.A1(new_n703), .A2(KEYINPUT105), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(KEYINPUT105), .B1(new_n703), .B2(new_n955), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n617), .A2(new_n628), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n696), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n665), .B1(new_n669), .B2(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n961), .B1(new_n665), .B2(new_n960), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n962), .A2(KEYINPUT43), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n958), .B(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n556), .B1(new_n955), .B2(new_n640), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n690), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n704), .A2(new_n952), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT42), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n966), .A2(new_n968), .B1(KEYINPUT43), .B2(new_n962), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n964), .B(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n203), .B1(new_n684), .B2(G45), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  OR3_X1    g0772(.A1(new_n707), .A2(KEYINPUT44), .A3(new_n954), .ZN(new_n973));
  OAI21_X1  g0773(.A(KEYINPUT44), .B1(new_n707), .B2(new_n954), .ZN(new_n974));
  XOR2_X1   g0774(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n975));
  NAND3_X1  g0775(.A1(new_n707), .A2(new_n954), .A3(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n975), .ZN(new_n977));
  INV_X1    g0777(.A(new_n954), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n977), .B1(new_n706), .B2(new_n978), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n973), .A2(new_n974), .A3(new_n976), .A4(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n695), .A2(new_n702), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n703), .A2(new_n704), .A3(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n760), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n710), .B(KEYINPUT41), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n972), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n962), .A2(new_n825), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n823), .B1(new_n207), .B2(new_n313), .C1(new_n247), .C2(new_n814), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n849), .A2(new_n780), .ZN(new_n989));
  AOI21_X1  g0789(.A(KEYINPUT46), .B1(new_n793), .B2(G116), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n990), .A2(new_n286), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n808), .A2(G283), .B1(new_n809), .B2(G97), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n804), .A2(G107), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n793), .A2(KEYINPUT46), .A3(G116), .ZN(new_n994));
  NAND4_X1  g0794(.A1(new_n991), .A2(new_n992), .A3(new_n993), .A4(new_n994), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n989), .B(new_n995), .C1(G294), .C2(new_n779), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n996), .B1(new_n564), .B2(new_n772), .C1(new_n798), .C2(new_n774), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n997), .B(KEYINPUT108), .Z(new_n998));
  AOI22_X1  g0798(.A1(new_n775), .A2(G143), .B1(new_n804), .B2(G68), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n265), .B2(new_n772), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT109), .ZN(new_n1001));
  AND2_X1   g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n799), .A2(new_n215), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n286), .B1(new_n407), .B2(new_n778), .C1(new_n849), .C2(new_n843), .ZN(new_n1005));
  NOR4_X1   g0805(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n1006), .B1(new_n210), .B2(new_n792), .C1(new_n212), .C2(new_n797), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n998), .A2(new_n1007), .ZN(new_n1008));
  XOR2_X1   g0808(.A(KEYINPUT110), .B(KEYINPUT47), .Z(new_n1009));
  XOR2_X1   g0809(.A(new_n1008), .B(new_n1009), .Z(new_n1010));
  OAI211_X1 g0810(.A(new_n763), .B(new_n988), .C1(new_n1010), .C2(new_n770), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n970), .A2(new_n986), .B1(new_n987), .B2(new_n1011), .ZN(G387));
  INV_X1    g0812(.A(new_n983), .ZN(new_n1013));
  AND2_X1   g0813(.A1(new_n760), .A2(new_n1013), .ZN(new_n1014));
  OR3_X1    g0814(.A1(new_n1014), .A2(KEYINPUT112), .A3(new_n711), .ZN(new_n1015));
  OAI21_X1  g0815(.A(KEYINPUT112), .B1(new_n1014), .B2(new_n711), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n1015), .B(new_n1016), .C1(new_n760), .C2(new_n1013), .ZN(new_n1017));
  OR2_X1    g0817(.A1(new_n700), .A2(new_n825), .ZN(new_n1018));
  NOR3_X1   g0818(.A1(new_n262), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1019), .A2(new_n713), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(G68), .A2(G77), .ZN(new_n1021));
  OAI21_X1  g0821(.A(KEYINPUT50), .B1(new_n262), .B2(G50), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1020), .A2(new_n815), .A3(new_n1021), .A4(new_n1022), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n813), .B(new_n1023), .C1(new_n244), .C2(new_n815), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n207), .A2(new_n713), .A3(new_n286), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1024), .B(new_n1025), .C1(G107), .C2(new_n207), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT111), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(new_n823), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1018), .A2(new_n763), .A3(new_n1028), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n849), .A2(new_n265), .B1(new_n225), .B2(new_n797), .ZN(new_n1030));
  AOI211_X1 g0830(.A(new_n321), .B(new_n1030), .C1(G159), .C2(new_n775), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n793), .A2(G77), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1032), .B1(new_n364), .B2(new_n799), .C1(new_n215), .C2(new_n772), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n263), .A2(new_n779), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n641), .A2(new_n804), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1031), .A2(new_n1034), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n773), .A2(G317), .B1(G311), .B2(new_n779), .ZN(new_n1038));
  INV_X1    g0838(.A(G322), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1038), .B1(new_n564), .B2(new_n799), .C1(new_n1039), .C2(new_n774), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT48), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1041), .B1(new_n796), .B2(new_n786), .C1(new_n784), .C2(new_n792), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT49), .ZN(new_n1043));
  OR2_X1    g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n809), .A2(G116), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n789), .A2(G326), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n1044), .A2(new_n321), .A3(new_n1045), .A4(new_n1046), .ZN(new_n1047));
  AND2_X1   g0847(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1037), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1029), .B1(new_n1049), .B2(new_n769), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(new_n1013), .B2(new_n972), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1017), .A2(new_n1051), .ZN(G393));
  XNOR2_X1  g0852(.A(new_n980), .B(new_n703), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n823), .B1(new_n225), .B2(new_n207), .C1(new_n814), .C2(new_n254), .ZN(new_n1054));
  AND2_X1   g0854(.A1(new_n955), .A2(new_n822), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n799), .A2(new_n262), .B1(new_n792), .B2(new_n368), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n265), .A2(new_n774), .B1(new_n772), .B2(new_n407), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT51), .Z(new_n1058));
  AOI211_X1 g0858(.A(new_n1056), .B(new_n1058), .C1(G50), .C2(new_n779), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n804), .A2(G77), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n789), .A2(G143), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n321), .B1(new_n809), .B2(G87), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(G311), .A2(new_n773), .B1(new_n775), .B2(G317), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n1064), .A2(new_n1065), .B1(new_n784), .B2(new_n799), .ZN(new_n1066));
  AND2_X1   g0866(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n321), .B1(new_n786), .B2(new_n217), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n849), .A2(new_n1039), .B1(new_n322), .B2(new_n797), .ZN(new_n1069));
  NOR4_X1   g0869(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .A4(new_n1069), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1070), .B1(new_n796), .B2(new_n792), .C1(new_n564), .C2(new_n778), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n770), .B1(new_n1063), .B2(new_n1071), .ZN(new_n1072));
  NOR3_X1   g0872(.A1(new_n1055), .A2(new_n764), .A3(new_n1072), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n1053), .A2(new_n972), .B1(new_n1054), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1014), .A2(new_n980), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1075), .B1(new_n1053), .B2(new_n1014), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1074), .B1(new_n1076), .B2(new_n711), .ZN(G390));
  NAND2_X1  g0877(.A1(new_n919), .A2(new_n898), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n829), .ZN(new_n1080));
  NOR3_X1   g0880(.A1(new_n680), .A2(new_n696), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n830), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n937), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n932), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n1083), .A2(new_n1084), .B1(new_n930), .B2(new_n927), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n887), .A2(new_n1084), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n721), .A2(new_n556), .B1(new_n723), .B2(new_n724), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n696), .B1(new_n1087), .B2(new_n652), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n829), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n830), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1086), .B1(new_n1090), .B2(new_n937), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1079), .B1(new_n1085), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1082), .B1(new_n1088), .B2(new_n829), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n937), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1084), .B(new_n887), .C1(new_n1093), .C2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n831), .B1(new_n756), .B2(new_n757), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n937), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n932), .B1(new_n936), .B2(new_n937), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1095), .B(new_n1097), .C1(new_n1098), .C2(new_n931), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1092), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n924), .A2(new_n664), .A3(new_n920), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1078), .B1(new_n1096), .B2(new_n937), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n936), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n894), .A2(G330), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1094), .B1(new_n1104), .B2(new_n831), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1097), .A2(new_n1093), .A3(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1101), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1100), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1092), .A2(new_n1107), .A3(new_n1099), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1109), .A2(new_n710), .A3(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1092), .A2(new_n972), .A3(new_n1099), .ZN(new_n1112));
  OR2_X1    g0912(.A1(new_n931), .A2(new_n821), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n854), .ZN(new_n1114));
  OR2_X1    g0914(.A1(new_n1114), .A2(new_n263), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1060), .B1(new_n796), .B2(new_n774), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n849), .A2(new_n784), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n847), .B1(new_n223), .B2(new_n792), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n321), .B1(new_n778), .B2(new_n322), .ZN(new_n1119));
  NOR4_X1   g0919(.A1(new_n1116), .A2(new_n1117), .A3(new_n1118), .A4(new_n1119), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n1120), .B1(new_n225), .B2(new_n799), .C1(new_n217), .C2(new_n772), .ZN(new_n1121));
  OAI21_X1  g0921(.A(KEYINPUT53), .B1(new_n792), .B2(new_n265), .ZN(new_n1122));
  INV_X1    g0922(.A(G128), .ZN(new_n1123));
  XOR2_X1   g0923(.A(KEYINPUT54), .B(G143), .Z(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n1122), .B1(new_n774), .B2(new_n1123), .C1(new_n799), .C2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1126), .B1(G159), .B2(new_n804), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n789), .A2(G125), .ZN(new_n1128));
  NOR3_X1   g0928(.A1(new_n792), .A2(KEYINPUT53), .A3(new_n265), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(G137), .B2(new_n779), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n286), .B1(new_n797), .B2(new_n215), .ZN(new_n1131));
  XOR2_X1   g0931(.A(new_n1131), .B(KEYINPUT114), .Z(new_n1132));
  NAND4_X1  g0932(.A1(new_n1127), .A2(new_n1128), .A3(new_n1130), .A4(new_n1132), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n772), .A2(new_n850), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1121), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT115), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n769), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1113), .A2(new_n763), .A3(new_n1115), .A4(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1111), .A2(new_n1112), .A3(new_n1138), .ZN(G378));
  NAND3_X1  g0939(.A1(new_n933), .A2(new_n938), .A3(new_n939), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n331), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n334), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n688), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n655), .A2(new_n306), .ZN(new_n1145));
  XOR2_X1   g0945(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1146));
  AND2_X1   g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1144), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  OR2_X1    g0949(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1144), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1150), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  AND2_X1   g0953(.A1(new_n1149), .A2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n917), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1149), .A2(new_n1153), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(new_n913), .B2(G330), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1140), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n917), .A2(new_n1154), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n913), .A2(G330), .A3(new_n1156), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1159), .A2(new_n940), .A3(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1158), .A2(new_n972), .A3(new_n1161), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1114), .A2(G50), .ZN(new_n1163));
  INV_X1    g0963(.A(G41), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT118), .ZN(new_n1165));
  OR2_X1    g0965(.A1(new_n1165), .A2(G124), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(G124), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n789), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n775), .A2(G125), .B1(new_n804), .B2(G150), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT117), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n1170), .B1(new_n850), .B2(new_n778), .C1(new_n792), .C2(new_n1125), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(G137), .B2(new_n808), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1172), .B1(new_n1123), .B2(new_n772), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1164), .B(new_n1168), .C1(new_n1173), .C2(KEYINPUT59), .ZN(new_n1174));
  AOI211_X1 g0974(.A(G33), .B(new_n1174), .C1(G159), .C2(new_n809), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1173), .A2(KEYINPUT59), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n321), .B1(new_n313), .B2(new_n799), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n1032), .B1(new_n225), .B2(new_n778), .C1(new_n322), .C2(new_n772), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n1177), .B(new_n1178), .C1(G68), .C2(new_n804), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n809), .A2(G58), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n789), .A2(G283), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1179), .A2(new_n1164), .A3(new_n1180), .A4(new_n1181), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n774), .A2(new_n217), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n1175), .A2(new_n1176), .B1(KEYINPUT58), .B2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1184), .A2(KEYINPUT58), .ZN(new_n1186));
  AOI21_X1  g0986(.A(G50), .B1(new_n285), .B2(new_n1164), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  XOR2_X1   g0988(.A(new_n1188), .B(KEYINPUT116), .Z(new_n1189));
  AOI21_X1  g0989(.A(new_n770), .B1(new_n1185), .B2(new_n1189), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n1163), .B(new_n1190), .C1(new_n1156), .C2(new_n820), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1191), .A2(new_n763), .ZN(new_n1192));
  AND2_X1   g0992(.A1(new_n1162), .A2(new_n1192), .ZN(new_n1193));
  AND3_X1   g0993(.A1(new_n1159), .A2(new_n940), .A3(new_n1160), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n940), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1101), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1110), .A2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(KEYINPUT57), .B1(new_n1196), .B2(new_n1198), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1158), .A2(KEYINPUT57), .A3(new_n1198), .A4(new_n1161), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(new_n710), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1193), .B1(new_n1199), .B2(new_n1201), .ZN(G375));
  NAND3_X1  g1002(.A1(new_n1103), .A2(new_n1101), .A3(new_n1106), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1108), .A2(new_n985), .A3(new_n1203), .ZN(new_n1204));
  XOR2_X1   g1004(.A(new_n1204), .B(KEYINPUT119), .Z(new_n1205));
  NOR2_X1   g1005(.A1(new_n774), .A2(new_n784), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1036), .B1(new_n796), .B2(new_n772), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n1207), .B(KEYINPUT120), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n778), .A2(new_n217), .B1(new_n797), .B2(new_n212), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n286), .B(new_n1209), .C1(G107), .C2(new_n808), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n1208), .B(new_n1210), .C1(new_n564), .C2(new_n849), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n1206), .B(new_n1211), .C1(G97), .C2(new_n793), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n1180), .B1(new_n407), .B2(new_n792), .C1(new_n215), .C2(new_n786), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT121), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(new_n774), .B2(new_n850), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n775), .A2(KEYINPUT121), .A3(G132), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1213), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n779), .A2(new_n1124), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n773), .A2(G137), .B1(new_n789), .B2(G128), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1217), .A2(new_n286), .A3(new_n1218), .A4(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(G150), .B2(new_n808), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n769), .B1(new_n1212), .B2(new_n1221), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1222), .B(new_n763), .C1(new_n821), .C2(new_n937), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(new_n364), .B2(new_n854), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1224), .B1(new_n1225), .B2(new_n972), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1205), .A2(new_n1226), .ZN(G381));
  OR2_X1    g1027(.A1(G375), .A2(G378), .ZN(new_n1228));
  OR2_X1    g1028(.A1(new_n1228), .A2(G384), .ZN(new_n1229));
  OR2_X1    g1029(.A1(G390), .A2(G387), .ZN(new_n1230));
  INV_X1    g1030(.A(G396), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1017), .A2(new_n1231), .A3(new_n1051), .ZN(new_n1232));
  OR4_X1    g1032(.A1(G381), .A2(new_n1229), .A3(new_n1230), .A4(new_n1232), .ZN(G407));
  INV_X1    g1033(.A(G343), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(G213), .ZN(new_n1235));
  OAI21_X1  g1035(.A(KEYINPUT122), .B1(new_n1228), .B2(new_n1235), .ZN(new_n1236));
  OR3_X1    g1036(.A1(new_n1228), .A2(KEYINPUT122), .A3(new_n1235), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(G407), .A2(G213), .A3(new_n1236), .A4(new_n1237), .ZN(G409));
  NAND4_X1  g1038(.A1(new_n1158), .A2(new_n985), .A3(new_n1198), .A4(new_n1161), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1239), .A2(new_n1162), .A3(new_n1192), .ZN(new_n1240));
  AND3_X1   g1040(.A1(new_n1111), .A2(new_n1112), .A3(new_n1138), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(KEYINPUT123), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1193), .B(G378), .C1(new_n1199), .C2(new_n1201), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT123), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1240), .A2(new_n1241), .A3(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1243), .A2(new_n1244), .A3(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT60), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1203), .A2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(new_n1108), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT124), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  OR2_X1    g1052(.A1(new_n1203), .A2(new_n1248), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1249), .A2(new_n1108), .A3(KEYINPUT124), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1252), .A2(new_n710), .A3(new_n1253), .A4(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1255), .A2(G384), .A3(new_n1226), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(G384), .B1(new_n1255), .B2(new_n1226), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1247), .A2(new_n1235), .A3(new_n1259), .ZN(new_n1260));
  AND2_X1   g1060(.A1(new_n1260), .A2(KEYINPUT62), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(G390), .A2(G387), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1230), .A2(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1231), .B1(new_n1017), .B2(new_n1051), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1263), .A2(new_n1232), .A3(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1232), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n1230), .B(new_n1262), .C1(new_n1267), .C2(new_n1264), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1266), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1260), .A2(KEYINPUT62), .ZN(new_n1271));
  NOR3_X1   g1071(.A1(new_n1261), .A2(new_n1270), .A3(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1247), .A2(new_n1235), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1258), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1235), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1274), .A2(G2897), .A3(new_n1275), .A4(new_n1256), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(G2897), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1277), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1276), .A2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1273), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT61), .ZN(new_n1281));
  AOI21_X1  g1081(.A(KEYINPUT126), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(new_n1247), .A2(new_n1235), .B1(new_n1276), .B2(new_n1278), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT126), .ZN(new_n1284));
  NOR3_X1   g1084(.A1(new_n1283), .A2(new_n1284), .A3(KEYINPUT61), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1282), .A2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1260), .A2(KEYINPUT63), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT63), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1247), .A2(new_n1288), .A3(new_n1259), .A4(new_n1235), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1287), .A2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1273), .A2(KEYINPUT125), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT125), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1247), .A2(new_n1292), .A3(new_n1235), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1291), .A2(new_n1279), .A3(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1290), .A2(new_n1294), .A3(new_n1281), .ZN(new_n1295));
  AOI22_X1  g1095(.A1(new_n1272), .A2(new_n1286), .B1(new_n1295), .B2(new_n1270), .ZN(G405));
  NAND2_X1  g1096(.A1(new_n1259), .A2(KEYINPUT127), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(G375), .A2(new_n1241), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1297), .A2(new_n1244), .A3(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1270), .A2(new_n1299), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1269), .A2(new_n1244), .A3(new_n1298), .A4(new_n1297), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1259), .A2(KEYINPUT127), .ZN(new_n1302));
  AND3_X1   g1102(.A1(new_n1300), .A2(new_n1301), .A3(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1302), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1303), .A2(new_n1304), .ZN(G402));
endmodule


