

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U558 ( .A1(n578), .A2(n541), .ZN(n812) );
  OR2_X1 U559 ( .A1(n628), .A2(n779), .ZN(n626) );
  INV_X1 U560 ( .A(KEYINPUT64), .ZN(n611) );
  INV_X1 U561 ( .A(KEYINPUT29), .ZN(n641) );
  XNOR2_X1 U562 ( .A(n642), .B(n641), .ZN(n649) );
  AND2_X1 U563 ( .A1(n721), .A2(n723), .ZN(n644) );
  INV_X1 U564 ( .A(n644), .ZN(n663) );
  NOR2_X1 U565 ( .A1(G164), .A2(G1384), .ZN(n723) );
  NOR2_X1 U566 ( .A1(n604), .A2(n603), .ZN(n605) );
  NOR2_X2 U567 ( .A1(n523), .A2(G2105), .ZN(n883) );
  NAND2_X1 U568 ( .A1(n609), .A2(n608), .ZN(n999) );
  NOR2_X1 U569 ( .A1(n537), .A2(n536), .ZN(G160) );
  INV_X1 U570 ( .A(G2104), .ZN(n523) );
  NAND2_X1 U571 ( .A1(n883), .A2(G102), .ZN(n522) );
  XNOR2_X1 U572 ( .A(n522), .B(KEYINPUT86), .ZN(n525) );
  AND2_X1 U573 ( .A1(n523), .A2(G2105), .ZN(n880) );
  NAND2_X1 U574 ( .A1(G126), .A2(n880), .ZN(n524) );
  NAND2_X1 U575 ( .A1(n525), .A2(n524), .ZN(n530) );
  NOR2_X1 U576 ( .A1(G2104), .A2(G2105), .ZN(n526) );
  XOR2_X2 U577 ( .A(KEYINPUT17), .B(n526), .Z(n884) );
  NAND2_X1 U578 ( .A1(G138), .A2(n884), .ZN(n528) );
  AND2_X1 U579 ( .A1(G2104), .A2(G2105), .ZN(n879) );
  NAND2_X1 U580 ( .A1(G114), .A2(n879), .ZN(n527) );
  NAND2_X1 U581 ( .A1(n528), .A2(n527), .ZN(n529) );
  NOR2_X1 U582 ( .A1(n530), .A2(n529), .ZN(G164) );
  NAND2_X1 U583 ( .A1(n884), .A2(G137), .ZN(n533) );
  NAND2_X1 U584 ( .A1(G101), .A2(n883), .ZN(n531) );
  XOR2_X1 U585 ( .A(KEYINPUT23), .B(n531), .Z(n532) );
  NAND2_X1 U586 ( .A1(n533), .A2(n532), .ZN(n537) );
  NAND2_X1 U587 ( .A1(G113), .A2(n879), .ZN(n535) );
  NAND2_X1 U588 ( .A1(G125), .A2(n880), .ZN(n534) );
  NAND2_X1 U589 ( .A1(n535), .A2(n534), .ZN(n536) );
  NOR2_X1 U590 ( .A1(G651), .A2(G543), .ZN(n809) );
  NAND2_X1 U591 ( .A1(G91), .A2(n809), .ZN(n540) );
  INV_X1 U592 ( .A(G651), .ZN(n541) );
  NOR2_X1 U593 ( .A1(G543), .A2(n541), .ZN(n538) );
  XOR2_X1 U594 ( .A(KEYINPUT1), .B(n538), .Z(n804) );
  NAND2_X1 U595 ( .A1(G65), .A2(n804), .ZN(n539) );
  NAND2_X1 U596 ( .A1(n540), .A2(n539), .ZN(n546) );
  XOR2_X1 U597 ( .A(KEYINPUT0), .B(G543), .Z(n578) );
  NAND2_X1 U598 ( .A1(G78), .A2(n812), .ZN(n544) );
  NOR2_X1 U599 ( .A1(G651), .A2(n578), .ZN(n542) );
  XOR2_X2 U600 ( .A(KEYINPUT65), .B(n542), .Z(n805) );
  NAND2_X1 U601 ( .A1(G53), .A2(n805), .ZN(n543) );
  NAND2_X1 U602 ( .A1(n544), .A2(n543), .ZN(n545) );
  NOR2_X1 U603 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U604 ( .A(KEYINPUT68), .B(n547), .Z(G299) );
  NAND2_X1 U605 ( .A1(G64), .A2(n804), .ZN(n549) );
  NAND2_X1 U606 ( .A1(G52), .A2(n805), .ZN(n548) );
  NAND2_X1 U607 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U608 ( .A(KEYINPUT66), .B(n550), .ZN(n556) );
  NAND2_X1 U609 ( .A1(G90), .A2(n809), .ZN(n552) );
  NAND2_X1 U610 ( .A1(G77), .A2(n812), .ZN(n551) );
  NAND2_X1 U611 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U612 ( .A(KEYINPUT9), .B(n553), .ZN(n554) );
  XNOR2_X1 U613 ( .A(KEYINPUT67), .B(n554), .ZN(n555) );
  NOR2_X1 U614 ( .A1(n556), .A2(n555), .ZN(G171) );
  NAND2_X1 U615 ( .A1(n809), .A2(G89), .ZN(n557) );
  XNOR2_X1 U616 ( .A(n557), .B(KEYINPUT4), .ZN(n559) );
  NAND2_X1 U617 ( .A1(G76), .A2(n812), .ZN(n558) );
  NAND2_X1 U618 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U619 ( .A(n560), .B(KEYINPUT5), .ZN(n566) );
  NAND2_X1 U620 ( .A1(n804), .A2(G63), .ZN(n561) );
  XOR2_X1 U621 ( .A(KEYINPUT75), .B(n561), .Z(n563) );
  NAND2_X1 U622 ( .A1(n805), .A2(G51), .ZN(n562) );
  NAND2_X1 U623 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U624 ( .A(KEYINPUT6), .B(n564), .Z(n565) );
  NAND2_X1 U625 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U626 ( .A(n567), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U627 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U628 ( .A1(G75), .A2(n812), .ZN(n569) );
  NAND2_X1 U629 ( .A1(G62), .A2(n804), .ZN(n568) );
  NAND2_X1 U630 ( .A1(n569), .A2(n568), .ZN(n572) );
  NAND2_X1 U631 ( .A1(n809), .A2(G88), .ZN(n570) );
  XOR2_X1 U632 ( .A(KEYINPUT82), .B(n570), .Z(n571) );
  NOR2_X1 U633 ( .A1(n572), .A2(n571), .ZN(n574) );
  NAND2_X1 U634 ( .A1(n805), .A2(G50), .ZN(n573) );
  NAND2_X1 U635 ( .A1(n574), .A2(n573), .ZN(G303) );
  NAND2_X1 U636 ( .A1(G49), .A2(n805), .ZN(n576) );
  NAND2_X1 U637 ( .A1(G74), .A2(G651), .ZN(n575) );
  NAND2_X1 U638 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U639 ( .A1(n804), .A2(n577), .ZN(n580) );
  NAND2_X1 U640 ( .A1(n578), .A2(G87), .ZN(n579) );
  NAND2_X1 U641 ( .A1(n580), .A2(n579), .ZN(G288) );
  NAND2_X1 U642 ( .A1(G73), .A2(n812), .ZN(n581) );
  XNOR2_X1 U643 ( .A(n581), .B(KEYINPUT2), .ZN(n588) );
  NAND2_X1 U644 ( .A1(G86), .A2(n809), .ZN(n583) );
  NAND2_X1 U645 ( .A1(G48), .A2(n805), .ZN(n582) );
  NAND2_X1 U646 ( .A1(n583), .A2(n582), .ZN(n586) );
  NAND2_X1 U647 ( .A1(G61), .A2(n804), .ZN(n584) );
  XNOR2_X1 U648 ( .A(KEYINPUT81), .B(n584), .ZN(n585) );
  NOR2_X1 U649 ( .A1(n586), .A2(n585), .ZN(n587) );
  NAND2_X1 U650 ( .A1(n588), .A2(n587), .ZN(G305) );
  NAND2_X1 U651 ( .A1(G85), .A2(n809), .ZN(n590) );
  NAND2_X1 U652 ( .A1(G60), .A2(n804), .ZN(n589) );
  NAND2_X1 U653 ( .A1(n590), .A2(n589), .ZN(n594) );
  NAND2_X1 U654 ( .A1(G72), .A2(n812), .ZN(n592) );
  NAND2_X1 U655 ( .A1(G47), .A2(n805), .ZN(n591) );
  NAND2_X1 U656 ( .A1(n592), .A2(n591), .ZN(n593) );
  OR2_X1 U657 ( .A1(n594), .A2(n593), .ZN(G290) );
  AND2_X1 U658 ( .A1(G160), .A2(G40), .ZN(n721) );
  AND2_X1 U659 ( .A1(G1996), .A2(n723), .ZN(n595) );
  AND2_X1 U660 ( .A1(n721), .A2(n595), .ZN(n596) );
  XOR2_X1 U661 ( .A(n596), .B(KEYINPUT26), .Z(n598) );
  NAND2_X1 U662 ( .A1(n663), .A2(G1341), .ZN(n597) );
  NAND2_X1 U663 ( .A1(n598), .A2(n597), .ZN(n610) );
  NAND2_X1 U664 ( .A1(G56), .A2(n804), .ZN(n599) );
  XOR2_X1 U665 ( .A(KEYINPUT14), .B(n599), .Z(n607) );
  XOR2_X1 U666 ( .A(KEYINPUT12), .B(KEYINPUT70), .Z(n601) );
  NAND2_X1 U667 ( .A1(G81), .A2(n809), .ZN(n600) );
  XNOR2_X1 U668 ( .A(n601), .B(n600), .ZN(n604) );
  NAND2_X1 U669 ( .A1(n812), .A2(G68), .ZN(n602) );
  XNOR2_X1 U670 ( .A(KEYINPUT71), .B(n602), .ZN(n603) );
  XNOR2_X1 U671 ( .A(n605), .B(KEYINPUT13), .ZN(n606) );
  NOR2_X1 U672 ( .A1(n607), .A2(n606), .ZN(n609) );
  NAND2_X1 U673 ( .A1(n805), .A2(G43), .ZN(n608) );
  NOR2_X1 U674 ( .A1(n610), .A2(n999), .ZN(n612) );
  XNOR2_X1 U675 ( .A(n612), .B(n611), .ZN(n628) );
  NAND2_X1 U676 ( .A1(G66), .A2(n804), .ZN(n619) );
  NAND2_X1 U677 ( .A1(G92), .A2(n809), .ZN(n614) );
  NAND2_X1 U678 ( .A1(G79), .A2(n812), .ZN(n613) );
  NAND2_X1 U679 ( .A1(n614), .A2(n613), .ZN(n617) );
  NAND2_X1 U680 ( .A1(n805), .A2(G54), .ZN(n615) );
  XOR2_X1 U681 ( .A(n615), .B(KEYINPUT74), .Z(n616) );
  NOR2_X1 U682 ( .A1(n617), .A2(n616), .ZN(n618) );
  NAND2_X1 U683 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X2 U684 ( .A(n620), .B(KEYINPUT15), .ZN(n1000) );
  INV_X1 U685 ( .A(n1000), .ZN(n779) );
  NAND2_X1 U686 ( .A1(G1348), .A2(n663), .ZN(n621) );
  XNOR2_X1 U687 ( .A(n621), .B(KEYINPUT94), .ZN(n623) );
  NAND2_X1 U688 ( .A1(G2067), .A2(n644), .ZN(n622) );
  NAND2_X1 U689 ( .A1(n623), .A2(n622), .ZN(n624) );
  XOR2_X1 U690 ( .A(KEYINPUT95), .B(n624), .Z(n625) );
  NAND2_X1 U691 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X1 U692 ( .A(n627), .B(KEYINPUT96), .ZN(n630) );
  NAND2_X1 U693 ( .A1(n628), .A2(n779), .ZN(n629) );
  NAND2_X1 U694 ( .A1(n630), .A2(n629), .ZN(n636) );
  NAND2_X1 U695 ( .A1(G1956), .A2(n663), .ZN(n631) );
  XNOR2_X1 U696 ( .A(KEYINPUT93), .B(n631), .ZN(n634) );
  NAND2_X1 U697 ( .A1(n644), .A2(G2072), .ZN(n632) );
  XNOR2_X1 U698 ( .A(KEYINPUT27), .B(n632), .ZN(n633) );
  NOR2_X1 U699 ( .A1(n634), .A2(n633), .ZN(n637) );
  INV_X1 U700 ( .A(G299), .ZN(n1005) );
  NAND2_X1 U701 ( .A1(n637), .A2(n1005), .ZN(n635) );
  NAND2_X1 U702 ( .A1(n636), .A2(n635), .ZN(n640) );
  NOR2_X1 U703 ( .A1(n637), .A2(n1005), .ZN(n638) );
  XOR2_X1 U704 ( .A(n638), .B(KEYINPUT28), .Z(n639) );
  NAND2_X1 U705 ( .A1(n640), .A2(n639), .ZN(n642) );
  XOR2_X1 U706 ( .A(KEYINPUT25), .B(G2078), .Z(n952) );
  NOR2_X1 U707 ( .A1(n952), .A2(n663), .ZN(n643) );
  XOR2_X1 U708 ( .A(KEYINPUT92), .B(n643), .Z(n647) );
  NOR2_X1 U709 ( .A1(n644), .A2(G1961), .ZN(n645) );
  XNOR2_X1 U710 ( .A(KEYINPUT91), .B(n645), .ZN(n646) );
  NAND2_X1 U711 ( .A1(n647), .A2(n646), .ZN(n652) );
  NAND2_X1 U712 ( .A1(G171), .A2(n652), .ZN(n648) );
  NAND2_X1 U713 ( .A1(n649), .A2(n648), .ZN(n651) );
  INV_X1 U714 ( .A(KEYINPUT97), .ZN(n650) );
  XNOR2_X1 U715 ( .A(n651), .B(n650), .ZN(n661) );
  NOR2_X1 U716 ( .A1(G171), .A2(n652), .ZN(n657) );
  NAND2_X1 U717 ( .A1(G8), .A2(n663), .ZN(n701) );
  NOR2_X1 U718 ( .A1(G1966), .A2(n701), .ZN(n674) );
  NOR2_X1 U719 ( .A1(G2084), .A2(n663), .ZN(n675) );
  NOR2_X1 U720 ( .A1(n674), .A2(n675), .ZN(n653) );
  NAND2_X1 U721 ( .A1(G8), .A2(n653), .ZN(n654) );
  XNOR2_X1 U722 ( .A(KEYINPUT30), .B(n654), .ZN(n655) );
  NOR2_X1 U723 ( .A1(G168), .A2(n655), .ZN(n656) );
  NOR2_X1 U724 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U725 ( .A(KEYINPUT31), .B(n658), .ZN(n659) );
  XOR2_X1 U726 ( .A(KEYINPUT98), .B(n659), .Z(n660) );
  NAND2_X1 U727 ( .A1(n661), .A2(n660), .ZN(n672) );
  NAND2_X1 U728 ( .A1(n672), .A2(G286), .ZN(n662) );
  XNOR2_X1 U729 ( .A(n662), .B(KEYINPUT100), .ZN(n669) );
  NOR2_X1 U730 ( .A1(G1971), .A2(n701), .ZN(n665) );
  NOR2_X1 U731 ( .A1(G2090), .A2(n663), .ZN(n664) );
  NOR2_X1 U732 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U733 ( .A1(n666), .A2(G303), .ZN(n667) );
  XOR2_X1 U734 ( .A(KEYINPUT101), .B(n667), .Z(n668) );
  NAND2_X1 U735 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U736 ( .A1(n670), .A2(G8), .ZN(n671) );
  XNOR2_X1 U737 ( .A(n671), .B(KEYINPUT32), .ZN(n680) );
  INV_X1 U738 ( .A(n672), .ZN(n673) );
  NOR2_X1 U739 ( .A1(n674), .A2(n673), .ZN(n677) );
  NAND2_X1 U740 ( .A1(G8), .A2(n675), .ZN(n676) );
  NAND2_X1 U741 ( .A1(n677), .A2(n676), .ZN(n678) );
  XOR2_X1 U742 ( .A(KEYINPUT99), .B(n678), .Z(n679) );
  NAND2_X1 U743 ( .A1(n680), .A2(n679), .ZN(n696) );
  NOR2_X1 U744 ( .A1(G2090), .A2(G303), .ZN(n681) );
  NAND2_X1 U745 ( .A1(G8), .A2(n681), .ZN(n682) );
  NAND2_X1 U746 ( .A1(n696), .A2(n682), .ZN(n683) );
  NAND2_X1 U747 ( .A1(n683), .A2(n701), .ZN(n708) );
  NOR2_X1 U748 ( .A1(G1976), .A2(G288), .ZN(n688) );
  NOR2_X1 U749 ( .A1(G1971), .A2(G303), .ZN(n684) );
  NOR2_X1 U750 ( .A1(n688), .A2(n684), .ZN(n1004) );
  XNOR2_X1 U751 ( .A(n1004), .B(KEYINPUT102), .ZN(n687) );
  NOR2_X1 U752 ( .A1(G1981), .A2(G305), .ZN(n685) );
  XNOR2_X1 U753 ( .A(KEYINPUT24), .B(n685), .ZN(n700) );
  INV_X1 U754 ( .A(n700), .ZN(n686) );
  AND2_X1 U755 ( .A1(n687), .A2(n686), .ZN(n694) );
  XNOR2_X1 U756 ( .A(KEYINPUT103), .B(n688), .ZN(n689) );
  NOR2_X1 U757 ( .A1(n701), .A2(n689), .ZN(n692) );
  XOR2_X1 U758 ( .A(KEYINPUT104), .B(G1981), .Z(n690) );
  XNOR2_X1 U759 ( .A(G305), .B(n690), .ZN(n1015) );
  NAND2_X1 U760 ( .A1(n1015), .A2(KEYINPUT33), .ZN(n691) );
  NOR2_X1 U761 ( .A1(n692), .A2(n691), .ZN(n704) );
  INV_X1 U762 ( .A(n704), .ZN(n693) );
  AND2_X1 U763 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U764 ( .A1(n696), .A2(n695), .ZN(n706) );
  NAND2_X1 U765 ( .A1(G1976), .A2(G288), .ZN(n1003) );
  AND2_X1 U766 ( .A1(n1003), .A2(n1015), .ZN(n698) );
  NOR2_X1 U767 ( .A1(KEYINPUT103), .A2(KEYINPUT33), .ZN(n697) );
  AND2_X1 U768 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U769 ( .A1(n700), .A2(n699), .ZN(n702) );
  NOR2_X1 U770 ( .A1(n702), .A2(n701), .ZN(n703) );
  OR2_X1 U771 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U772 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U773 ( .A1(n708), .A2(n707), .ZN(n710) );
  INV_X1 U774 ( .A(KEYINPUT105), .ZN(n709) );
  XNOR2_X1 U775 ( .A(n710), .B(n709), .ZN(n747) );
  XOR2_X1 U776 ( .A(G2067), .B(KEYINPUT37), .Z(n748) );
  NAND2_X1 U777 ( .A1(G116), .A2(n879), .ZN(n712) );
  NAND2_X1 U778 ( .A1(G128), .A2(n880), .ZN(n711) );
  NAND2_X1 U779 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U780 ( .A(n713), .B(KEYINPUT35), .ZN(n718) );
  NAND2_X1 U781 ( .A1(G104), .A2(n883), .ZN(n715) );
  NAND2_X1 U782 ( .A1(G140), .A2(n884), .ZN(n714) );
  NAND2_X1 U783 ( .A1(n715), .A2(n714), .ZN(n716) );
  XOR2_X1 U784 ( .A(KEYINPUT34), .B(n716), .Z(n717) );
  NAND2_X1 U785 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U786 ( .A(n719), .B(KEYINPUT36), .ZN(n892) );
  NAND2_X1 U787 ( .A1(n748), .A2(n892), .ZN(n720) );
  XNOR2_X1 U788 ( .A(n720), .B(KEYINPUT88), .ZN(n941) );
  INV_X1 U789 ( .A(n721), .ZN(n722) );
  NOR2_X1 U790 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U791 ( .A(KEYINPUT87), .B(n724), .Z(n761) );
  INV_X1 U792 ( .A(n761), .ZN(n725) );
  NOR2_X1 U793 ( .A1(n941), .A2(n725), .ZN(n757) );
  INV_X1 U794 ( .A(n757), .ZN(n743) );
  NAND2_X1 U795 ( .A1(G105), .A2(n883), .ZN(n726) );
  XNOR2_X1 U796 ( .A(n726), .B(KEYINPUT38), .ZN(n733) );
  NAND2_X1 U797 ( .A1(G141), .A2(n884), .ZN(n728) );
  NAND2_X1 U798 ( .A1(G117), .A2(n879), .ZN(n727) );
  NAND2_X1 U799 ( .A1(n728), .A2(n727), .ZN(n731) );
  NAND2_X1 U800 ( .A1(n880), .A2(G129), .ZN(n729) );
  XOR2_X1 U801 ( .A(KEYINPUT90), .B(n729), .Z(n730) );
  NOR2_X1 U802 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U803 ( .A1(n733), .A2(n732), .ZN(n864) );
  NAND2_X1 U804 ( .A1(G1996), .A2(n864), .ZN(n742) );
  NAND2_X1 U805 ( .A1(G95), .A2(n883), .ZN(n735) );
  NAND2_X1 U806 ( .A1(G119), .A2(n880), .ZN(n734) );
  NAND2_X1 U807 ( .A1(n735), .A2(n734), .ZN(n738) );
  NAND2_X1 U808 ( .A1(G131), .A2(n884), .ZN(n736) );
  XNOR2_X1 U809 ( .A(KEYINPUT89), .B(n736), .ZN(n737) );
  NOR2_X1 U810 ( .A1(n738), .A2(n737), .ZN(n740) );
  NAND2_X1 U811 ( .A1(n879), .A2(G107), .ZN(n739) );
  NAND2_X1 U812 ( .A1(n740), .A2(n739), .ZN(n876) );
  NAND2_X1 U813 ( .A1(G1991), .A2(n876), .ZN(n741) );
  NAND2_X1 U814 ( .A1(n742), .A2(n741), .ZN(n933) );
  NAND2_X1 U815 ( .A1(n761), .A2(n933), .ZN(n751) );
  NAND2_X1 U816 ( .A1(n743), .A2(n751), .ZN(n745) );
  XNOR2_X1 U817 ( .A(G1986), .B(G290), .ZN(n1014) );
  AND2_X1 U818 ( .A1(n1014), .A2(n761), .ZN(n744) );
  NOR2_X1 U819 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U820 ( .A1(n747), .A2(n746), .ZN(n764) );
  NOR2_X1 U821 ( .A1(n892), .A2(n748), .ZN(n926) );
  NOR2_X1 U822 ( .A1(G1986), .A2(G290), .ZN(n749) );
  NOR2_X1 U823 ( .A1(G1991), .A2(n876), .ZN(n928) );
  NOR2_X1 U824 ( .A1(n749), .A2(n928), .ZN(n750) );
  XNOR2_X1 U825 ( .A(KEYINPUT107), .B(n750), .ZN(n752) );
  NAND2_X1 U826 ( .A1(n752), .A2(n751), .ZN(n754) );
  NOR2_X1 U827 ( .A1(G1996), .A2(n864), .ZN(n753) );
  XOR2_X1 U828 ( .A(KEYINPUT106), .B(n753), .Z(n922) );
  NAND2_X1 U829 ( .A1(n754), .A2(n922), .ZN(n755) );
  XNOR2_X1 U830 ( .A(KEYINPUT39), .B(n755), .ZN(n756) );
  NOR2_X1 U831 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U832 ( .A(n758), .B(KEYINPUT108), .ZN(n759) );
  NOR2_X1 U833 ( .A1(n926), .A2(n759), .ZN(n760) );
  XNOR2_X1 U834 ( .A(KEYINPUT109), .B(n760), .ZN(n762) );
  NAND2_X1 U835 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U836 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U837 ( .A(n765), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U838 ( .A(G2451), .B(G2454), .Z(n767) );
  XNOR2_X1 U839 ( .A(G2430), .B(KEYINPUT110), .ZN(n766) );
  XNOR2_X1 U840 ( .A(n767), .B(n766), .ZN(n768) );
  XOR2_X1 U841 ( .A(n768), .B(G2446), .Z(n770) );
  XNOR2_X1 U842 ( .A(G1341), .B(G1348), .ZN(n769) );
  XNOR2_X1 U843 ( .A(n770), .B(n769), .ZN(n774) );
  XOR2_X1 U844 ( .A(G2438), .B(G2427), .Z(n772) );
  XNOR2_X1 U845 ( .A(G2443), .B(G2435), .ZN(n771) );
  XNOR2_X1 U846 ( .A(n772), .B(n771), .ZN(n773) );
  XOR2_X1 U847 ( .A(n774), .B(n773), .Z(n775) );
  AND2_X1 U848 ( .A1(G14), .A2(n775), .ZN(G401) );
  AND2_X1 U849 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U850 ( .A(G57), .ZN(G237) );
  INV_X1 U851 ( .A(G82), .ZN(G220) );
  NAND2_X1 U852 ( .A1(G7), .A2(G661), .ZN(n776) );
  XNOR2_X1 U853 ( .A(n776), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U854 ( .A(G223), .ZN(n837) );
  NAND2_X1 U855 ( .A1(n837), .A2(G567), .ZN(n777) );
  XOR2_X1 U856 ( .A(KEYINPUT11), .B(n777), .Z(G234) );
  INV_X1 U857 ( .A(G860), .ZN(n784) );
  NOR2_X1 U858 ( .A1(n999), .A2(n784), .ZN(n778) );
  XOR2_X1 U859 ( .A(KEYINPUT72), .B(n778), .Z(G153) );
  XNOR2_X1 U860 ( .A(G171), .B(KEYINPUT73), .ZN(G301) );
  NAND2_X1 U861 ( .A1(G868), .A2(G301), .ZN(n781) );
  INV_X1 U862 ( .A(G868), .ZN(n821) );
  NAND2_X1 U863 ( .A1(n779), .A2(n821), .ZN(n780) );
  NAND2_X1 U864 ( .A1(n781), .A2(n780), .ZN(G284) );
  NOR2_X1 U865 ( .A1(G286), .A2(n821), .ZN(n783) );
  NOR2_X1 U866 ( .A1(G299), .A2(G868), .ZN(n782) );
  NOR2_X1 U867 ( .A1(n783), .A2(n782), .ZN(G297) );
  NAND2_X1 U868 ( .A1(n784), .A2(G559), .ZN(n785) );
  NAND2_X1 U869 ( .A1(n785), .A2(n1000), .ZN(n786) );
  XNOR2_X1 U870 ( .A(n786), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U871 ( .A1(G868), .A2(n999), .ZN(n789) );
  NAND2_X1 U872 ( .A1(G868), .A2(n1000), .ZN(n787) );
  NOR2_X1 U873 ( .A1(G559), .A2(n787), .ZN(n788) );
  NOR2_X1 U874 ( .A1(n789), .A2(n788), .ZN(G282) );
  XOR2_X1 U875 ( .A(G2100), .B(KEYINPUT76), .Z(n798) );
  NAND2_X1 U876 ( .A1(G123), .A2(n880), .ZN(n790) );
  XNOR2_X1 U877 ( .A(n790), .B(KEYINPUT18), .ZN(n792) );
  NAND2_X1 U878 ( .A1(n883), .A2(G99), .ZN(n791) );
  NAND2_X1 U879 ( .A1(n792), .A2(n791), .ZN(n796) );
  NAND2_X1 U880 ( .A1(G135), .A2(n884), .ZN(n794) );
  NAND2_X1 U881 ( .A1(G111), .A2(n879), .ZN(n793) );
  NAND2_X1 U882 ( .A1(n794), .A2(n793), .ZN(n795) );
  NOR2_X1 U883 ( .A1(n796), .A2(n795), .ZN(n927) );
  XNOR2_X1 U884 ( .A(G2096), .B(n927), .ZN(n797) );
  NAND2_X1 U885 ( .A1(n798), .A2(n797), .ZN(G156) );
  XNOR2_X1 U886 ( .A(KEYINPUT83), .B(KEYINPUT19), .ZN(n800) );
  XNOR2_X1 U887 ( .A(G305), .B(KEYINPUT84), .ZN(n799) );
  XNOR2_X1 U888 ( .A(n800), .B(n799), .ZN(n803) );
  XNOR2_X1 U889 ( .A(G299), .B(G303), .ZN(n801) );
  XNOR2_X1 U890 ( .A(n801), .B(G290), .ZN(n802) );
  XNOR2_X1 U891 ( .A(n803), .B(n802), .ZN(n818) );
  NAND2_X1 U892 ( .A1(G67), .A2(n804), .ZN(n807) );
  NAND2_X1 U893 ( .A1(G55), .A2(n805), .ZN(n806) );
  NAND2_X1 U894 ( .A1(n807), .A2(n806), .ZN(n808) );
  XNOR2_X1 U895 ( .A(n808), .B(KEYINPUT79), .ZN(n811) );
  NAND2_X1 U896 ( .A1(G93), .A2(n809), .ZN(n810) );
  NAND2_X1 U897 ( .A1(n811), .A2(n810), .ZN(n815) );
  NAND2_X1 U898 ( .A1(n812), .A2(G80), .ZN(n813) );
  XOR2_X1 U899 ( .A(KEYINPUT78), .B(n813), .Z(n814) );
  NOR2_X1 U900 ( .A1(n815), .A2(n814), .ZN(n816) );
  XOR2_X1 U901 ( .A(KEYINPUT80), .B(n816), .Z(n844) );
  XNOR2_X1 U902 ( .A(G288), .B(n844), .ZN(n817) );
  XNOR2_X1 U903 ( .A(n818), .B(n817), .ZN(n850) );
  NAND2_X1 U904 ( .A1(G559), .A2(n1000), .ZN(n819) );
  XOR2_X1 U905 ( .A(n999), .B(n819), .Z(n841) );
  XOR2_X1 U906 ( .A(n850), .B(n841), .Z(n820) );
  NOR2_X1 U907 ( .A1(n821), .A2(n820), .ZN(n823) );
  NOR2_X1 U908 ( .A1(n844), .A2(G868), .ZN(n822) );
  NOR2_X1 U909 ( .A1(n823), .A2(n822), .ZN(G295) );
  NAND2_X1 U910 ( .A1(G2084), .A2(G2078), .ZN(n824) );
  XOR2_X1 U911 ( .A(KEYINPUT20), .B(n824), .Z(n825) );
  NAND2_X1 U912 ( .A1(G2090), .A2(n825), .ZN(n826) );
  XNOR2_X1 U913 ( .A(KEYINPUT21), .B(n826), .ZN(n827) );
  NAND2_X1 U914 ( .A1(n827), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U915 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U916 ( .A(KEYINPUT69), .B(G132), .ZN(G219) );
  NOR2_X1 U917 ( .A1(G220), .A2(G219), .ZN(n828) );
  XOR2_X1 U918 ( .A(KEYINPUT22), .B(n828), .Z(n829) );
  NOR2_X1 U919 ( .A1(G218), .A2(n829), .ZN(n830) );
  NAND2_X1 U920 ( .A1(G96), .A2(n830), .ZN(n845) );
  NAND2_X1 U921 ( .A1(n845), .A2(G2106), .ZN(n834) );
  NAND2_X1 U922 ( .A1(G69), .A2(G120), .ZN(n831) );
  NOR2_X1 U923 ( .A1(G237), .A2(n831), .ZN(n832) );
  NAND2_X1 U924 ( .A1(G108), .A2(n832), .ZN(n846) );
  NAND2_X1 U925 ( .A1(n846), .A2(G567), .ZN(n833) );
  NAND2_X1 U926 ( .A1(n834), .A2(n833), .ZN(n921) );
  NAND2_X1 U927 ( .A1(G661), .A2(G483), .ZN(n835) );
  NOR2_X1 U928 ( .A1(n921), .A2(n835), .ZN(n840) );
  NAND2_X1 U929 ( .A1(G36), .A2(n840), .ZN(n836) );
  XOR2_X1 U930 ( .A(KEYINPUT85), .B(n836), .Z(G176) );
  INV_X1 U931 ( .A(G303), .ZN(G166) );
  NAND2_X1 U932 ( .A1(G2106), .A2(n837), .ZN(G217) );
  AND2_X1 U933 ( .A1(G15), .A2(G2), .ZN(n838) );
  NAND2_X1 U934 ( .A1(G661), .A2(n838), .ZN(G259) );
  NAND2_X1 U935 ( .A1(G3), .A2(G1), .ZN(n839) );
  NAND2_X1 U936 ( .A1(n840), .A2(n839), .ZN(G188) );
  XNOR2_X1 U938 ( .A(KEYINPUT77), .B(n841), .ZN(n842) );
  NOR2_X1 U939 ( .A1(G860), .A2(n842), .ZN(n843) );
  XOR2_X1 U940 ( .A(n844), .B(n843), .Z(G145) );
  INV_X1 U941 ( .A(G120), .ZN(G236) );
  INV_X1 U942 ( .A(G96), .ZN(G221) );
  INV_X1 U943 ( .A(G69), .ZN(G235) );
  NOR2_X1 U944 ( .A1(n846), .A2(n845), .ZN(G325) );
  INV_X1 U945 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U946 ( .A(n999), .B(G286), .ZN(n848) );
  XNOR2_X1 U947 ( .A(G171), .B(n1000), .ZN(n847) );
  XNOR2_X1 U948 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U949 ( .A(n850), .B(n849), .Z(n851) );
  NOR2_X1 U950 ( .A1(G37), .A2(n851), .ZN(G397) );
  NAND2_X1 U951 ( .A1(G124), .A2(n880), .ZN(n852) );
  XOR2_X1 U952 ( .A(KEYINPUT111), .B(n852), .Z(n853) );
  XNOR2_X1 U953 ( .A(n853), .B(KEYINPUT44), .ZN(n855) );
  NAND2_X1 U954 ( .A1(G136), .A2(n884), .ZN(n854) );
  NAND2_X1 U955 ( .A1(n855), .A2(n854), .ZN(n856) );
  XNOR2_X1 U956 ( .A(KEYINPUT112), .B(n856), .ZN(n860) );
  NAND2_X1 U957 ( .A1(G100), .A2(n883), .ZN(n858) );
  NAND2_X1 U958 ( .A1(G112), .A2(n879), .ZN(n857) );
  NAND2_X1 U959 ( .A1(n858), .A2(n857), .ZN(n859) );
  NOR2_X1 U960 ( .A1(n860), .A2(n859), .ZN(G162) );
  XOR2_X1 U961 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n862) );
  XNOR2_X1 U962 ( .A(G164), .B(KEYINPUT115), .ZN(n861) );
  XNOR2_X1 U963 ( .A(n862), .B(n861), .ZN(n866) );
  XOR2_X1 U964 ( .A(G160), .B(n927), .Z(n863) );
  XNOR2_X1 U965 ( .A(n864), .B(n863), .ZN(n865) );
  XNOR2_X1 U966 ( .A(n866), .B(n865), .ZN(n878) );
  NAND2_X1 U967 ( .A1(G103), .A2(n883), .ZN(n868) );
  NAND2_X1 U968 ( .A1(G139), .A2(n884), .ZN(n867) );
  NAND2_X1 U969 ( .A1(n868), .A2(n867), .ZN(n874) );
  NAND2_X1 U970 ( .A1(n880), .A2(G127), .ZN(n869) );
  XOR2_X1 U971 ( .A(KEYINPUT113), .B(n869), .Z(n871) );
  NAND2_X1 U972 ( .A1(n879), .A2(G115), .ZN(n870) );
  NAND2_X1 U973 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U974 ( .A(KEYINPUT47), .B(n872), .Z(n873) );
  NOR2_X1 U975 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U976 ( .A(KEYINPUT114), .B(n875), .Z(n937) );
  XNOR2_X1 U977 ( .A(n876), .B(n937), .ZN(n877) );
  XNOR2_X1 U978 ( .A(n878), .B(n877), .ZN(n891) );
  NAND2_X1 U979 ( .A1(G118), .A2(n879), .ZN(n882) );
  NAND2_X1 U980 ( .A1(G130), .A2(n880), .ZN(n881) );
  NAND2_X1 U981 ( .A1(n882), .A2(n881), .ZN(n889) );
  NAND2_X1 U982 ( .A1(G106), .A2(n883), .ZN(n886) );
  NAND2_X1 U983 ( .A1(G142), .A2(n884), .ZN(n885) );
  NAND2_X1 U984 ( .A1(n886), .A2(n885), .ZN(n887) );
  XOR2_X1 U985 ( .A(KEYINPUT45), .B(n887), .Z(n888) );
  NOR2_X1 U986 ( .A1(n889), .A2(n888), .ZN(n890) );
  XOR2_X1 U987 ( .A(n891), .B(n890), .Z(n894) );
  XNOR2_X1 U988 ( .A(n892), .B(G162), .ZN(n893) );
  XNOR2_X1 U989 ( .A(n894), .B(n893), .ZN(n895) );
  NOR2_X1 U990 ( .A1(n895), .A2(G37), .ZN(n896) );
  XNOR2_X1 U991 ( .A(n896), .B(KEYINPUT116), .ZN(G395) );
  XOR2_X1 U992 ( .A(G2096), .B(G2100), .Z(n898) );
  XNOR2_X1 U993 ( .A(KEYINPUT42), .B(G2678), .ZN(n897) );
  XNOR2_X1 U994 ( .A(n898), .B(n897), .ZN(n902) );
  XOR2_X1 U995 ( .A(KEYINPUT43), .B(G2090), .Z(n900) );
  XNOR2_X1 U996 ( .A(G2067), .B(G2072), .ZN(n899) );
  XNOR2_X1 U997 ( .A(n900), .B(n899), .ZN(n901) );
  XOR2_X1 U998 ( .A(n902), .B(n901), .Z(n904) );
  XNOR2_X1 U999 ( .A(G2084), .B(G2078), .ZN(n903) );
  XNOR2_X1 U1000 ( .A(n904), .B(n903), .ZN(G227) );
  XOR2_X1 U1001 ( .A(G1981), .B(G1971), .Z(n906) );
  XNOR2_X1 U1002 ( .A(G1966), .B(G1956), .ZN(n905) );
  XNOR2_X1 U1003 ( .A(n906), .B(n905), .ZN(n907) );
  XOR2_X1 U1004 ( .A(n907), .B(KEYINPUT41), .Z(n909) );
  XNOR2_X1 U1005 ( .A(G1976), .B(G1986), .ZN(n908) );
  XNOR2_X1 U1006 ( .A(n909), .B(n908), .ZN(n913) );
  XOR2_X1 U1007 ( .A(G2474), .B(G1991), .Z(n911) );
  XNOR2_X1 U1008 ( .A(G1961), .B(G1996), .ZN(n910) );
  XNOR2_X1 U1009 ( .A(n911), .B(n910), .ZN(n912) );
  XNOR2_X1 U1010 ( .A(n913), .B(n912), .ZN(G229) );
  NOR2_X1 U1011 ( .A1(G397), .A2(G395), .ZN(n914) );
  XNOR2_X1 U1012 ( .A(KEYINPUT118), .B(n914), .ZN(n920) );
  NOR2_X1 U1013 ( .A1(n921), .A2(G401), .ZN(n915) );
  XNOR2_X1 U1014 ( .A(n915), .B(KEYINPUT117), .ZN(n918) );
  NOR2_X1 U1015 ( .A1(G227), .A2(G229), .ZN(n916) );
  XNOR2_X1 U1016 ( .A(KEYINPUT49), .B(n916), .ZN(n917) );
  NOR2_X1 U1017 ( .A1(n918), .A2(n917), .ZN(n919) );
  NAND2_X1 U1018 ( .A1(n920), .A2(n919), .ZN(G225) );
  INV_X1 U1019 ( .A(G225), .ZN(G308) );
  INV_X1 U1020 ( .A(n921), .ZN(G319) );
  INV_X1 U1021 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1022 ( .A(G2090), .B(G162), .ZN(n923) );
  NAND2_X1 U1023 ( .A1(n923), .A2(n922), .ZN(n924) );
  XNOR2_X1 U1024 ( .A(n924), .B(KEYINPUT51), .ZN(n935) );
  XOR2_X1 U1025 ( .A(G2084), .B(G160), .Z(n925) );
  NOR2_X1 U1026 ( .A1(n926), .A2(n925), .ZN(n931) );
  NOR2_X1 U1027 ( .A1(n928), .A2(n927), .ZN(n929) );
  XOR2_X1 U1028 ( .A(KEYINPUT119), .B(n929), .Z(n930) );
  NAND2_X1 U1029 ( .A1(n931), .A2(n930), .ZN(n932) );
  NOR2_X1 U1030 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(n944) );
  XOR2_X1 U1032 ( .A(G164), .B(G2078), .Z(n936) );
  XNOR2_X1 U1033 ( .A(KEYINPUT120), .B(n936), .ZN(n939) );
  XNOR2_X1 U1034 ( .A(n937), .B(G2072), .ZN(n938) );
  NOR2_X1 U1035 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1036 ( .A(KEYINPUT50), .B(n940), .ZN(n942) );
  NAND2_X1 U1037 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1038 ( .A1(n944), .A2(n943), .ZN(n945) );
  XOR2_X1 U1039 ( .A(KEYINPUT52), .B(n945), .Z(n946) );
  NOR2_X1 U1040 ( .A1(KEYINPUT55), .A2(n946), .ZN(n947) );
  XNOR2_X1 U1041 ( .A(KEYINPUT121), .B(n947), .ZN(n948) );
  NAND2_X1 U1042 ( .A1(n948), .A2(G29), .ZN(n998) );
  XOR2_X1 U1043 ( .A(G1991), .B(G25), .Z(n949) );
  NAND2_X1 U1044 ( .A1(n949), .A2(G28), .ZN(n958) );
  XNOR2_X1 U1045 ( .A(G1996), .B(G32), .ZN(n951) );
  XNOR2_X1 U1046 ( .A(G33), .B(G2072), .ZN(n950) );
  NOR2_X1 U1047 ( .A1(n951), .A2(n950), .ZN(n956) );
  XNOR2_X1 U1048 ( .A(n952), .B(G27), .ZN(n954) );
  XNOR2_X1 U1049 ( .A(G2067), .B(G26), .ZN(n953) );
  NOR2_X1 U1050 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n957) );
  NOR2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1053 ( .A(KEYINPUT53), .B(n959), .Z(n962) );
  XOR2_X1 U1054 ( .A(KEYINPUT54), .B(G34), .Z(n960) );
  XNOR2_X1 U1055 ( .A(G2084), .B(n960), .ZN(n961) );
  NAND2_X1 U1056 ( .A1(n962), .A2(n961), .ZN(n964) );
  XNOR2_X1 U1057 ( .A(G35), .B(G2090), .ZN(n963) );
  NOR2_X1 U1058 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1059 ( .A(KEYINPUT55), .B(n965), .ZN(n967) );
  INV_X1 U1060 ( .A(G29), .ZN(n966) );
  NAND2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1062 ( .A1(n968), .A2(G11), .ZN(n969) );
  XNOR2_X1 U1063 ( .A(n969), .B(KEYINPUT122), .ZN(n996) );
  XOR2_X1 U1064 ( .A(KEYINPUT61), .B(KEYINPUT127), .Z(n993) );
  XOR2_X1 U1065 ( .A(G1961), .B(G5), .Z(n981) );
  XOR2_X1 U1066 ( .A(G4), .B(KEYINPUT125), .Z(n971) );
  XNOR2_X1 U1067 ( .A(G1348), .B(KEYINPUT59), .ZN(n970) );
  XNOR2_X1 U1068 ( .A(n971), .B(n970), .ZN(n975) );
  XNOR2_X1 U1069 ( .A(G1341), .B(G19), .ZN(n973) );
  XNOR2_X1 U1070 ( .A(G6), .B(G1981), .ZN(n972) );
  NOR2_X1 U1071 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1072 ( .A1(n975), .A2(n974), .ZN(n978) );
  XNOR2_X1 U1073 ( .A(KEYINPUT124), .B(G1956), .ZN(n976) );
  XNOR2_X1 U1074 ( .A(G20), .B(n976), .ZN(n977) );
  NOR2_X1 U1075 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1076 ( .A(KEYINPUT60), .B(n979), .ZN(n980) );
  NAND2_X1 U1077 ( .A1(n981), .A2(n980), .ZN(n988) );
  XNOR2_X1 U1078 ( .A(G1971), .B(G22), .ZN(n983) );
  XNOR2_X1 U1079 ( .A(G23), .B(G1976), .ZN(n982) );
  NOR2_X1 U1080 ( .A1(n983), .A2(n982), .ZN(n985) );
  XOR2_X1 U1081 ( .A(G1986), .B(G24), .Z(n984) );
  NAND2_X1 U1082 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1083 ( .A(KEYINPUT58), .B(n986), .ZN(n987) );
  NOR2_X1 U1084 ( .A1(n988), .A2(n987), .ZN(n991) );
  XOR2_X1 U1085 ( .A(G1966), .B(KEYINPUT126), .Z(n989) );
  XNOR2_X1 U1086 ( .A(G21), .B(n989), .ZN(n990) );
  NAND2_X1 U1087 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1088 ( .A(n993), .B(n992), .ZN(n994) );
  NOR2_X1 U1089 ( .A1(G16), .A2(n994), .ZN(n995) );
  NOR2_X1 U1090 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1091 ( .A1(n998), .A2(n997), .ZN(n1025) );
  XOR2_X1 U1092 ( .A(G16), .B(KEYINPUT56), .Z(n1023) );
  XNOR2_X1 U1093 ( .A(G1341), .B(n999), .ZN(n1002) );
  XOR2_X1 U1094 ( .A(G1348), .B(n1000), .Z(n1001) );
  NOR2_X1 U1095 ( .A1(n1002), .A2(n1001), .ZN(n1012) );
  NAND2_X1 U1096 ( .A1(n1004), .A2(n1003), .ZN(n1009) );
  XNOR2_X1 U1097 ( .A(n1005), .B(G1956), .ZN(n1007) );
  NAND2_X1 U1098 ( .A1(G1971), .A2(G303), .ZN(n1006) );
  NAND2_X1 U1099 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1100 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1101 ( .A(KEYINPUT123), .B(n1010), .Z(n1011) );
  NAND2_X1 U1102 ( .A1(n1012), .A2(n1011), .ZN(n1021) );
  XOR2_X1 U1103 ( .A(G171), .B(G1961), .Z(n1013) );
  NOR2_X1 U1104 ( .A1(n1014), .A2(n1013), .ZN(n1019) );
  XNOR2_X1 U1105 ( .A(G1966), .B(G168), .ZN(n1016) );
  NAND2_X1 U1106 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1107 ( .A(n1017), .B(KEYINPUT57), .ZN(n1018) );
  NAND2_X1 U1108 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NOR2_X1 U1109 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NOR2_X1 U1110 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1111 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1112 ( .A(n1026), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1113 ( .A(G311), .ZN(G150) );
endmodule

