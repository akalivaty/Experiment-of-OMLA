//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 1 1 0 1 0 0 1 0 0 0 1 1 1 1 0 0 1 1 1 1 0 1 1 1 1 1 0 1 0 1 0 0 0 1 1 0 0 1 1 1 0 0 1 1 1 1 1 1 1 0 1 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:39 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(G125), .B(G140), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT16), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT16), .ZN(new_n192));
  INV_X1    g006(.A(G140), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(new_n193), .A3(G125), .ZN(new_n194));
  AND3_X1   g008(.A1(new_n191), .A2(G146), .A3(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT23), .ZN(new_n197));
  INV_X1    g011(.A(G119), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n197), .B1(new_n198), .B2(G128), .ZN(new_n199));
  INV_X1    g013(.A(G128), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n200), .A2(KEYINPUT23), .A3(G119), .ZN(new_n201));
  OAI211_X1 g015(.A(new_n199), .B(new_n201), .C1(G119), .C2(new_n200), .ZN(new_n202));
  XNOR2_X1  g016(.A(G119), .B(G128), .ZN(new_n203));
  XOR2_X1   g017(.A(KEYINPUT24), .B(G110), .Z(new_n204));
  OAI22_X1  g018(.A1(new_n202), .A2(G110), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n193), .A2(G125), .ZN(new_n206));
  INV_X1    g020(.A(G125), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G140), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n196), .B(new_n205), .C1(G146), .C2(new_n209), .ZN(new_n210));
  AOI22_X1  g024(.A1(new_n202), .A2(G110), .B1(new_n203), .B2(new_n204), .ZN(new_n211));
  AOI21_X1  g025(.A(G146), .B1(new_n191), .B2(new_n194), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n211), .B1(new_n195), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G953), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(G221), .A3(G234), .ZN(new_n216));
  XNOR2_X1  g030(.A(new_n216), .B(KEYINPUT78), .ZN(new_n217));
  XNOR2_X1  g031(.A(KEYINPUT22), .B(G137), .ZN(new_n218));
  XNOR2_X1  g032(.A(new_n217), .B(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(new_n214), .B(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(KEYINPUT25), .B1(new_n221), .B2(new_n188), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n214), .A2(new_n220), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n219), .B1(new_n210), .B2(new_n213), .ZN(new_n224));
  OAI211_X1 g038(.A(KEYINPUT25), .B(new_n188), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n189), .B1(new_n222), .B2(new_n226), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n189), .A2(G902), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n221), .A2(new_n228), .ZN(new_n229));
  AND2_X1   g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT77), .ZN(new_n232));
  INV_X1    g046(.A(G472), .ZN(new_n233));
  INV_X1    g047(.A(G146), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G143), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(KEYINPUT1), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G128), .ZN(new_n237));
  INV_X1    g051(.A(G143), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G146), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n235), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT66), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n242), .B1(new_n238), .B2(G146), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n234), .A2(KEYINPUT66), .A3(G143), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n200), .A2(KEYINPUT1), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n243), .A2(new_n244), .A3(new_n245), .A4(new_n239), .ZN(new_n246));
  AND2_X1   g060(.A1(new_n246), .A2(KEYINPUT68), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n246), .A2(KEYINPUT68), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n241), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G134), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G137), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n250), .A2(G137), .ZN(new_n253));
  OAI21_X1  g067(.A(G131), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT11), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n255), .B1(new_n250), .B2(G137), .ZN(new_n256));
  INV_X1    g070(.A(G137), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n257), .A2(KEYINPUT11), .A3(G134), .ZN(new_n258));
  INV_X1    g072(.A(G131), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n256), .A2(new_n258), .A3(new_n259), .A4(new_n251), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n254), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  AND3_X1   g076(.A1(new_n243), .A2(new_n244), .A3(new_n239), .ZN(new_n263));
  AND2_X1   g077(.A1(KEYINPUT0), .A2(G128), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT0), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n265), .A2(new_n200), .A3(KEYINPUT65), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT65), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n267), .B1(KEYINPUT0), .B2(G128), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n264), .B1(new_n235), .B2(new_n239), .ZN(new_n270));
  AOI22_X1  g084(.A1(new_n263), .A2(new_n264), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n256), .A2(new_n251), .A3(new_n258), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G131), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(new_n260), .ZN(new_n274));
  AOI22_X1  g088(.A1(new_n249), .A2(new_n262), .B1(new_n271), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G113), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(KEYINPUT2), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT2), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G113), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT69), .ZN(new_n281));
  INV_X1    g095(.A(G116), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(KEYINPUT69), .A2(G116), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n283), .A2(G119), .A3(new_n284), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n282), .A2(G119), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n280), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT70), .ZN(new_n290));
  AND2_X1   g104(.A1(KEYINPUT69), .A2(G116), .ZN(new_n291));
  NOR2_X1   g105(.A1(KEYINPUT69), .A2(G116), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n286), .B1(new_n293), .B2(G119), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n290), .B1(new_n294), .B2(new_n280), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n285), .A2(new_n280), .A3(new_n290), .A4(new_n287), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n289), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(KEYINPUT71), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n285), .A2(new_n287), .A3(new_n280), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(KEYINPUT70), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n296), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT71), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n302), .A2(new_n303), .A3(new_n289), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n275), .A2(new_n299), .A3(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT28), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT76), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n305), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n303), .B1(new_n302), .B2(new_n289), .ZN(new_n311));
  AOI211_X1 g125(.A(KEYINPUT71), .B(new_n288), .C1(new_n301), .C2(new_n296), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n313), .A2(KEYINPUT76), .A3(new_n275), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n299), .A2(new_n304), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n271), .A2(new_n274), .ZN(new_n316));
  AND2_X1   g130(.A1(new_n244), .A2(new_n239), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT68), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n317), .A2(new_n318), .A3(new_n243), .A4(new_n245), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n246), .A2(KEYINPUT68), .ZN(new_n320));
  AOI22_X1  g134(.A1(new_n319), .A2(new_n320), .B1(new_n240), .B2(new_n237), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n316), .B1(new_n321), .B2(new_n261), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n315), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n310), .A2(new_n314), .A3(new_n323), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n308), .B1(new_n324), .B2(KEYINPUT28), .ZN(new_n325));
  XNOR2_X1  g139(.A(KEYINPUT72), .B(KEYINPUT27), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT73), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n326), .B(new_n327), .ZN(new_n328));
  NOR2_X1   g142(.A1(G237), .A2(G953), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n328), .A2(G210), .A3(new_n329), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n326), .B(KEYINPUT73), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n329), .A2(G210), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT26), .B(G101), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n330), .A2(new_n335), .A3(new_n333), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  AND2_X1   g153(.A1(new_n339), .A2(KEYINPUT29), .ZN(new_n340));
  AOI21_X1  g154(.A(G902), .B1(new_n325), .B2(new_n340), .ZN(new_n341));
  OAI211_X1 g155(.A(KEYINPUT30), .B(new_n316), .C1(new_n321), .C2(new_n261), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n271), .A2(KEYINPUT67), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n270), .A2(new_n269), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n243), .A2(new_n244), .A3(new_n239), .A4(new_n264), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT67), .ZN(new_n347));
  AOI22_X1  g161(.A1(new_n346), .A2(new_n347), .B1(new_n260), .B2(new_n273), .ZN(new_n348));
  AOI22_X1  g162(.A1(new_n343), .A2(new_n348), .B1(new_n249), .B2(new_n262), .ZN(new_n349));
  XOR2_X1   g163(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n342), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n305), .B1(new_n352), .B2(new_n313), .ZN(new_n353));
  INV_X1    g167(.A(new_n339), .ZN(new_n354));
  AOI21_X1  g168(.A(KEYINPUT29), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n313), .A2(KEYINPUT28), .A3(new_n275), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n274), .B1(new_n271), .B2(KEYINPUT67), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n346), .A2(new_n347), .ZN(new_n358));
  OAI22_X1  g172(.A1(new_n357), .A2(new_n358), .B1(new_n321), .B2(new_n261), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n315), .A2(new_n359), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n307), .A2(new_n339), .A3(new_n356), .A4(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(KEYINPUT75), .ZN(new_n362));
  NOR3_X1   g176(.A1(new_n322), .A2(new_n311), .A3(new_n312), .ZN(new_n363));
  AOI22_X1  g177(.A1(new_n363), .A2(KEYINPUT28), .B1(new_n315), .B2(new_n359), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT75), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n364), .A2(new_n365), .A3(new_n339), .A4(new_n307), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n355), .A2(new_n362), .A3(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n233), .B1(new_n341), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(KEYINPUT74), .B1(new_n337), .B2(new_n338), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n369), .B(new_n305), .C1(new_n352), .C2(new_n313), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT31), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n315), .B(new_n342), .C1(new_n349), .C2(new_n351), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n373), .A2(KEYINPUT31), .A3(new_n305), .A4(new_n369), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n364), .A2(new_n307), .ZN(new_n375));
  AOI22_X1  g189(.A1(new_n372), .A2(new_n374), .B1(new_n375), .B2(new_n354), .ZN(new_n376));
  NOR2_X1   g190(.A1(G472), .A2(G902), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(KEYINPUT32), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n375), .A2(new_n354), .ZN(new_n380));
  AOI22_X1  g194(.A1(new_n359), .A2(new_n350), .B1(new_n275), .B2(KEYINPUT30), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n363), .B1(new_n381), .B2(new_n315), .ZN(new_n382));
  AOI21_X1  g196(.A(KEYINPUT31), .B1(new_n382), .B2(new_n369), .ZN(new_n383));
  AND4_X1   g197(.A1(KEYINPUT31), .A2(new_n373), .A3(new_n305), .A4(new_n369), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n380), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT32), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(new_n386), .A3(new_n377), .ZN(new_n387));
  AOI22_X1  g201(.A1(new_n232), .A2(new_n368), .B1(new_n379), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n324), .A2(KEYINPUT28), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(new_n307), .A3(new_n340), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n367), .A2(new_n188), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(G472), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(KEYINPUT77), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n231), .B1(new_n388), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(G214), .B1(G237), .B2(G902), .ZN(new_n395));
  NAND2_X1  g209(.A1(G234), .A2(G237), .ZN(new_n396));
  AND3_X1   g210(.A1(new_n396), .A2(G952), .A3(new_n215), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n396), .A2(G902), .A3(G953), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n398), .B(KEYINPUT94), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(KEYINPUT21), .B(G898), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n397), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G224), .ZN(new_n404));
  OAI21_X1  g218(.A(KEYINPUT7), .B1(new_n404), .B2(G953), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n404), .A2(G953), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n249), .A2(G125), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n271), .A2(new_n207), .ZN(new_n408));
  OAI221_X1 g222(.A(new_n405), .B1(KEYINPUT87), .B2(new_n406), .C1(new_n407), .C2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT86), .ZN(new_n410));
  XNOR2_X1  g224(.A(G110), .B(G122), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n411), .B(KEYINPUT8), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT81), .ZN(new_n413));
  INV_X1    g227(.A(G104), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n413), .B1(new_n414), .B2(G107), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(G107), .ZN(new_n416));
  INV_X1    g230(.A(G107), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n417), .A2(KEYINPUT81), .A3(G104), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n415), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G101), .ZN(new_n420));
  OAI21_X1  g234(.A(KEYINPUT3), .B1(new_n414), .B2(G107), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT3), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n422), .A2(new_n417), .A3(G104), .ZN(new_n423));
  INV_X1    g237(.A(G101), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n421), .A2(new_n423), .A3(new_n424), .A4(new_n416), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n420), .A2(KEYINPUT82), .A3(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT82), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n419), .A2(new_n427), .A3(G101), .ZN(new_n428));
  AND2_X1   g242(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n285), .A2(KEYINPUT5), .A3(new_n287), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT5), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n276), .B1(new_n286), .B2(new_n431), .ZN(new_n432));
  AOI22_X1  g246(.A1(new_n301), .A2(new_n296), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n412), .B1(new_n429), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n430), .A2(new_n432), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n302), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n426), .A2(new_n428), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n410), .B1(new_n434), .B2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n405), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n408), .B1(new_n207), .B2(new_n321), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n406), .A2(KEYINPUT87), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n440), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n436), .A2(new_n437), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n429), .A2(new_n433), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n444), .A2(new_n445), .A3(KEYINPUT86), .A4(new_n412), .ZN(new_n446));
  AND4_X1   g260(.A1(new_n409), .A2(new_n439), .A3(new_n443), .A4(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT84), .ZN(new_n448));
  AND3_X1   g262(.A1(new_n426), .A2(new_n448), .A3(new_n428), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n448), .B1(new_n426), .B2(new_n428), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n433), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n421), .A2(new_n423), .A3(new_n416), .ZN(new_n453));
  NAND2_X1  g267(.A1(KEYINPUT80), .A2(KEYINPUT4), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n453), .A2(G101), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n453), .A2(G101), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n456), .A2(KEYINPUT80), .A3(KEYINPUT4), .A4(new_n425), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n455), .B(new_n457), .C1(new_n311), .C2(new_n312), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n452), .A2(new_n458), .A3(new_n411), .ZN(new_n459));
  AOI21_X1  g273(.A(G902), .B1(new_n447), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(G210), .B1(G237), .B2(G902), .ZN(new_n461));
  INV_X1    g275(.A(new_n411), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n457), .A2(new_n455), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n463), .B1(new_n299), .B2(new_n304), .ZN(new_n464));
  NOR3_X1   g278(.A1(new_n449), .A2(new_n436), .A3(new_n450), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n462), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n466), .A2(new_n459), .A3(KEYINPUT6), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n406), .B(KEYINPUT85), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n441), .B(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT6), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n470), .B(new_n462), .C1(new_n464), .C2(new_n465), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n467), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  AND3_X1   g286(.A1(new_n460), .A2(new_n461), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n461), .B1(new_n460), .B2(new_n472), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n395), .B(new_n403), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(G469), .ZN(new_n477));
  XNOR2_X1  g291(.A(G110), .B(G140), .ZN(new_n478));
  AND2_X1   g292(.A1(new_n215), .A2(G227), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n478), .B(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT83), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n243), .A2(new_n244), .A3(new_n239), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n237), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n484), .B1(new_n247), .B2(new_n248), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n437), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT10), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n482), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AOI211_X1 g302(.A(KEYINPUT83), .B(KEYINPUT10), .C1(new_n485), .C2(new_n437), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n321), .A2(new_n487), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n437), .A2(KEYINPUT84), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n426), .A2(new_n448), .A3(new_n428), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n494), .B1(new_n346), .B2(new_n463), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n274), .B1(new_n490), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n463), .A2(new_n346), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n497), .B1(new_n451), .B2(new_n491), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n319), .A2(new_n320), .ZN(new_n499));
  AOI22_X1  g313(.A1(new_n499), .A2(new_n484), .B1(new_n426), .B2(new_n428), .ZN(new_n500));
  OAI21_X1  g314(.A(KEYINPUT83), .B1(new_n500), .B2(KEYINPUT10), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n486), .A2(new_n482), .A3(new_n487), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n274), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n498), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n481), .B1(new_n496), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n249), .A2(new_n437), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n274), .B1(new_n507), .B2(new_n500), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT12), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n321), .A2(new_n426), .A3(new_n428), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(new_n486), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n512), .A2(KEYINPUT12), .A3(new_n274), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  AND3_X1   g328(.A1(new_n505), .A2(new_n514), .A3(new_n481), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n477), .B(new_n188), .C1(new_n506), .C2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(G469), .A2(G902), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n480), .B(KEYINPUT79), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  AND3_X1   g333(.A1(new_n498), .A2(new_n503), .A3(new_n504), .ZN(new_n520));
  AOI21_X1  g334(.A(KEYINPUT12), .B1(new_n512), .B2(new_n274), .ZN(new_n521));
  AOI211_X1 g335(.A(new_n509), .B(new_n504), .C1(new_n511), .C2(new_n486), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n519), .B1(new_n520), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n496), .A2(new_n505), .A3(new_n481), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(new_n525), .A3(G469), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n516), .A2(new_n517), .A3(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(KEYINPUT9), .B(G234), .ZN(new_n528));
  OAI21_X1  g342(.A(G221), .B1(new_n528), .B2(G902), .ZN(new_n529));
  NOR2_X1   g343(.A1(G475), .A2(G902), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT90), .ZN(new_n531));
  AND2_X1   g345(.A1(KEYINPUT88), .A2(G143), .ZN(new_n532));
  NOR2_X1   g346(.A1(KEYINPUT88), .A2(G143), .ZN(new_n533));
  OAI211_X1 g347(.A(G214), .B(new_n329), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n329), .A2(G214), .ZN(new_n535));
  NAND2_X1  g349(.A1(KEYINPUT88), .A2(G143), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(KEYINPUT18), .A2(G131), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n531), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n534), .A2(new_n537), .A3(KEYINPUT90), .A4(new_n539), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT89), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n534), .A2(new_n537), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n544), .B1(new_n534), .B2(new_n537), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n540), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n190), .B(new_n234), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n543), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n195), .A2(new_n212), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n538), .A2(G131), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT17), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n534), .A2(new_n537), .A3(new_n259), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n538), .A2(KEYINPUT17), .A3(G131), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n550), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  XNOR2_X1  g370(.A(G113), .B(G122), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n557), .B(new_n414), .ZN(new_n558));
  AND3_X1   g372(.A1(new_n549), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n551), .A2(new_n553), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n209), .B(KEYINPUT19), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n560), .B(new_n196), .C1(G146), .C2(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n558), .B1(new_n549), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n530), .B1(new_n559), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(KEYINPUT20), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT20), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n566), .B(new_n530), .C1(new_n559), .C2(new_n563), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n558), .B1(new_n549), .B2(new_n556), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n188), .B1(new_n559), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(G475), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n283), .A2(G122), .A3(new_n284), .ZN(new_n573));
  INV_X1    g387(.A(G122), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(G116), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT14), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(KEYINPUT93), .B1(new_n573), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n573), .A2(KEYINPUT14), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT93), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n573), .A2(new_n577), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(G107), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n238), .A2(G128), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n200), .A2(G143), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n587), .B(G134), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n573), .A2(new_n417), .A3(new_n575), .ZN(new_n589));
  AND2_X1   g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n584), .A2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT92), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT13), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n586), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n587), .A2(new_n594), .A3(G134), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n585), .B(new_n586), .C1(new_n593), .C2(new_n250), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NOR3_X1   g411(.A1(new_n291), .A2(new_n292), .A3(new_n574), .ZN(new_n598));
  INV_X1    g412(.A(new_n575), .ZN(new_n599));
  OAI21_X1  g413(.A(G107), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n589), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT91), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n597), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n600), .A2(new_n589), .A3(KEYINPUT91), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n592), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  AND3_X1   g419(.A1(new_n573), .A2(new_n417), .A3(new_n575), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n417), .B1(new_n573), .B2(new_n575), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n602), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n597), .ZN(new_n609));
  AND4_X1   g423(.A1(new_n592), .A2(new_n608), .A3(new_n604), .A4(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n591), .B1(new_n605), .B2(new_n610), .ZN(new_n611));
  NOR3_X1   g425(.A1(new_n528), .A2(new_n187), .A3(G953), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  OAI211_X1 g428(.A(new_n591), .B(new_n612), .C1(new_n605), .C2(new_n610), .ZN(new_n615));
  AOI21_X1  g429(.A(G902), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(G478), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n617), .A2(KEYINPUT15), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  AOI211_X1 g434(.A(G902), .B(new_n618), .C1(new_n614), .C2(new_n615), .ZN(new_n621));
  NOR3_X1   g435(.A1(new_n572), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  AND3_X1   g436(.A1(new_n527), .A2(new_n529), .A3(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n394), .A2(new_n476), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(G101), .ZN(G3));
  AND3_X1   g439(.A1(new_n527), .A2(new_n230), .A3(new_n529), .ZN(new_n626));
  OAI21_X1  g440(.A(G472), .B1(new_n376), .B2(G902), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n385), .A2(new_n377), .ZN(new_n628));
  AND2_X1   g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n395), .ZN(new_n631));
  INV_X1    g445(.A(new_n461), .ZN(new_n632));
  AND3_X1   g446(.A1(new_n467), .A2(new_n469), .A3(new_n471), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n409), .A2(new_n439), .A3(new_n443), .A4(new_n446), .ZN(new_n634));
  INV_X1    g448(.A(new_n459), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n188), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n632), .B1(new_n633), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n460), .A2(new_n472), .A3(new_n461), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n631), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n617), .A2(new_n188), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n640), .B1(new_n616), .B2(new_n617), .ZN(new_n641));
  INV_X1    g455(.A(new_n615), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n608), .A2(new_n604), .A3(new_n609), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(KEYINPUT92), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n603), .A2(new_n592), .A3(new_n604), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n612), .B1(new_n646), .B2(new_n591), .ZN(new_n647));
  OAI21_X1  g461(.A(KEYINPUT33), .B1(new_n642), .B2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT33), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n614), .A2(new_n649), .A3(new_n615), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n648), .A2(G478), .A3(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n572), .A2(new_n641), .A3(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n639), .A2(KEYINPUT95), .A3(new_n403), .A4(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT95), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n655), .B1(new_n475), .B2(new_n652), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n630), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(KEYINPUT96), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT34), .B(G104), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G6));
  AOI22_X1  g474(.A1(new_n565), .A2(new_n567), .B1(G475), .B2(new_n570), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n661), .B1(new_n620), .B2(new_n621), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n630), .A2(new_n475), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G107), .ZN(new_n664));
  XNOR2_X1  g478(.A(KEYINPUT97), .B(KEYINPUT35), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G9));
  NOR2_X1   g480(.A1(new_n219), .A2(KEYINPUT36), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n214), .B(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n228), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n227), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n627), .A2(new_n628), .A3(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT98), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n627), .A2(new_n628), .A3(KEYINPUT98), .A4(new_n670), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n623), .A2(new_n673), .A3(new_n476), .A4(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT37), .B(G110), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G12));
  INV_X1    g491(.A(KEYINPUT100), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n504), .B1(new_n498), .B2(new_n503), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n480), .B1(new_n520), .B2(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n505), .A2(new_n514), .A3(new_n481), .ZN(new_n681));
  AOI211_X1 g495(.A(G469), .B(G902), .C1(new_n680), .C2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n526), .A2(new_n517), .ZN(new_n683));
  OAI211_X1 g497(.A(new_n529), .B(new_n670), .C1(new_n682), .C2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n395), .B1(new_n473), .B2(new_n474), .ZN(new_n686));
  INV_X1    g500(.A(G900), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n397), .B1(new_n400), .B2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(KEYINPUT99), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  OAI211_X1 g504(.A(new_n661), .B(new_n690), .C1(new_n620), .C2(new_n621), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n686), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n685), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n379), .A2(new_n387), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n391), .A2(new_n232), .A3(G472), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n368), .A2(new_n232), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n678), .B1(new_n693), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n637), .A2(new_n638), .ZN(new_n700));
  INV_X1    g514(.A(new_n691), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n700), .A2(new_n701), .A3(new_n395), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n702), .A2(new_n684), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n393), .A2(new_n694), .A3(new_n695), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n703), .A2(KEYINPUT100), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n699), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G128), .ZN(G30));
  OAI21_X1  g521(.A(new_n529), .B1(new_n682), .B2(new_n683), .ZN(new_n708));
  XOR2_X1   g522(.A(new_n689), .B(KEYINPUT39), .Z(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(KEYINPUT40), .ZN(new_n712));
  XOR2_X1   g526(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n713));
  XNOR2_X1  g527(.A(new_n700), .B(new_n713), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n188), .B1(new_n324), .B2(new_n339), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n382), .A2(new_n354), .ZN(new_n716));
  OAI21_X1  g530(.A(G472), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT102), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n694), .ZN(new_n720));
  INV_X1    g534(.A(new_n670), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n620), .A2(new_n621), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n722), .A2(new_n661), .ZN(new_n723));
  AND4_X1   g537(.A1(new_n395), .A2(new_n720), .A3(new_n721), .A4(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n712), .A2(new_n714), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G143), .ZN(G45));
  NOR2_X1   g540(.A1(new_n652), .A2(new_n689), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n704), .A2(new_n639), .A3(new_n685), .A4(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G146), .ZN(G48));
  NAND2_X1  g543(.A1(new_n656), .A2(new_n654), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n506), .A2(new_n515), .ZN(new_n731));
  OAI21_X1  g545(.A(G469), .B1(new_n731), .B2(G902), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n732), .A2(new_n529), .A3(new_n516), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n730), .A2(new_n394), .A3(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(KEYINPUT41), .B(G113), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n735), .B(new_n736), .ZN(G15));
  NOR2_X1   g551(.A1(new_n475), .A2(new_n662), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n394), .A2(new_n734), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G116), .ZN(G18));
  AOI21_X1  g554(.A(new_n402), .B1(new_n227), .B2(new_n669), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n622), .A2(new_n741), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n733), .A2(new_n686), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n704), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G119), .ZN(G21));
  NOR2_X1   g559(.A1(new_n325), .A2(new_n339), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n383), .A2(new_n384), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n377), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n748), .A2(new_n627), .A3(new_n230), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT103), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n748), .A2(new_n627), .A3(new_n230), .A4(KEYINPUT103), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n639), .A2(new_n723), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n732), .A2(new_n403), .A3(new_n529), .A4(new_n516), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G122), .ZN(G24));
  NOR2_X1   g572(.A1(new_n733), .A2(new_n686), .ZN(new_n759));
  AND3_X1   g573(.A1(new_n748), .A2(new_n627), .A3(new_n670), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n759), .A2(new_n727), .A3(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G125), .ZN(G27));
  NAND3_X1  g576(.A1(new_n637), .A2(new_n395), .A3(new_n638), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n708), .A2(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n704), .A2(new_n764), .A3(new_n230), .A4(new_n727), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT42), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n394), .A2(KEYINPUT42), .A3(new_n727), .A4(new_n764), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G131), .ZN(G33));
  NAND3_X1  g584(.A1(new_n394), .A2(new_n701), .A3(new_n764), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G134), .ZN(G36));
  NAND2_X1  g586(.A1(new_n524), .A2(new_n525), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT45), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n477), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n775), .B1(new_n774), .B2(new_n773), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(KEYINPUT104), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n517), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT46), .ZN(new_n779));
  OAI21_X1  g593(.A(KEYINPUT105), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n682), .B1(new_n778), .B2(new_n779), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT105), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n777), .A2(new_n782), .A3(KEYINPUT46), .A4(new_n517), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n780), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n529), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n785), .A2(new_n710), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n629), .A2(new_n721), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n641), .A2(new_n651), .A3(new_n661), .ZN(new_n788));
  XOR2_X1   g602(.A(new_n788), .B(KEYINPUT43), .Z(new_n789));
  INV_X1    g603(.A(KEYINPUT106), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n789), .A2(new_n790), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n787), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(KEYINPUT44), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n794), .A2(KEYINPUT44), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n796), .A2(new_n763), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n786), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(KEYINPUT107), .B(G137), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n799), .B(new_n800), .ZN(G39));
  INV_X1    g615(.A(KEYINPUT47), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n785), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n784), .A2(KEYINPUT47), .A3(new_n529), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR4_X1   g619(.A1(new_n763), .A2(new_n230), .A3(new_n652), .A4(new_n689), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n805), .A2(new_n698), .A3(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(KEYINPUT108), .B(G140), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n807), .B(new_n808), .ZN(G42));
  NOR2_X1   g623(.A1(new_n714), .A2(new_n720), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n230), .A2(new_n395), .A3(new_n529), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n732), .A2(new_n516), .ZN(new_n812));
  AOI211_X1 g626(.A(new_n788), .B(new_n811), .C1(new_n812), .C2(KEYINPUT49), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n810), .B(new_n813), .C1(KEYINPUT49), .C2(new_n812), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n789), .A2(new_n397), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n733), .A2(new_n763), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(new_n394), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(KEYINPUT48), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n815), .A2(new_n753), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n820), .A2(new_n639), .A3(new_n734), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n215), .A2(G952), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n230), .A2(new_n397), .ZN(new_n823));
  NOR4_X1   g637(.A1(new_n720), .A2(new_n733), .A3(new_n763), .A4(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n822), .B1(new_n824), .B2(new_n653), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n819), .A2(new_n821), .A3(new_n825), .ZN(new_n826));
  OR2_X1    g640(.A1(new_n812), .A2(new_n529), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n803), .A2(new_n804), .A3(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(new_n820), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n829), .A2(new_n763), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n714), .A2(new_n395), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n820), .A2(new_n734), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(KEYINPUT118), .A2(KEYINPUT50), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(KEYINPUT117), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n817), .A2(new_n760), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n572), .B1(new_n651), .B2(new_n641), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n824), .A2(new_n838), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n820), .A2(KEYINPUT117), .A3(new_n734), .A4(new_n832), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n841), .A2(KEYINPUT118), .ZN(new_n842));
  OAI211_X1 g656(.A(new_n836), .B(new_n840), .C1(new_n842), .C2(KEYINPUT50), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n831), .A2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT51), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n826), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n843), .B1(new_n828), .B2(new_n830), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n848), .A2(KEYINPUT119), .A3(KEYINPUT51), .ZN(new_n849));
  AOI21_X1  g663(.A(KEYINPUT119), .B1(new_n848), .B2(KEYINPUT51), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n847), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT53), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT112), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT111), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n722), .A2(new_n661), .A3(new_n690), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n854), .B1(new_n763), .B2(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n473), .A2(new_n474), .ZN(new_n857));
  NOR4_X1   g671(.A1(new_n572), .A2(new_n620), .A3(new_n621), .A4(new_n689), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n857), .A2(new_n858), .A3(KEYINPUT111), .A4(new_n395), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n704), .A2(new_n685), .A3(new_n856), .A4(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n764), .A2(new_n727), .A3(new_n760), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AND4_X1   g676(.A1(new_n704), .A2(new_n764), .A3(new_n230), .A4(new_n701), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n853), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n771), .A2(KEYINPUT112), .A3(new_n860), .A4(new_n861), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT109), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n652), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n572), .A2(new_n641), .A3(new_n651), .A4(KEYINPUT109), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n867), .A2(new_n662), .A3(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n626), .A2(new_n476), .A3(new_n629), .A4(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n704), .A2(new_n230), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n623), .A2(new_n476), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n675), .B(new_n870), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(KEYINPUT110), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT110), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n624), .A2(new_n875), .A3(new_n675), .A4(new_n870), .ZN(new_n876));
  AOI22_X1  g690(.A1(new_n864), .A2(new_n865), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  AOI22_X1  g691(.A1(new_n753), .A2(new_n756), .B1(new_n743), .B2(new_n704), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n878), .A2(new_n735), .A3(new_n739), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n877), .A2(new_n769), .A3(new_n879), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n703), .A2(KEYINPUT100), .A3(new_n704), .ZN(new_n881));
  AOI21_X1  g695(.A(KEYINPUT100), .B1(new_n703), .B2(new_n704), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n761), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(KEYINPUT113), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT113), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n706), .A2(new_n885), .A3(new_n761), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n708), .A2(new_n670), .A3(new_n689), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n887), .A2(new_n639), .A3(new_n720), .A4(new_n723), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n888), .A2(KEYINPUT52), .A3(new_n728), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n884), .A2(new_n886), .A3(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT114), .ZN(new_n891));
  INV_X1    g705(.A(new_n761), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n892), .B1(new_n699), .B2(new_n705), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n888), .A2(new_n728), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT52), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n890), .A2(new_n891), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n891), .B1(new_n890), .B2(new_n897), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n852), .B(new_n880), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n895), .B(KEYINPUT52), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n877), .A2(new_n769), .A3(new_n879), .ZN(new_n902));
  OAI21_X1  g716(.A(KEYINPUT53), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(KEYINPUT54), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n767), .A2(new_n768), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n878), .A2(new_n735), .A3(new_n739), .ZN(new_n907));
  OAI21_X1  g721(.A(KEYINPUT116), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT116), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n879), .A2(new_n909), .A3(new_n769), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n864), .A2(new_n865), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n874), .A2(new_n876), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n912), .A2(new_n913), .A3(KEYINPUT53), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n915), .B1(new_n898), .B2(new_n899), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT54), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n852), .B1(new_n901), .B2(new_n902), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n905), .A2(KEYINPUT115), .A3(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT115), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n904), .A2(new_n921), .A3(KEYINPUT54), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n851), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(G952), .A2(G953), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n814), .B1(new_n923), .B2(new_n924), .ZN(G75));
  NAND4_X1  g739(.A1(new_n877), .A2(new_n908), .A3(new_n910), .A4(KEYINPUT53), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n890), .A2(new_n897), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(KEYINPUT114), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n890), .A2(new_n897), .A3(new_n891), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n926), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n895), .B(new_n896), .ZN(new_n931));
  AOI21_X1  g745(.A(KEYINPUT53), .B1(new_n880), .B2(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n933), .A2(new_n188), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(G210), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT56), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n467), .A2(new_n471), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(new_n469), .ZN(new_n938));
  XNOR2_X1  g752(.A(KEYINPUT120), .B(KEYINPUT55), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n938), .B(new_n939), .ZN(new_n940));
  AND3_X1   g754(.A1(new_n935), .A2(new_n936), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n940), .B1(new_n935), .B2(new_n936), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n215), .A2(G952), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(G51));
  INV_X1    g758(.A(KEYINPUT122), .ZN(new_n945));
  AOI211_X1 g759(.A(new_n188), .B(new_n777), .C1(new_n916), .C2(new_n918), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n517), .B(KEYINPUT121), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT57), .ZN(new_n948));
  AND3_X1   g762(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n917), .B1(new_n916), .B2(new_n918), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n948), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(new_n731), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n946), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n945), .B1(new_n953), .B2(new_n943), .ZN(new_n954));
  INV_X1    g768(.A(new_n943), .ZN(new_n955));
  OAI21_X1  g769(.A(KEYINPUT54), .B1(new_n930), .B2(new_n932), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(new_n919), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n731), .B1(new_n957), .B2(new_n948), .ZN(new_n958));
  OAI211_X1 g772(.A(KEYINPUT122), .B(new_n955), .C1(new_n958), .C2(new_n946), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n954), .A2(new_n959), .ZN(G54));
  NAND3_X1  g774(.A1(new_n934), .A2(KEYINPUT58), .A3(G475), .ZN(new_n961));
  OR2_X1    g775(.A1(new_n559), .A2(new_n563), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n961), .A2(new_n963), .ZN(new_n965));
  NOR3_X1   g779(.A1(new_n964), .A2(new_n965), .A3(new_n943), .ZN(G60));
  NAND2_X1  g780(.A1(new_n648), .A2(new_n650), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n640), .B(KEYINPUT59), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n957), .A2(new_n967), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(new_n955), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n920), .A2(new_n922), .A3(new_n969), .ZN(new_n972));
  INV_X1    g786(.A(new_n967), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n971), .B1(new_n972), .B2(new_n973), .ZN(G63));
  NAND2_X1  g788(.A1(G217), .A2(G902), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT60), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n976), .B1(new_n916), .B2(new_n918), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n943), .B1(new_n977), .B2(new_n668), .ZN(new_n978));
  INV_X1    g792(.A(new_n221), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n979), .B1(new_n933), .B2(new_n976), .ZN(new_n980));
  AOI21_X1  g794(.A(KEYINPUT123), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT61), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n981), .B(new_n982), .ZN(G66));
  OAI21_X1  g797(.A(G953), .B1(new_n401), .B2(new_n404), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n913), .A2(new_n879), .ZN(new_n985));
  INV_X1    g799(.A(new_n985), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n984), .B1(new_n986), .B2(G953), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n937), .B1(G898), .B2(new_n215), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n987), .B(new_n988), .ZN(G69));
  AOI21_X1  g803(.A(new_n215), .B1(G227), .B2(G900), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT126), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g806(.A(new_n992), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n884), .A2(new_n886), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(new_n728), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n871), .A2(new_n754), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n995), .B1(new_n786), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n769), .A2(new_n771), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n998), .B1(new_n786), .B2(new_n798), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n807), .A2(new_n997), .A3(new_n215), .A4(new_n999), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n381), .B(KEYINPUT124), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n1001), .B(new_n561), .Z(new_n1002));
  INV_X1    g816(.A(new_n1002), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n1003), .B1(G900), .B2(G953), .ZN(new_n1004));
  AOI22_X1  g818(.A1(new_n1000), .A2(new_n1004), .B1(new_n991), .B2(new_n990), .ZN(new_n1005));
  INV_X1    g819(.A(new_n995), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1006), .A2(new_n725), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1007), .A2(KEYINPUT62), .ZN(new_n1008));
  INV_X1    g822(.A(KEYINPUT62), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n1006), .A2(new_n1009), .A3(new_n725), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n710), .B1(new_n869), .B2(KEYINPUT125), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n1011), .B1(KEYINPUT125), .B2(new_n869), .ZN(new_n1012));
  NOR4_X1   g826(.A1(new_n1012), .A2(new_n871), .A3(new_n708), .A4(new_n763), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1013), .B1(new_n786), .B2(new_n798), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n1008), .A2(new_n807), .A3(new_n1010), .A4(new_n1014), .ZN(new_n1015));
  AND2_X1   g829(.A1(new_n1015), .A2(new_n215), .ZN(new_n1016));
  OAI211_X1 g830(.A(new_n993), .B(new_n1005), .C1(new_n1016), .C2(new_n1002), .ZN(new_n1017));
  INV_X1    g831(.A(new_n990), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1002), .B1(new_n1015), .B2(new_n215), .ZN(new_n1019));
  AND2_X1   g833(.A1(new_n1000), .A2(new_n1004), .ZN(new_n1020));
  OAI211_X1 g834(.A(KEYINPUT126), .B(new_n1018), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1021));
  AND2_X1   g835(.A1(new_n1017), .A2(new_n1021), .ZN(G72));
  NOR2_X1   g836(.A1(new_n353), .A2(new_n339), .ZN(new_n1023));
  AND4_X1   g837(.A1(new_n807), .A2(new_n997), .A3(new_n986), .A4(new_n999), .ZN(new_n1024));
  NAND2_X1  g838(.A1(G472), .A2(G902), .ZN(new_n1025));
  XOR2_X1   g839(.A(new_n1025), .B(KEYINPUT63), .Z(new_n1026));
  INV_X1    g840(.A(new_n1026), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n1023), .B1(new_n1024), .B2(new_n1027), .ZN(new_n1028));
  NOR3_X1   g842(.A1(new_n716), .A2(new_n1023), .A3(new_n1027), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n943), .B1(new_n904), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g845(.A(KEYINPUT127), .ZN(new_n1032));
  OAI211_X1 g846(.A(new_n1032), .B(new_n1026), .C1(new_n1015), .C2(new_n985), .ZN(new_n1033));
  AND2_X1   g847(.A1(new_n1033), .A2(new_n716), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n1026), .B1(new_n1015), .B2(new_n985), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1035), .A2(KEYINPUT127), .ZN(new_n1036));
  AOI21_X1  g850(.A(new_n1031), .B1(new_n1034), .B2(new_n1036), .ZN(G57));
endmodule


