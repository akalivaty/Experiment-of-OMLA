//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 1 0 0 1 0 1 1 0 1 1 0 1 1 1 1 1 1 0 0 0 1 0 0 1 1 0 0 1 0 1 1 1 0 1 1 0 0 1 0 0 1 1 1 1 0 1 1 0 1 0 1 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n748, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n870, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n880, new_n881, new_n882, new_n883, new_n884, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n959, new_n960, new_n961, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1005, new_n1006;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT31), .B(G50gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G228gat), .ZN(new_n206));
  INV_X1    g005(.A(G233gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  AND2_X1   g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210));
  OAI21_X1  g009(.A(KEYINPUT75), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G155gat), .ZN(new_n212));
  INV_X1    g011(.A(G162gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT75), .ZN(new_n215));
  NAND2_X1  g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT2), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n209), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(G141gat), .B(G148gat), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n211), .B(new_n217), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  XOR2_X1   g020(.A(G141gat), .B(G148gat), .Z(new_n222));
  INV_X1    g021(.A(KEYINPUT76), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n223), .B1(new_n209), .B2(new_n218), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n216), .A2(KEYINPUT76), .A3(KEYINPUT2), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n214), .A2(new_n216), .ZN(new_n226));
  NAND4_X1  g025(.A1(new_n222), .A2(new_n224), .A3(new_n225), .A4(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n221), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G218gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(KEYINPUT73), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT73), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G218gat), .ZN(new_n232));
  AOI21_X1  g031(.A(KEYINPUT22), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(G204gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(G197gat), .ZN(new_n235));
  INV_X1    g034(.A(G197gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(G204gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(G211gat), .B1(new_n233), .B2(new_n238), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n235), .A2(new_n237), .ZN(new_n240));
  INV_X1    g039(.A(G211gat), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n240), .A2(KEYINPUT22), .A3(new_n241), .ZN(new_n242));
  AND3_X1   g041(.A1(new_n239), .A2(new_n229), .A3(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n229), .B1(new_n239), .B2(new_n242), .ZN(new_n244));
  NOR3_X1   g043(.A1(new_n243), .A2(new_n244), .A3(KEYINPUT29), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n228), .B1(new_n245), .B2(KEYINPUT3), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT22), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n231), .A2(G218gat), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n229), .A2(KEYINPUT73), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n241), .B1(new_n250), .B2(new_n240), .ZN(new_n251));
  NOR3_X1   g050(.A1(new_n238), .A2(new_n247), .A3(G211gat), .ZN(new_n252));
  OAI21_X1  g051(.A(G218gat), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n239), .A2(new_n229), .A3(new_n242), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT3), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n221), .A2(new_n227), .A3(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT29), .ZN(new_n257));
  AOI22_X1  g056(.A1(new_n253), .A2(new_n254), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n208), .B1(new_n246), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n228), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n253), .A2(new_n257), .A3(new_n254), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n261), .B1(new_n262), .B2(new_n255), .ZN(new_n263));
  INV_X1    g062(.A(new_n208), .ZN(new_n264));
  NOR3_X1   g063(.A1(new_n263), .A2(new_n264), .A3(new_n258), .ZN(new_n265));
  OAI211_X1 g064(.A(KEYINPUT78), .B(G22gat), .C1(new_n260), .C2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n246), .A2(new_n208), .A3(new_n259), .ZN(new_n267));
  INV_X1    g066(.A(G22gat), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n264), .B1(new_n263), .B2(new_n258), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n266), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n267), .A2(new_n269), .ZN(new_n272));
  AOI21_X1  g071(.A(KEYINPUT78), .B1(new_n272), .B2(G22gat), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n205), .B1(new_n271), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(KEYINPUT79), .A2(G22gat), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n267), .A2(new_n269), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(new_n204), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n275), .B1(new_n267), .B2(new_n269), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n274), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(G227gat), .A2(G233gat), .ZN(new_n282));
  XOR2_X1   g081(.A(new_n282), .B(KEYINPUT64), .Z(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  OR2_X1    g083(.A1(new_n284), .A2(KEYINPUT34), .ZN(new_n285));
  NOR2_X1   g084(.A1(G169gat), .A2(G176gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT23), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT25), .ZN(new_n288));
  AOI22_X1  g087(.A1(new_n288), .A2(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT24), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n290), .A2(G183gat), .A3(G190gat), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT23), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n292), .B1(G169gat), .B2(G176gat), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n287), .A2(new_n289), .A3(new_n291), .A4(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(G183gat), .ZN(new_n295));
  INV_X1    g094(.A(G190gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(G183gat), .A2(G190gat), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n297), .A2(KEYINPUT24), .A3(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  OAI22_X1  g099(.A1(new_n294), .A2(new_n300), .B1(KEYINPUT65), .B2(new_n288), .ZN(new_n301));
  AND2_X1   g100(.A1(new_n287), .A2(new_n293), .ZN(new_n302));
  AND2_X1   g101(.A1(new_n289), .A2(new_n291), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n288), .A2(KEYINPUT65), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n302), .A2(new_n303), .A3(new_n304), .A4(new_n299), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(KEYINPUT27), .B(G183gat), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n307), .A2(KEYINPUT28), .A3(new_n296), .ZN(new_n308));
  OAI21_X1  g107(.A(KEYINPUT27), .B1(new_n295), .B2(KEYINPUT66), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT66), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT27), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n310), .A2(new_n311), .A3(G183gat), .ZN(new_n312));
  AND3_X1   g111(.A1(new_n309), .A2(new_n312), .A3(new_n296), .ZN(new_n313));
  XOR2_X1   g112(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n314));
  OAI21_X1  g113(.A(new_n308), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(G169gat), .A2(G176gat), .ZN(new_n317));
  AND2_X1   g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT26), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n286), .A2(new_n319), .ZN(new_n320));
  AOI22_X1  g119(.A1(new_n318), .A2(new_n320), .B1(G183gat), .B2(G190gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n315), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(G127gat), .ZN(new_n324));
  OAI21_X1  g123(.A(KEYINPUT68), .B1(new_n324), .B2(G134gat), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT1), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n326), .B1(G113gat), .B2(G120gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(G113gat), .A2(G120gat), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n325), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(G127gat), .B(G134gat), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(G113gat), .ZN(new_n334));
  INV_X1    g133(.A(G120gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n336), .A2(new_n326), .A3(new_n328), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n337), .A2(new_n331), .A3(new_n325), .ZN(new_n338));
  AND3_X1   g137(.A1(new_n333), .A2(KEYINPUT69), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(KEYINPUT69), .B1(new_n333), .B2(new_n338), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n323), .A2(new_n341), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n306), .B(new_n322), .C1(new_n339), .C2(new_n340), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n285), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n342), .A2(new_n343), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(new_n282), .ZN(new_n346));
  XNOR2_X1  g145(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n344), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n342), .A2(new_n343), .A3(new_n284), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT33), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(G15gat), .B(G43gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(G71gat), .B(G99gat), .ZN(new_n353));
  XOR2_X1   g152(.A(new_n352), .B(new_n353), .Z(new_n354));
  NAND2_X1  g153(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n348), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n347), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n357), .B1(new_n345), .B2(new_n282), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n351), .B(new_n354), .C1(new_n358), .C2(new_n344), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT71), .ZN(new_n361));
  AND3_X1   g160(.A1(new_n349), .A2(new_n361), .A3(KEYINPUT32), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n361), .B1(new_n349), .B2(KEYINPUT32), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n360), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n356), .A2(new_n364), .A3(new_n359), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n243), .A2(new_n244), .ZN(new_n369));
  NAND2_X1  g168(.A1(G226gat), .A2(G233gat), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n371), .B1(new_n323), .B2(new_n257), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n370), .B1(new_n306), .B2(new_n322), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n369), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n323), .A2(new_n371), .ZN(new_n375));
  INV_X1    g174(.A(new_n369), .ZN(new_n376));
  AOI21_X1  g175(.A(KEYINPUT29), .B1(new_n306), .B2(new_n322), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n375), .B(new_n376), .C1(new_n371), .C2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n374), .A2(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(G8gat), .B(G36gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(G64gat), .B(G92gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n380), .B(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT30), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n379), .A2(KEYINPUT30), .A3(new_n383), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n388), .B1(new_n383), .B2(new_n379), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(G225gat), .A2(G233gat), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n330), .A2(new_n332), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n331), .B1(new_n337), .B2(new_n325), .ZN(new_n394));
  OAI211_X1 g193(.A(new_n227), .B(new_n221), .C1(new_n393), .C2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT4), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n392), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n228), .A2(KEYINPUT3), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n393), .A2(new_n394), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n398), .A2(new_n399), .A3(new_n256), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT69), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n401), .B1(new_n393), .B2(new_n394), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n333), .A2(new_n338), .A3(KEYINPUT69), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n261), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n397), .B(new_n400), .C1(new_n404), .C2(new_n396), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT5), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n399), .A2(new_n228), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(new_n395), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n406), .B1(new_n408), .B2(new_n392), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n404), .A2(new_n396), .ZN(new_n411));
  OR2_X1    g210(.A1(new_n395), .A2(new_n396), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n392), .A2(KEYINPUT5), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n411), .A2(new_n400), .A3(new_n412), .A4(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n410), .A2(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(G1gat), .B(G29gat), .ZN(new_n416));
  INV_X1    g215(.A(G85gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n416), .B(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(KEYINPUT0), .B(G57gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n418), .B(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n415), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT6), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n410), .A2(new_n420), .A3(new_n414), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n420), .B1(new_n410), .B2(new_n414), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(KEYINPUT6), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT35), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  AND4_X1   g227(.A1(new_n281), .A2(new_n368), .A3(new_n390), .A4(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(G22gat), .B1(new_n260), .B2(new_n265), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT78), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n432), .A2(new_n270), .A3(new_n266), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n279), .B1(new_n433), .B2(new_n205), .ZN(new_n434));
  AND3_X1   g233(.A1(new_n356), .A2(new_n359), .A3(new_n364), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n364), .B1(new_n356), .B2(new_n359), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(KEYINPUT81), .B1(new_n434), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT81), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n281), .A2(new_n439), .A3(new_n368), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT74), .ZN(new_n441));
  AOI211_X1 g240(.A(new_n385), .B(new_n382), .C1(new_n374), .C2(new_n378), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n379), .A2(new_n383), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n388), .B(KEYINPUT74), .C1(new_n383), .C2(new_n379), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n444), .A2(new_n445), .A3(new_n386), .ZN(new_n446));
  INV_X1    g245(.A(new_n427), .ZN(new_n447));
  AND3_X1   g246(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT77), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n426), .A2(KEYINPUT6), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n449), .B1(new_n451), .B2(new_n424), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n446), .B1(new_n450), .B2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n438), .A2(new_n440), .A3(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n429), .B1(new_n455), .B2(KEYINPUT35), .ZN(new_n456));
  AND3_X1   g255(.A1(new_n425), .A2(new_n427), .A3(new_n384), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT80), .ZN(new_n458));
  AOI21_X1  g257(.A(KEYINPUT37), .B1(new_n379), .B2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT37), .ZN(new_n460));
  AOI211_X1 g259(.A(KEYINPUT80), .B(new_n460), .C1(new_n374), .C2(new_n378), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n382), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT38), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT38), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n464), .B(new_n382), .C1(new_n459), .C2(new_n461), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n457), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT39), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n412), .A2(new_n400), .ZN(new_n468));
  AOI21_X1  g267(.A(KEYINPUT4), .B1(new_n341), .B2(new_n261), .ZN(new_n469));
  OAI211_X1 g268(.A(new_n467), .B(new_n392), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n468), .A2(new_n469), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n471), .A2(new_n391), .ZN(new_n472));
  OAI21_X1  g271(.A(KEYINPUT39), .B1(new_n408), .B2(new_n392), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n470), .B(new_n420), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT40), .ZN(new_n475));
  OR2_X1    g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n426), .B1(new_n474), .B2(new_n475), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n476), .B(new_n477), .C1(new_n389), .C2(new_n387), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n466), .A2(new_n478), .A3(new_n281), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n427), .B1(new_n425), .B2(KEYINPUT77), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n480), .A2(new_n452), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n434), .B1(new_n481), .B2(new_n446), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT72), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n437), .A2(new_n483), .A3(KEYINPUT36), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT36), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n485), .B1(new_n368), .B2(KEYINPUT72), .ZN(new_n486));
  AND4_X1   g285(.A1(new_n479), .A2(new_n482), .A3(new_n484), .A4(new_n486), .ZN(new_n487));
  OR2_X1    g286(.A1(new_n456), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(G8gat), .ZN(new_n489));
  XNOR2_X1  g288(.A(G15gat), .B(G22gat), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT16), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n490), .B1(new_n491), .B2(G1gat), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n489), .B1(new_n492), .B2(KEYINPUT88), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n492), .B1(G1gat), .B2(new_n490), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI221_X1 g294(.A(new_n492), .B1(KEYINPUT88), .B2(new_n489), .C1(G1gat), .C2(new_n490), .ZN(new_n496));
  AND2_X1   g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT14), .ZN(new_n498));
  INV_X1    g297(.A(G29gat), .ZN(new_n499));
  INV_X1    g298(.A(G36gat), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n502));
  AOI22_X1  g301(.A1(new_n501), .A2(new_n502), .B1(G29gat), .B2(G36gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT85), .ZN(new_n504));
  INV_X1    g303(.A(G43gat), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n505), .A2(G50gat), .ZN(new_n506));
  INV_X1    g305(.A(G50gat), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n507), .A2(G43gat), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT15), .ZN(new_n509));
  NOR3_X1   g308(.A1(new_n506), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n504), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n510), .A2(new_n503), .A3(KEYINPUT85), .ZN(new_n513));
  XOR2_X1   g312(.A(KEYINPUT86), .B(KEYINPUT15), .Z(new_n514));
  OAI21_X1  g313(.A(KEYINPUT87), .B1(new_n507), .B2(G43gat), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n515), .B1(new_n505), .B2(G50gat), .ZN(new_n516));
  NOR3_X1   g315(.A1(new_n507), .A2(KEYINPUT87), .A3(G43gat), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n503), .B(new_n514), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n512), .A2(new_n513), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT17), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT17), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n512), .A2(new_n521), .A3(new_n518), .A4(new_n513), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n497), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT89), .ZN(new_n524));
  NAND2_X1  g323(.A1(G229gat), .A2(G233gat), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT89), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n497), .A2(new_n520), .A3(new_n526), .A4(new_n522), .ZN(new_n527));
  INV_X1    g326(.A(new_n519), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n495), .A2(new_n496), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n524), .A2(new_n525), .A3(new_n527), .A4(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT18), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n497), .A2(new_n519), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(new_n530), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n525), .B(KEYINPUT13), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(KEYINPUT90), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT90), .ZN(new_n539));
  AOI211_X1 g338(.A(new_n539), .B(new_n536), .C1(new_n534), .C2(new_n530), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  AOI22_X1  g340(.A1(new_n523), .A2(KEYINPUT89), .B1(new_n529), .B2(new_n528), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n542), .A2(KEYINPUT18), .A3(new_n525), .A4(new_n527), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n533), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(KEYINPUT82), .B(KEYINPUT11), .ZN(new_n545));
  XOR2_X1   g344(.A(G169gat), .B(G197gat), .Z(new_n546));
  XNOR2_X1  g345(.A(G113gat), .B(G141gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  XOR2_X1   g347(.A(KEYINPUT83), .B(KEYINPUT84), .Z(new_n549));
  OR2_X1    g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n548), .A2(new_n549), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n545), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n550), .A2(new_n545), .A3(new_n551), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT12), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(KEYINPUT12), .B1(new_n553), .B2(new_n554), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n544), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n557), .A2(new_n558), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n560), .A2(new_n533), .A3(new_n541), .A4(new_n543), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  AND2_X1   g361(.A1(new_n488), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT96), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT93), .ZN(new_n565));
  NAND2_X1  g364(.A1(G99gat), .A2(G106gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(KEYINPUT8), .ZN(new_n567));
  NAND2_X1  g366(.A1(G85gat), .A2(G92gat), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT7), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(G92gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n417), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n567), .A2(new_n570), .A3(new_n572), .A4(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G99gat), .B(G106gat), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  AOI22_X1  g376(.A1(KEYINPUT8), .A2(new_n566), .B1(new_n417), .B2(new_n571), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n578), .A2(new_n575), .A3(new_n570), .A4(new_n573), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n565), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  AND2_X1   g379(.A1(new_n579), .A2(new_n565), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n528), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(G232gat), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n584), .A2(new_n207), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(KEYINPUT41), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  AND2_X1   g386(.A1(new_n520), .A2(new_n522), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT94), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n589), .B1(new_n580), .B2(new_n581), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n582), .A2(KEYINPUT94), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n588), .A2(KEYINPUT95), .A3(new_n590), .A4(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT95), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n590), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n520), .A2(new_n522), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n587), .B1(new_n592), .B2(new_n596), .ZN(new_n597));
  XOR2_X1   g396(.A(G190gat), .B(G218gat), .Z(new_n598));
  AOI21_X1  g397(.A(new_n564), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n585), .A2(KEYINPUT41), .ZN(new_n600));
  XNOR2_X1  g399(.A(G134gat), .B(G162gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n597), .A2(new_n598), .ZN(new_n604));
  INV_X1    g403(.A(new_n598), .ZN(new_n605));
  AOI211_X1 g404(.A(new_n605), .B(new_n587), .C1(new_n592), .C2(new_n596), .ZN(new_n606));
  OAI22_X1  g405(.A1(new_n599), .A2(new_n603), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  AND2_X1   g406(.A1(new_n592), .A2(new_n596), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n605), .B1(new_n608), .B2(new_n587), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n597), .A2(new_n598), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n609), .A2(new_n564), .A3(new_n610), .A4(new_n602), .ZN(new_n611));
  AND2_X1   g410(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT97), .ZN(new_n613));
  AND2_X1   g412(.A1(KEYINPUT91), .A2(G57gat), .ZN(new_n614));
  NOR2_X1   g413(.A1(KEYINPUT91), .A2(G57gat), .ZN(new_n615));
  OAI21_X1  g414(.A(G64gat), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(G64gat), .ZN(new_n617));
  AND2_X1   g416(.A1(new_n617), .A2(G57gat), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(G71gat), .A2(G78gat), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(KEYINPUT9), .ZN(new_n622));
  NAND2_X1  g421(.A1(G71gat), .A2(G78gat), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n617), .A2(G57gat), .ZN(new_n625));
  OAI21_X1  g424(.A(KEYINPUT9), .B1(new_n618), .B2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n623), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n627), .A2(new_n621), .ZN(new_n628));
  AOI22_X1  g427(.A1(new_n620), .A2(new_n624), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(KEYINPUT21), .ZN(new_n630));
  OR2_X1    g429(.A1(new_n629), .A2(KEYINPUT21), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n529), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n632), .B1(new_n529), .B2(new_n631), .ZN(new_n633));
  NAND2_X1  g432(.A1(G231gat), .A2(G233gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT92), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(new_n295), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(G211gat), .ZN(new_n637));
  OR2_X1    g436(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n633), .A2(new_n637), .ZN(new_n639));
  XNOR2_X1  g438(.A(G127gat), .B(G155gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  AND3_X1   g441(.A1(new_n638), .A2(new_n639), .A3(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n642), .B1(new_n638), .B2(new_n639), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(G230gat), .A2(G233gat), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n577), .A2(new_n579), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(KEYINPUT93), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n579), .A2(new_n565), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n620), .A2(new_n624), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n626), .A2(new_n628), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n648), .A2(new_n649), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n629), .A2(new_n647), .ZN(new_n654));
  AOI21_X1  g453(.A(KEYINPUT10), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT10), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n582), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n646), .B1(new_n655), .B2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n646), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n653), .A2(new_n661), .A3(new_n654), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(G120gat), .B(G148gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(G176gat), .B(G204gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n666), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n660), .A2(new_n662), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n612), .A2(new_n613), .A3(new_n645), .A4(new_n671), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n645), .A2(new_n607), .A3(new_n611), .A4(new_n671), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(KEYINPUT97), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n563), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(new_n481), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g478(.A1(new_n676), .A2(new_n390), .ZN(new_n680));
  NOR2_X1   g479(.A1(KEYINPUT98), .A2(KEYINPUT42), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(new_n491), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(G8gat), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n680), .A2(new_n489), .A3(new_n682), .ZN(new_n685));
  OR2_X1    g484(.A1(new_n680), .A2(KEYINPUT42), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(KEYINPUT99), .ZN(G1325gat));
  INV_X1    g487(.A(G15gat), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n486), .A2(new_n484), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n676), .A2(new_n689), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n368), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n692), .B1(new_n689), .B2(new_n693), .ZN(G1326gat));
  NOR2_X1   g493(.A1(new_n676), .A2(new_n281), .ZN(new_n695));
  XOR2_X1   g494(.A(KEYINPUT43), .B(G22gat), .Z(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(G1327gat));
  NOR2_X1   g496(.A1(new_n645), .A2(new_n670), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n607), .A2(new_n611), .ZN(new_n699));
  AND2_X1   g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n563), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n481), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n701), .A2(G29gat), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT100), .ZN(new_n704));
  OR2_X1    g503(.A1(new_n704), .A2(KEYINPUT45), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(KEYINPUT45), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n699), .B1(new_n456), .B2(new_n487), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(KEYINPUT44), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n709));
  OAI211_X1 g508(.A(new_n709), .B(new_n699), .C1(new_n456), .C2(new_n487), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n711), .A2(new_n562), .A3(new_n698), .ZN(new_n712));
  OAI21_X1  g511(.A(G29gat), .B1(new_n712), .B2(new_n702), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n705), .A2(new_n706), .A3(new_n713), .ZN(G1328gat));
  NOR3_X1   g513(.A1(new_n701), .A2(G36gat), .A3(new_n390), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT46), .ZN(new_n716));
  OAI21_X1  g515(.A(G36gat), .B1(new_n712), .B2(new_n390), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(G1329gat));
  INV_X1    g517(.A(new_n712), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n719), .A2(G43gat), .A3(new_n690), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT101), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(KEYINPUT47), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n701), .A2(new_n437), .ZN(new_n723));
  OAI211_X1 g522(.A(new_n720), .B(new_n722), .C1(G43gat), .C2(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n721), .A2(KEYINPUT47), .ZN(new_n725));
  XOR2_X1   g524(.A(new_n724), .B(new_n725), .Z(G1330gat));
  NOR3_X1   g525(.A1(new_n701), .A2(G50gat), .A3(new_n281), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n719), .A2(new_n434), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n727), .B1(new_n728), .B2(G50gat), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g529(.A(new_n645), .ZN(new_n731));
  NOR4_X1   g530(.A1(new_n699), .A2(new_n562), .A3(new_n731), .A4(new_n671), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n488), .A2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(new_n481), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n614), .A2(new_n615), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n735), .B(new_n736), .ZN(G1332gat));
  XOR2_X1   g536(.A(new_n733), .B(KEYINPUT102), .Z(new_n738));
  NOR2_X1   g537(.A1(new_n738), .A2(new_n390), .ZN(new_n739));
  NOR2_X1   g538(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n740));
  AND2_X1   g539(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n742), .B1(new_n739), .B2(new_n740), .ZN(G1333gat));
  OAI21_X1  g542(.A(G71gat), .B1(new_n738), .B2(new_n691), .ZN(new_n744));
  OR3_X1    g543(.A1(new_n733), .A2(G71gat), .A3(new_n437), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  XOR2_X1   g545(.A(new_n746), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g546(.A1(new_n738), .A2(new_n281), .ZN(new_n748));
  XOR2_X1   g547(.A(new_n748), .B(G78gat), .Z(G1335gat));
  INV_X1    g548(.A(new_n562), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n488), .A2(new_n750), .A3(new_n699), .A4(new_n731), .ZN(new_n751));
  OR2_X1    g550(.A1(new_n751), .A2(KEYINPUT51), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(KEYINPUT51), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n752), .A2(new_n670), .A3(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  AOI21_X1  g554(.A(G85gat), .B1(new_n755), .B2(new_n481), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n750), .A2(new_n731), .A3(new_n670), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT103), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(KEYINPUT104), .B1(new_n711), .B2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT104), .ZN(new_n761));
  AOI211_X1 g560(.A(new_n761), .B(new_n758), .C1(new_n708), .C2(new_n710), .ZN(new_n762));
  OR2_X1    g561(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n702), .A2(new_n417), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n756), .B1(new_n763), .B2(new_n764), .ZN(G1336gat));
  NOR2_X1   g564(.A1(new_n390), .A2(G92gat), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n752), .A2(new_n670), .A3(new_n753), .A4(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(KEYINPUT52), .B1(new_n767), .B2(KEYINPUT106), .ZN(new_n768));
  INV_X1    g567(.A(new_n390), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n711), .A2(new_n769), .A3(new_n759), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT107), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(G92gat), .B1(new_n770), .B2(new_n771), .ZN(new_n773));
  OAI221_X1 g572(.A(new_n768), .B1(KEYINPUT106), .B2(new_n767), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n769), .B1(new_n760), .B2(new_n762), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT105), .ZN(new_n776));
  AND3_X1   g575(.A1(new_n775), .A2(new_n776), .A3(G92gat), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n776), .B1(new_n775), .B2(G92gat), .ZN(new_n778));
  INV_X1    g577(.A(new_n767), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n777), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT52), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n774), .B1(new_n780), .B2(new_n781), .ZN(G1337gat));
  OR3_X1    g581(.A1(new_n754), .A2(G99gat), .A3(new_n437), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n763), .A2(new_n690), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n784), .A2(KEYINPUT108), .ZN(new_n785));
  OAI21_X1  g584(.A(G99gat), .B1(new_n784), .B2(KEYINPUT108), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n783), .B1(new_n785), .B2(new_n786), .ZN(G1338gat));
  NOR3_X1   g586(.A1(new_n754), .A2(G106gat), .A3(new_n281), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n788), .A2(KEYINPUT53), .ZN(new_n789));
  INV_X1    g588(.A(G106gat), .ZN(new_n790));
  AOI211_X1 g589(.A(new_n281), .B(new_n758), .C1(new_n708), .C2(new_n710), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n790), .B1(new_n763), .B2(new_n434), .ZN(new_n793));
  OAI21_X1  g592(.A(KEYINPUT53), .B1(new_n793), .B2(new_n788), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(G1339gat));
  INV_X1    g594(.A(KEYINPUT110), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n666), .B1(new_n660), .B2(KEYINPUT54), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT54), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n580), .A2(new_n581), .A3(new_n629), .ZN(new_n800));
  INV_X1    g599(.A(new_n654), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n656), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n658), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n799), .B1(new_n803), .B2(new_n646), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n802), .A2(new_n661), .A3(new_n658), .ZN(new_n805));
  AOI21_X1  g604(.A(KEYINPUT109), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n660), .A2(new_n805), .A3(KEYINPUT109), .A4(KEYINPUT54), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  OAI211_X1 g607(.A(KEYINPUT55), .B(new_n798), .C1(new_n806), .C2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n669), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n660), .A2(new_n805), .A3(KEYINPUT54), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT109), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n797), .B1(new_n813), .B2(new_n807), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n814), .A2(KEYINPUT55), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n796), .B1(new_n810), .B2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(new_n669), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n817), .B1(new_n814), .B2(KEYINPUT55), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n798), .B1(new_n806), .B2(new_n808), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n818), .A2(KEYINPUT110), .A3(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n750), .B1(new_n816), .B2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT111), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n535), .A2(new_n537), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n524), .A2(new_n527), .A3(new_n530), .ZN(new_n826));
  INV_X1    g625(.A(new_n525), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n825), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(new_n555), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n824), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n525), .B1(new_n542), .B2(new_n527), .ZN(new_n831));
  OAI211_X1 g630(.A(KEYINPUT111), .B(new_n555), .C1(new_n831), .C2(new_n825), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n561), .A2(new_n830), .A3(new_n670), .A4(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT112), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n833), .B(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n612), .B1(new_n823), .B2(new_n835), .ZN(new_n836));
  AND3_X1   g635(.A1(new_n561), .A2(new_n830), .A3(new_n832), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n810), .A2(new_n815), .A3(new_n796), .ZN(new_n838));
  AOI21_X1  g637(.A(KEYINPUT110), .B1(new_n818), .B2(new_n821), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n699), .B(new_n837), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n645), .B1(new_n836), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n673), .A2(new_n562), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n438), .A2(new_n440), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n481), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT114), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n845), .A2(KEYINPUT114), .A3(new_n481), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n848), .A2(new_n390), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n562), .A2(new_n334), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n851), .B(KEYINPUT115), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n562), .B1(new_n838), .B2(new_n839), .ZN(new_n853));
  XNOR2_X1  g652(.A(new_n833), .B(KEYINPUT112), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n699), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n840), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n731), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(new_n842), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(KEYINPUT113), .B1(new_n859), .B2(new_n281), .ZN(new_n860));
  OAI211_X1 g659(.A(KEYINPUT113), .B(new_n281), .C1(new_n841), .C2(new_n842), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n702), .A2(new_n769), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(new_n368), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n863), .A2(new_n750), .A3(new_n865), .ZN(new_n866));
  OAI22_X1  g665(.A1(new_n850), .A2(new_n852), .B1(new_n866), .B2(new_n334), .ZN(G1340gat));
  INV_X1    g666(.A(new_n850), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n868), .A2(new_n335), .A3(new_n670), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n863), .A2(new_n671), .A3(new_n865), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n869), .B1(new_n870), .B2(new_n335), .ZN(G1341gat));
  NAND2_X1  g670(.A1(new_n645), .A2(new_n324), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n850), .A2(new_n872), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n863), .A2(new_n731), .A3(new_n865), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n874), .A2(new_n324), .ZN(new_n875));
  OAI21_X1  g674(.A(KEYINPUT116), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT116), .ZN(new_n877));
  OAI221_X1 g676(.A(new_n877), .B1(new_n874), .B2(new_n324), .C1(new_n850), .C2(new_n872), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n876), .A2(new_n878), .ZN(G1342gat));
  INV_X1    g678(.A(G134gat), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n699), .A2(new_n880), .ZN(new_n881));
  OR3_X1    g680(.A1(new_n850), .A2(KEYINPUT56), .A3(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(KEYINPUT56), .B1(new_n850), .B2(new_n881), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n863), .A2(new_n612), .A3(new_n865), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n882), .B(new_n883), .C1(new_n880), .C2(new_n884), .ZN(G1343gat));
  NOR2_X1   g684(.A1(new_n843), .A2(new_n281), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n886), .A2(new_n691), .A3(new_n864), .ZN(new_n887));
  INV_X1    g686(.A(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(G141gat), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n888), .A2(new_n889), .A3(new_n562), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n886), .A2(KEYINPUT57), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n562), .A2(new_n818), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT117), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n819), .A2(new_n893), .A3(new_n820), .ZN(new_n894));
  OAI21_X1  g693(.A(KEYINPUT117), .B1(new_n814), .B2(KEYINPUT55), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n833), .B1(new_n892), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n612), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n840), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n842), .B1(new_n899), .B2(new_n731), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT57), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n900), .A2(new_n901), .A3(new_n281), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n891), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n691), .A2(new_n864), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n903), .A2(new_n750), .A3(new_n904), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n890), .B1(new_n905), .B2(new_n889), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(KEYINPUT58), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT58), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n908), .B(new_n890), .C1(new_n905), .C2(new_n889), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n907), .A2(new_n909), .ZN(G1344gat));
  INV_X1    g709(.A(G148gat), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n888), .A2(new_n911), .A3(new_n670), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n903), .A2(new_n904), .ZN(new_n913));
  AOI211_X1 g712(.A(KEYINPUT59), .B(new_n911), .C1(new_n913), .C2(new_n670), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT59), .ZN(new_n915));
  OAI211_X1 g714(.A(KEYINPUT57), .B(new_n434), .C1(new_n841), .C2(new_n842), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(KEYINPUT119), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT119), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n859), .A2(new_n918), .A3(KEYINPUT57), .A4(new_n434), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n672), .A2(new_n750), .A3(new_n674), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT120), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n672), .A2(KEYINPUT120), .A3(new_n750), .A4(new_n674), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT121), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n818), .A2(new_n821), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n925), .B1(new_n612), .B2(new_n926), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n699), .A2(KEYINPUT121), .A3(new_n818), .A4(new_n821), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n927), .A2(new_n837), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n645), .B1(new_n929), .B2(new_n898), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n434), .B1(new_n924), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(new_n901), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n917), .A2(new_n919), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n671), .B1(new_n904), .B2(KEYINPUT118), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n933), .B(new_n934), .C1(KEYINPUT118), .C2(new_n904), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n915), .B1(new_n935), .B2(G148gat), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n912), .B1(new_n914), .B2(new_n936), .ZN(G1345gat));
  AOI21_X1  g736(.A(G155gat), .B1(new_n888), .B2(new_n645), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n731), .A2(new_n212), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n938), .B1(new_n913), .B2(new_n939), .ZN(G1346gat));
  NAND3_X1  g739(.A1(new_n888), .A2(new_n213), .A3(new_n699), .ZN(new_n941));
  NOR3_X1   g740(.A1(new_n903), .A2(new_n612), .A3(new_n904), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n941), .B1(new_n942), .B2(new_n213), .ZN(G1347gat));
  NOR2_X1   g742(.A1(new_n481), .A2(new_n390), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n845), .A2(new_n944), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n945), .A2(G169gat), .A3(new_n750), .ZN(new_n946));
  XOR2_X1   g745(.A(new_n946), .B(KEYINPUT122), .Z(new_n947));
  NAND2_X1  g746(.A1(new_n944), .A2(new_n368), .ZN(new_n948));
  XOR2_X1   g747(.A(new_n948), .B(KEYINPUT123), .Z(new_n949));
  NOR2_X1   g748(.A1(new_n863), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(new_n562), .ZN(new_n951));
  AND3_X1   g750(.A1(new_n951), .A2(KEYINPUT124), .A3(G169gat), .ZN(new_n952));
  AOI21_X1  g751(.A(KEYINPUT124), .B1(new_n951), .B2(G169gat), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n947), .B1(new_n952), .B2(new_n953), .ZN(G1348gat));
  INV_X1    g753(.A(new_n945), .ZN(new_n955));
  AOI21_X1  g754(.A(G176gat), .B1(new_n955), .B2(new_n670), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n670), .A2(G176gat), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n956), .B1(new_n950), .B2(new_n957), .ZN(G1349gat));
  NAND3_X1  g757(.A1(new_n955), .A2(new_n307), .A3(new_n645), .ZN(new_n959));
  NOR3_X1   g758(.A1(new_n863), .A2(new_n731), .A3(new_n949), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n959), .B1(new_n960), .B2(new_n295), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n961), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g761(.A1(new_n955), .A2(new_n296), .A3(new_n699), .ZN(new_n963));
  INV_X1    g762(.A(new_n949), .ZN(new_n964));
  OAI211_X1 g763(.A(new_n699), .B(new_n964), .C1(new_n860), .C2(new_n862), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT61), .ZN(new_n966));
  AND3_X1   g765(.A1(new_n965), .A2(new_n966), .A3(G190gat), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n966), .B1(new_n965), .B2(G190gat), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n963), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(KEYINPUT125), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT125), .ZN(new_n971));
  OAI211_X1 g770(.A(new_n971), .B(new_n963), .C1(new_n967), .C2(new_n968), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n970), .A2(new_n972), .ZN(G1351gat));
  NAND2_X1  g772(.A1(new_n691), .A2(new_n944), .ZN(new_n974));
  AOI22_X1  g773(.A1(new_n916), .A2(KEYINPUT119), .B1(new_n931), .B2(new_n901), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n974), .B1(new_n975), .B2(new_n919), .ZN(new_n976));
  INV_X1    g775(.A(new_n976), .ZN(new_n977));
  OAI21_X1  g776(.A(G197gat), .B1(new_n977), .B2(new_n750), .ZN(new_n978));
  INV_X1    g777(.A(new_n974), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n886), .A2(new_n979), .ZN(new_n980));
  INV_X1    g779(.A(new_n980), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n981), .A2(new_n236), .A3(new_n562), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n978), .A2(new_n982), .ZN(G1352gat));
  NOR2_X1   g782(.A1(new_n671), .A2(G204gat), .ZN(new_n984));
  INV_X1    g783(.A(new_n984), .ZN(new_n985));
  OAI21_X1  g784(.A(KEYINPUT62), .B1(new_n980), .B2(new_n985), .ZN(new_n986));
  INV_X1    g785(.A(KEYINPUT62), .ZN(new_n987));
  NAND4_X1  g786(.A1(new_n886), .A2(new_n987), .A3(new_n979), .A4(new_n984), .ZN(new_n988));
  AND2_X1   g787(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  INV_X1    g788(.A(KEYINPUT126), .ZN(new_n990));
  NAND4_X1  g789(.A1(new_n933), .A2(new_n990), .A3(new_n670), .A4(new_n979), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n991), .A2(G204gat), .ZN(new_n992));
  AOI21_X1  g791(.A(new_n990), .B1(new_n976), .B2(new_n670), .ZN(new_n993));
  OAI21_X1  g792(.A(new_n989), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n994), .A2(KEYINPUT127), .ZN(new_n995));
  INV_X1    g794(.A(KEYINPUT127), .ZN(new_n996));
  OAI211_X1 g795(.A(new_n996), .B(new_n989), .C1(new_n992), .C2(new_n993), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n995), .A2(new_n997), .ZN(G1353gat));
  NAND3_X1  g797(.A1(new_n981), .A2(new_n241), .A3(new_n645), .ZN(new_n999));
  OAI21_X1  g798(.A(G211gat), .B1(new_n977), .B2(new_n731), .ZN(new_n1000));
  INV_X1    g799(.A(KEYINPUT63), .ZN(new_n1001));
  AND2_X1   g800(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1003));
  OAI21_X1  g802(.A(new_n999), .B1(new_n1002), .B2(new_n1003), .ZN(G1354gat));
  AOI21_X1  g803(.A(G218gat), .B1(new_n981), .B2(new_n699), .ZN(new_n1005));
  NOR3_X1   g804(.A1(new_n612), .A2(new_n248), .A3(new_n249), .ZN(new_n1006));
  AOI21_X1  g805(.A(new_n1005), .B1(new_n976), .B2(new_n1006), .ZN(G1355gat));
endmodule


