//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1 0 0 1 1 1 0 1 0 0 1 0 0 0 1 1 0 1 0 1 1 0 0 0 1 1 1 1 1 0 1 0 1 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:47 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n559, new_n560, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n627, new_n628, new_n629, new_n630,
    new_n633, new_n635, new_n636, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT64), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT66), .ZN(G259));
  XOR2_X1   g020(.A(KEYINPUT67), .B(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT68), .Z(new_n455));
  NAND2_X1  g030(.A1(new_n453), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(new_n453), .ZN(new_n458));
  INV_X1    g033(.A(new_n455), .ZN(new_n459));
  AOI22_X1  g034(.A1(new_n458), .A2(G2106), .B1(G567), .B2(new_n459), .ZN(G319));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G137), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n465), .A2(new_n468), .B1(G101), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  INV_X1    g047(.A(G125), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n472), .B1(new_n463), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n468), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n471), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  NOR2_X1   g053(.A1(new_n463), .A2(new_n468), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n463), .A2(G2105), .ZN(new_n480));
  AOI22_X1  g055(.A1(G124), .A2(new_n479), .B1(new_n480), .B2(G136), .ZN(new_n481));
  OAI221_X1 g056(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n468), .C2(G112), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT70), .ZN(G162));
  INV_X1    g059(.A(G114), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT71), .ZN(new_n487));
  XNOR2_X1  g062(.A(new_n486), .B(new_n487), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n463), .ZN(new_n491));
  AND2_X1   g066(.A1(G126), .A2(G2105), .ZN(new_n492));
  AOI22_X1  g067(.A1(new_n488), .A2(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n491), .A2(G138), .A3(new_n468), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n491), .A2(KEYINPUT4), .A3(G138), .A4(new_n468), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n493), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  XNOR2_X1  g074(.A(KEYINPUT6), .B(G651), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G543), .ZN(new_n501));
  INV_X1    g076(.A(G50), .ZN(new_n502));
  NOR2_X1   g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  AND2_X1   g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  AND2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  OAI22_X1  g081(.A1(new_n503), .A2(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G88), .ZN(new_n508));
  OAI22_X1  g083(.A1(new_n501), .A2(new_n502), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  OR2_X1    g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G62), .ZN(new_n514));
  NAND2_X1  g089(.A1(G75), .A2(G543), .ZN(new_n515));
  XNOR2_X1  g090(.A(new_n515), .B(KEYINPUT72), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n510), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n509), .A2(new_n517), .ZN(G166));
  OAI211_X1 g093(.A(G51), .B(G543), .C1(new_n505), .C2(new_n506), .ZN(new_n519));
  AND2_X1   g094(.A1(G63), .A2(G651), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n520), .B1(new_n504), .B2(new_n503), .ZN(new_n521));
  INV_X1    g096(.A(G89), .ZN(new_n522));
  OAI211_X1 g097(.A(new_n519), .B(new_n521), .C1(new_n507), .C2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(KEYINPUT73), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT73), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n527), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n528));
  AND3_X1   g103(.A1(new_n526), .A2(KEYINPUT7), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g104(.A(KEYINPUT7), .B1(new_n526), .B2(new_n528), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n524), .A2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(G168));
  NOR2_X1   g108(.A1(new_n504), .A2(new_n503), .ZN(new_n534));
  INV_X1    g109(.A(G64), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AND2_X1   g111(.A1(G77), .A2(G543), .ZN(new_n537));
  OAI21_X1  g112(.A(G651), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  OR2_X1    g113(.A1(KEYINPUT6), .A2(G651), .ZN(new_n539));
  NAND2_X1  g114(.A1(KEYINPUT6), .A2(G651), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n511), .A2(new_n512), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(G543), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n542), .B1(new_n539), .B2(new_n540), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n541), .A2(G90), .B1(new_n543), .B2(G52), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n538), .A2(new_n544), .ZN(G301));
  INV_X1    g120(.A(G301), .ZN(G171));
  NAND2_X1  g121(.A1(G68), .A2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G56), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n534), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G651), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n513), .A2(new_n500), .A3(G81), .ZN(new_n551));
  OAI211_X1 g126(.A(G43), .B(G543), .C1(new_n505), .C2(new_n506), .ZN(new_n552));
  AND3_X1   g127(.A1(new_n551), .A2(KEYINPUT74), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g128(.A(KEYINPUT74), .B1(new_n551), .B2(new_n552), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n550), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND4_X1  g135(.A1(G319), .A2(G483), .A3(G661), .A4(new_n560), .ZN(G188));
  INV_X1    g136(.A(KEYINPUT77), .ZN(new_n562));
  OAI21_X1  g137(.A(G65), .B1(new_n504), .B2(new_n503), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n563), .A2(KEYINPUT76), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G651), .ZN(new_n566));
  AOI21_X1  g141(.A(KEYINPUT76), .B1(new_n563), .B2(new_n564), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n562), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n563), .A2(new_n564), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT76), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n571), .A2(KEYINPUT77), .A3(G651), .A4(new_n565), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(G53), .ZN(new_n574));
  OR3_X1    g149(.A1(new_n501), .A2(KEYINPUT9), .A3(new_n574), .ZN(new_n575));
  OAI21_X1  g150(.A(KEYINPUT9), .B1(new_n501), .B2(new_n574), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT75), .ZN(new_n577));
  INV_X1    g152(.A(G91), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n507), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n541), .A2(KEYINPUT75), .A3(G91), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n575), .A2(new_n576), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n573), .A2(new_n581), .ZN(G299));
  AOI22_X1  g157(.A1(new_n541), .A2(G89), .B1(new_n513), .B2(new_n520), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT78), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n583), .A2(new_n531), .A3(new_n584), .A4(new_n519), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n526), .A2(new_n528), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT7), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n526), .A2(KEYINPUT7), .A3(new_n528), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g165(.A(KEYINPUT78), .B1(new_n590), .B2(new_n523), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n585), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(G286));
  INV_X1    g168(.A(G166), .ZN(G303));
  OAI21_X1  g169(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n543), .A2(G49), .ZN(new_n596));
  INV_X1    g171(.A(G87), .ZN(new_n597));
  OAI211_X1 g172(.A(new_n595), .B(new_n596), .C1(new_n597), .C2(new_n507), .ZN(G288));
  AOI22_X1  g173(.A1(new_n513), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n599), .A2(new_n510), .ZN(new_n600));
  INV_X1    g175(.A(G48), .ZN(new_n601));
  INV_X1    g176(.A(G86), .ZN(new_n602));
  OAI22_X1  g177(.A1(new_n501), .A2(new_n601), .B1(new_n507), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(G305));
  AOI22_X1  g180(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n606));
  OR2_X1    g181(.A1(new_n606), .A2(new_n510), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n541), .A2(G85), .B1(new_n543), .B2(G47), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(G290));
  NAND2_X1  g184(.A1(G301), .A2(G868), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT10), .ZN(new_n611));
  INV_X1    g186(.A(G92), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n507), .B2(new_n612), .ZN(new_n613));
  NAND4_X1  g188(.A1(new_n513), .A2(new_n500), .A3(KEYINPUT10), .A4(G92), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(G66), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(KEYINPUT79), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT79), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(G66), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n617), .B(new_n619), .C1(new_n504), .C2(new_n503), .ZN(new_n620));
  NAND2_X1  g195(.A1(G79), .A2(G543), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AOI22_X1  g197(.A1(new_n622), .A2(G651), .B1(G54), .B2(new_n543), .ZN(new_n623));
  AND2_X1   g198(.A1(new_n615), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n610), .B1(new_n624), .B2(G868), .ZN(G284));
  OAI21_X1  g200(.A(new_n610), .B1(new_n624), .B2(G868), .ZN(G321));
  AND3_X1   g201(.A1(G286), .A2(KEYINPUT80), .A3(G868), .ZN(new_n627));
  INV_X1    g202(.A(G868), .ZN(new_n628));
  NAND2_X1  g203(.A1(G299), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g204(.A(KEYINPUT80), .B1(G286), .B2(G868), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n627), .B1(new_n629), .B2(new_n630), .ZN(G297));
  AOI21_X1  g206(.A(new_n627), .B1(new_n629), .B2(new_n630), .ZN(G280));
  INV_X1    g207(.A(G559), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n624), .B1(new_n633), .B2(G860), .ZN(G148));
  NAND2_X1  g209(.A1(new_n624), .A2(new_n633), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(KEYINPUT81), .Z(new_n636));
  MUX2_X1   g211(.A(new_n555), .B(new_n636), .S(G868), .Z(G323));
  XNOR2_X1  g212(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g213(.A1(new_n491), .A2(new_n470), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT12), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT13), .ZN(new_n641));
  INV_X1    g216(.A(G2100), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT82), .Z(new_n644));
  AOI22_X1  g219(.A1(G123), .A2(new_n479), .B1(new_n480), .B2(G135), .ZN(new_n645));
  OAI21_X1  g220(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n646), .A2(KEYINPUT83), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(KEYINPUT83), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n648), .B1(new_n468), .B2(G111), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n645), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(G2096), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  OAI211_X1 g227(.A(new_n644), .B(new_n652), .C1(new_n642), .C2(new_n641), .ZN(G156));
  XOR2_X1   g228(.A(KEYINPUT15), .B(G2435), .Z(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT84), .B(G2438), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2427), .B(G2430), .Z(new_n657));
  OAI21_X1  g232(.A(KEYINPUT14), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT85), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n656), .A2(new_n657), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2443), .B(G2446), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1341), .B(G1348), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2451), .B(G2454), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT16), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n668), .A2(G14), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n665), .A2(new_n667), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT86), .ZN(G401));
  INV_X1    g247(.A(KEYINPUT18), .ZN(new_n673));
  XOR2_X1   g248(.A(G2084), .B(G2090), .Z(new_n674));
  XNOR2_X1  g249(.A(G2067), .B(G2678), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n676), .A2(KEYINPUT17), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n674), .A2(new_n675), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n673), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(new_n642), .ZN(new_n680));
  XOR2_X1   g255(.A(G2072), .B(G2078), .Z(new_n681));
  AOI21_X1  g256(.A(new_n681), .B1(new_n676), .B2(KEYINPUT18), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(new_n651), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n680), .B(new_n683), .ZN(G227));
  XOR2_X1   g259(.A(G1971), .B(G1976), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT19), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1956), .B(G2474), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1961), .B(G1966), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT20), .ZN(new_n691));
  AND2_X1   g266(.A1(new_n687), .A2(new_n688), .ZN(new_n692));
  NOR3_X1   g267(.A1(new_n686), .A2(new_n689), .A3(new_n692), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n693), .B1(new_n686), .B2(new_n692), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT87), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n695), .B(new_n697), .Z(new_n698));
  XNOR2_X1  g273(.A(G1991), .B(G1996), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1981), .B(G1986), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(G229));
  AND2_X1   g278(.A1(G288), .A2(KEYINPUT89), .ZN(new_n704));
  NOR2_X1   g279(.A1(G288), .A2(KEYINPUT89), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(new_n707), .B2(G23), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT33), .B(G1976), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n707), .A2(G22), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G166), .B2(new_n707), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT90), .Z(new_n713));
  AOI22_X1  g288(.A1(new_n709), .A2(new_n710), .B1(new_n713), .B2(G1971), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G1971), .B2(new_n713), .ZN(new_n715));
  NOR2_X1   g290(.A1(G6), .A2(G16), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(new_n604), .B2(G16), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT32), .B(G1981), .Z(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(new_n709), .B2(new_n710), .ZN(new_n720));
  OR3_X1    g295(.A1(new_n715), .A2(KEYINPUT34), .A3(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(KEYINPUT34), .B1(new_n715), .B2(new_n720), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n707), .A2(G24), .ZN(new_n723));
  INV_X1    g298(.A(G290), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n723), .B1(new_n724), .B2(new_n707), .ZN(new_n725));
  INV_X1    g300(.A(G1986), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G29), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G25), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n479), .A2(G119), .ZN(new_n730));
  OAI221_X1 g305(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n468), .C2(G107), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n480), .A2(G131), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n730), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT88), .Z(new_n734));
  OAI21_X1  g309(.A(new_n729), .B1(new_n734), .B2(new_n728), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT35), .B(G1991), .Z(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n727), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(new_n735), .B2(new_n737), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n721), .A2(new_n722), .A3(new_n739), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT36), .Z(new_n741));
  NAND2_X1  g316(.A1(new_n728), .A2(G35), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G162), .B2(new_n728), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT29), .ZN(new_n744));
  INV_X1    g319(.A(G2090), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n728), .A2(G26), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT28), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n480), .A2(G140), .ZN(new_n749));
  NOR2_X1   g324(.A1(G104), .A2(G2105), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT93), .ZN(new_n751));
  OAI21_X1  g326(.A(G2104), .B1(new_n468), .B2(G116), .ZN(new_n752));
  AND3_X1   g327(.A1(new_n479), .A2(KEYINPUT92), .A3(G128), .ZN(new_n753));
  AOI21_X1  g328(.A(KEYINPUT92), .B1(new_n479), .B2(G128), .ZN(new_n754));
  OAI221_X1 g329(.A(new_n749), .B1(new_n751), .B2(new_n752), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(G29), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n756), .A2(KEYINPUT94), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n756), .A2(KEYINPUT94), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n748), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(G2067), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n556), .A2(new_n707), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n707), .B2(G19), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  AND2_X1   g339(.A1(new_n764), .A2(G1341), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n764), .A2(G1341), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n707), .A2(G4), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(new_n624), .B2(new_n707), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT91), .B(G1348), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n768), .B(new_n769), .Z(new_n770));
  INV_X1    g345(.A(G34), .ZN(new_n771));
  AOI21_X1  g346(.A(G29), .B1(new_n771), .B2(KEYINPUT24), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(KEYINPUT24), .B2(new_n771), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(new_n477), .B2(new_n728), .ZN(new_n774));
  INV_X1    g349(.A(G2084), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT96), .ZN(new_n777));
  NOR4_X1   g352(.A1(new_n765), .A2(new_n766), .A3(new_n770), .A4(new_n777), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n746), .A2(new_n761), .A3(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(G171), .A2(new_n707), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G5), .B2(new_n707), .ZN(new_n781));
  INV_X1    g356(.A(G1961), .ZN(new_n782));
  AND2_X1   g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT97), .B(KEYINPUT26), .ZN(new_n784));
  NAND3_X1  g359(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G105), .B2(new_n470), .ZN(new_n787));
  AOI22_X1  g362(.A1(G129), .A2(new_n479), .B1(new_n480), .B2(G141), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n790), .A2(new_n728), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(new_n728), .B2(G32), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT27), .B(G1996), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AOI211_X1 g369(.A(new_n783), .B(new_n794), .C1(new_n775), .C2(new_n774), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n795), .A2(KEYINPUT100), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n728), .A2(G27), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G164), .B2(new_n728), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT101), .Z(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n800), .A2(G2078), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT25), .Z(new_n803));
  NAND2_X1  g378(.A1(new_n480), .A2(G139), .ZN(new_n804));
  AOI22_X1  g379(.A1(new_n491), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n805));
  OAI211_X1 g380(.A(new_n803), .B(new_n804), .C1(new_n468), .C2(new_n805), .ZN(new_n806));
  MUX2_X1   g381(.A(G33), .B(new_n806), .S(G29), .Z(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT95), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n808), .A2(G2072), .ZN(new_n809));
  NOR3_X1   g384(.A1(new_n796), .A2(new_n801), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n707), .A2(G20), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT23), .Z(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(G299), .B2(G16), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(G1956), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT31), .B(G11), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT30), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n728), .B1(new_n816), .B2(G28), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n817), .A2(KEYINPUT99), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n816), .A2(G28), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(new_n817), .B2(KEYINPUT99), .ZN(new_n820));
  OAI221_X1 g395(.A(new_n815), .B1(new_n818), .B2(new_n820), .C1(new_n650), .C2(new_n728), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(new_n792), .B2(new_n793), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n707), .A2(G21), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(G168), .B2(new_n707), .ZN(new_n824));
  XNOR2_X1  g399(.A(KEYINPUT98), .B(G1966), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n822), .B(new_n826), .C1(new_n782), .C2(new_n781), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(G2078), .B2(new_n800), .ZN(new_n828));
  AOI22_X1  g403(.A1(new_n795), .A2(KEYINPUT100), .B1(G2072), .B2(new_n808), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n810), .A2(new_n814), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  NOR3_X1   g405(.A1(new_n741), .A2(new_n779), .A3(new_n830), .ZN(G311));
  INV_X1    g406(.A(G311), .ZN(G150));
  NAND2_X1  g407(.A1(new_n624), .A2(G559), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT103), .ZN(new_n834));
  INV_X1    g409(.A(G55), .ZN(new_n835));
  INV_X1    g410(.A(G93), .ZN(new_n836));
  OAI22_X1  g411(.A1(new_n501), .A2(new_n835), .B1(new_n507), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(G67), .B1(new_n504), .B2(new_n503), .ZN(new_n838));
  NAND2_X1  g413(.A1(G80), .A2(G543), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n510), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n555), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n837), .A2(new_n840), .ZN(new_n843));
  OAI211_X1 g418(.A(new_n843), .B(new_n550), .C1(new_n554), .C2(new_n553), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n834), .B(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT39), .ZN(new_n850));
  AOI21_X1  g425(.A(G860), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n851), .B1(new_n850), .B2(new_n849), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n841), .A2(G860), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(KEYINPUT37), .Z(new_n854));
  NAND2_X1  g429(.A1(new_n852), .A2(new_n854), .ZN(G145));
  XOR2_X1   g430(.A(new_n733), .B(KEYINPUT105), .Z(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n640), .ZN(new_n857));
  AOI22_X1  g432(.A1(G130), .A2(new_n479), .B1(new_n480), .B2(G142), .ZN(new_n858));
  OAI221_X1 g433(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n468), .C2(G118), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n857), .B(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(KEYINPUT106), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n861), .A2(KEYINPUT106), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n755), .B(new_n789), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(new_n806), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n498), .B(KEYINPUT104), .Z(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n866), .A2(new_n867), .ZN(new_n870));
  OAI22_X1  g445(.A1(new_n863), .A2(new_n864), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OR2_X1    g446(.A1(new_n861), .A2(KEYINPUT106), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n869), .A2(new_n870), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n872), .A2(new_n873), .A3(new_n862), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(G162), .B(G160), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(new_n650), .ZN(new_n877));
  AOI21_X1  g452(.A(G37), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n863), .A2(new_n864), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n877), .B1(new_n879), .B2(new_n873), .ZN(new_n880));
  NOR3_X1   g455(.A1(new_n869), .A2(KEYINPUT107), .A3(new_n870), .ZN(new_n881));
  OAI21_X1  g456(.A(KEYINPUT107), .B1(new_n869), .B2(new_n870), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n857), .B(new_n860), .Z(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n880), .B1(new_n881), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n878), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g462(.A(KEYINPUT108), .B1(new_n843), .B2(G868), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n636), .B(new_n845), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n624), .B1(new_n573), .B2(new_n581), .ZN(new_n890));
  AND3_X1   g465(.A1(new_n573), .A2(new_n581), .A3(new_n624), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n636), .B(new_n846), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT41), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n894), .B1(new_n891), .B2(new_n890), .ZN(new_n895));
  INV_X1    g470(.A(new_n624), .ZN(new_n896));
  NAND2_X1  g471(.A1(G299), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n573), .A2(new_n624), .A3(new_n581), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n897), .A2(KEYINPUT41), .A3(new_n898), .ZN(new_n899));
  AND2_X1   g474(.A1(new_n895), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n893), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n892), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(KEYINPUT42), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT42), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n892), .A2(new_n905), .A3(new_n902), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n706), .A2(G305), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n604), .B1(new_n704), .B2(new_n705), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n724), .A2(G303), .ZN(new_n911));
  NAND2_X1  g486(.A1(G290), .A2(G166), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n908), .A2(new_n912), .A3(new_n911), .A4(new_n909), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n907), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n904), .A2(new_n916), .A3(new_n906), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n918), .A2(G868), .A3(new_n919), .ZN(new_n920));
  MUX2_X1   g495(.A(KEYINPUT108), .B(new_n888), .S(new_n920), .Z(G295));
  MUX2_X1   g496(.A(KEYINPUT108), .B(new_n888), .S(new_n920), .Z(G331));
  AOI21_X1  g497(.A(new_n584), .B1(new_n524), .B2(new_n531), .ZN(new_n923));
  NOR3_X1   g498(.A1(new_n590), .A2(new_n523), .A3(KEYINPUT78), .ZN(new_n924));
  OAI21_X1  g499(.A(G171), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  AOI22_X1  g500(.A1(new_n524), .A2(new_n531), .B1(new_n538), .B2(new_n544), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n925), .A2(new_n842), .A3(new_n844), .A4(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT109), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(G301), .B1(new_n585), .B2(new_n591), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n845), .B1(new_n931), .B2(new_n926), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n926), .B1(new_n592), .B2(G171), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n933), .A2(KEYINPUT109), .A3(new_n842), .A4(new_n844), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n930), .A2(new_n932), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(new_n900), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n891), .A2(new_n890), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n937), .A2(new_n932), .A3(new_n928), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n916), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n930), .A2(new_n937), .A3(new_n932), .A4(new_n934), .ZN(new_n940));
  NOR3_X1   g515(.A1(new_n845), .A2(new_n931), .A3(new_n926), .ZN(new_n941));
  AOI22_X1  g516(.A1(new_n925), .A2(new_n927), .B1(new_n842), .B2(new_n844), .ZN(new_n942));
  OAI211_X1 g517(.A(new_n895), .B(new_n899), .C1(new_n941), .C2(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n940), .A2(new_n943), .A3(new_n916), .ZN(new_n944));
  INV_X1    g519(.A(G37), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(KEYINPUT43), .B1(new_n939), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n940), .A2(new_n943), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n917), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n949), .A2(KEYINPUT110), .A3(new_n945), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT110), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n916), .B1(new_n940), .B2(new_n943), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n951), .B1(new_n952), .B2(G37), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n950), .A2(new_n953), .A3(new_n944), .ZN(new_n954));
  OAI211_X1 g529(.A(KEYINPUT44), .B(new_n947), .C1(new_n954), .C2(KEYINPUT43), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT111), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n957));
  NOR3_X1   g532(.A1(new_n939), .A2(new_n946), .A3(KEYINPUT43), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT44), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n956), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n958), .B1(new_n954), .B2(KEYINPUT43), .ZN(new_n963));
  NOR3_X1   g538(.A1(new_n963), .A2(KEYINPUT111), .A3(KEYINPUT44), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n955), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT112), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT112), .ZN(new_n967));
  OAI211_X1 g542(.A(new_n967), .B(new_n955), .C1(new_n962), .C2(new_n964), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n966), .A2(new_n968), .ZN(G397));
  XOR2_X1   g544(.A(KEYINPUT113), .B(G1384), .Z(new_n970));
  NAND2_X1  g545(.A1(new_n498), .A2(new_n970), .ZN(new_n971));
  XOR2_X1   g546(.A(KEYINPUT114), .B(KEYINPUT45), .Z(new_n972));
  AND2_X1   g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT115), .ZN(new_n975));
  NAND3_X1  g550(.A1(G160), .A2(new_n975), .A3(G40), .ZN(new_n976));
  INV_X1    g551(.A(G40), .ZN(new_n977));
  OAI21_X1  g552(.A(KEYINPUT115), .B1(new_n477), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n974), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(G1996), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n982), .B(KEYINPUT117), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n983), .A2(new_n789), .ZN(new_n984));
  INV_X1    g559(.A(new_n980), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n755), .B(new_n760), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n789), .A2(G1996), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n985), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n984), .A2(new_n988), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n733), .B(new_n736), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n989), .B1(new_n985), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n724), .A2(new_n726), .ZN(new_n992));
  XOR2_X1   g567(.A(new_n992), .B(KEYINPUT116), .Z(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n994), .B1(new_n726), .B2(new_n724), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n991), .B1(new_n980), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G1384), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n498), .A2(new_n997), .ZN(new_n998));
  OR2_X1    g573(.A1(new_n979), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT119), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n1000), .B1(G305), .B2(G1981), .ZN(new_n1001));
  INV_X1    g576(.A(G1981), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n604), .A2(KEYINPUT119), .A3(new_n1002), .ZN(new_n1003));
  AOI22_X1  g578(.A1(new_n1001), .A2(new_n1003), .B1(G1981), .B2(G305), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n999), .B(G8), .C1(KEYINPUT49), .C2(new_n1004), .ZN(new_n1005));
  AND2_X1   g580(.A1(new_n1004), .A2(KEYINPUT49), .ZN(new_n1006));
  OR2_X1    g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g582(.A1(G288), .A2(G1976), .ZN(new_n1008));
  AOI22_X1  g583(.A1(new_n1007), .A2(new_n1008), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n999), .A2(G8), .ZN(new_n1010));
  INV_X1    g585(.A(G8), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n998), .A2(KEYINPUT50), .ZN(new_n1012));
  AND3_X1   g587(.A1(new_n1012), .A2(new_n978), .A3(new_n976), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT50), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n498), .A2(new_n1014), .A3(new_n997), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1013), .A2(new_n745), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n998), .A2(new_n972), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n498), .A2(KEYINPUT45), .A3(new_n970), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1017), .A2(new_n978), .A3(new_n976), .A4(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g594(.A(KEYINPUT118), .B(G1971), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1011), .B1(new_n1016), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(G303), .A2(G8), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n1023), .B(KEYINPUT55), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1022), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n706), .A2(G1976), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n999), .A2(G8), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(KEYINPUT52), .ZN(new_n1029));
  INV_X1    g604(.A(G1976), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT52), .B1(G288), .B2(new_n1030), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n999), .A2(G8), .A3(new_n1027), .A4(new_n1031), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n1029), .B(new_n1032), .C1(new_n1006), .C2(new_n1005), .ZN(new_n1033));
  OAI22_X1  g608(.A1(new_n1009), .A2(new_n1010), .B1(new_n1026), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1033), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1012), .A2(new_n978), .A3(new_n976), .A4(new_n1015), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1036), .A2(G2084), .ZN(new_n1037));
  AND2_X1   g612(.A1(new_n976), .A2(new_n978), .ZN(new_n1038));
  OR2_X1    g613(.A1(new_n998), .A2(new_n972), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT45), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n998), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1038), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(G1966), .ZN(new_n1043));
  AOI22_X1  g618(.A1(new_n1037), .A2(KEYINPUT121), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT121), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1045), .B1(new_n1036), .B2(G2084), .ZN(new_n1046));
  AOI211_X1 g621(.A(new_n1011), .B(G286), .C1(new_n1044), .C2(new_n1046), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1035), .B(new_n1047), .C1(new_n1025), .C2(new_n1022), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1034), .B1(KEYINPUT63), .B2(new_n1048), .ZN(new_n1049));
  XOR2_X1   g624(.A(KEYINPUT122), .B(G1956), .Z(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1038), .A2(new_n1012), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT120), .ZN(new_n1053));
  XNOR2_X1  g628(.A(new_n1015), .B(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1051), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  XOR2_X1   g630(.A(G299), .B(KEYINPUT57), .Z(new_n1056));
  AND3_X1   g631(.A1(new_n976), .A2(new_n978), .A3(new_n1018), .ZN(new_n1057));
  XNOR2_X1  g632(.A(KEYINPUT56), .B(G2072), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1057), .A2(new_n1017), .A3(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1055), .A2(new_n1056), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1038), .A2(new_n997), .A3(new_n760), .A4(new_n498), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1036), .A2(new_n769), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1062), .A2(new_n1063), .A3(KEYINPUT123), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT123), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1065));
  OR3_X1    g640(.A1(new_n1064), .A2(new_n1065), .A3(new_n896), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1056), .ZN(new_n1067));
  XNOR2_X1  g642(.A(new_n1015), .B(KEYINPUT120), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1050), .B1(new_n1068), .B2(new_n1013), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1059), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1067), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1061), .B1(new_n1066), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1060), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT61), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1071), .A2(new_n1060), .A3(KEYINPUT61), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(KEYINPUT60), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1078));
  AND2_X1   g653(.A1(new_n896), .A2(KEYINPUT126), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n896), .A2(KEYINPUT126), .ZN(new_n1080));
  OR3_X1    g655(.A1(new_n1078), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  NOR3_X1   g656(.A1(new_n1064), .A2(new_n1065), .A3(KEYINPUT60), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1082), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1077), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT124), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1085), .B1(new_n1019), .B2(G1996), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1057), .A2(KEYINPUT124), .A3(new_n981), .A4(new_n1017), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  XOR2_X1   g663(.A(KEYINPUT58), .B(G1341), .Z(new_n1089));
  NAND2_X1  g664(.A1(new_n999), .A2(new_n1089), .ZN(new_n1090));
  AND3_X1   g665(.A1(new_n1088), .A2(KEYINPUT125), .A3(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(KEYINPUT125), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n556), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT59), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT59), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n1095), .B(new_n556), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1072), .B1(new_n1084), .B2(new_n1097), .ZN(new_n1098));
  OR2_X1    g673(.A1(new_n1019), .A2(G2078), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT53), .ZN(new_n1100));
  AOI22_X1  g675(.A1(new_n1099), .A2(new_n1100), .B1(new_n782), .B2(new_n1036), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1100), .A2(G2078), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  OR2_X1    g678(.A1(new_n1042), .A2(new_n1103), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n1101), .A2(G301), .A3(new_n1104), .ZN(new_n1105));
  NOR3_X1   g680(.A1(new_n477), .A2(new_n977), .A3(new_n1103), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n974), .A2(new_n1018), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(G301), .B1(new_n1101), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT54), .ZN(new_n1109));
  NOR3_X1   g684(.A1(new_n1105), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1068), .A2(new_n1013), .A3(new_n745), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n1111), .A2(new_n1021), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1024), .B1(new_n1112), .B2(new_n1011), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1035), .A2(new_n1113), .A3(new_n1026), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1110), .A2(new_n1114), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1013), .A2(KEYINPUT121), .A3(new_n775), .A4(new_n1015), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1116), .A2(new_n1117), .A3(G168), .A4(new_n1046), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(G8), .ZN(new_n1119));
  OR2_X1    g694(.A1(new_n1119), .A2(KEYINPUT51), .ZN(new_n1120));
  AOI21_X1  g695(.A(G168), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1121));
  OAI21_X1  g696(.A(KEYINPUT51), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  AND3_X1   g698(.A1(new_n1101), .A2(G301), .A3(new_n1107), .ZN(new_n1124));
  AOI21_X1  g699(.A(G301), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1109), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1115), .A2(new_n1123), .A3(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1049), .B1(new_n1098), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1123), .A2(KEYINPUT62), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT62), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1120), .A2(new_n1122), .A3(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1129), .A2(new_n1125), .A3(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT63), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1047), .A2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1114), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n996), .B1(new_n1128), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n734), .A2(new_n736), .ZN(new_n1137));
  NOR3_X1   g712(.A1(new_n984), .A2(new_n988), .A3(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n755), .A2(G2067), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n980), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n993), .A2(new_n980), .ZN(new_n1141));
  XOR2_X1   g716(.A(new_n1141), .B(KEYINPUT48), .Z(new_n1142));
  AOI21_X1  g717(.A(new_n985), .B1(new_n986), .B2(new_n790), .ZN(new_n1143));
  OR2_X1    g718(.A1(new_n983), .A2(KEYINPUT46), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n983), .A2(KEYINPUT46), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1143), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT47), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  AOI211_X1 g723(.A(KEYINPUT47), .B(new_n1143), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1149));
  OAI221_X1 g724(.A(new_n1140), .B1(new_n991), .B2(new_n1142), .C1(new_n1148), .C2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1136), .A2(new_n1151), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g727(.A(new_n671), .ZN(new_n1154));
  INV_X1    g728(.A(G227), .ZN(new_n1155));
  NAND2_X1  g729(.A1(new_n1155), .A2(G319), .ZN(new_n1156));
  XNOR2_X1  g730(.A(new_n1156), .B(KEYINPUT127), .ZN(new_n1157));
  NOR2_X1   g731(.A1(G229), .A2(new_n1157), .ZN(new_n1158));
  NAND4_X1  g732(.A1(new_n886), .A2(new_n1154), .A3(new_n960), .A4(new_n1158), .ZN(G225));
  INV_X1    g733(.A(G225), .ZN(G308));
endmodule


