

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X2 U552 ( .A(n528), .B(KEYINPUT90), .ZN(G164) );
  NOR2_X1 U553 ( .A1(n763), .A2(n762), .ZN(n764) );
  XOR2_X1 U554 ( .A(KEYINPUT1), .B(n530), .Z(n641) );
  NOR2_X1 U555 ( .A1(n733), .A2(n732), .ZN(n735) );
  XOR2_X1 U556 ( .A(KEYINPUT76), .B(n531), .Z(n519) );
  INV_X1 U557 ( .A(KEYINPUT26), .ZN(n703) );
  XNOR2_X1 U558 ( .A(KEYINPUT99), .B(KEYINPUT31), .ZN(n734) );
  XNOR2_X1 U559 ( .A(n735), .B(n734), .ZN(n736) );
  AND2_X1 U560 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U561 ( .A1(n697), .A2(n696), .ZN(n738) );
  NAND2_X1 U562 ( .A1(G8), .A2(n738), .ZN(n774) );
  INV_X1 U563 ( .A(KEYINPUT13), .ZN(n565) );
  NOR2_X1 U564 ( .A1(G1384), .A2(G164), .ZN(n697) );
  XNOR2_X1 U565 ( .A(n565), .B(KEYINPUT71), .ZN(n566) );
  NOR2_X1 U566 ( .A1(G2104), .A2(G2105), .ZN(n522) );
  XNOR2_X1 U567 ( .A(n567), .B(n566), .ZN(n568) );
  NOR2_X1 U568 ( .A1(G651), .A2(G543), .ZN(n647) );
  NOR2_X1 U569 ( .A1(G651), .A2(n535), .ZN(n642) );
  NAND2_X1 U570 ( .A1(n571), .A2(n570), .ZN(n929) );
  XNOR2_X1 U571 ( .A(KEYINPUT7), .B(n546), .ZN(G168) );
  INV_X1 U572 ( .A(G2105), .ZN(n523) );
  NOR2_X1 U573 ( .A1(G2104), .A2(n523), .ZN(n887) );
  NAND2_X1 U574 ( .A1(G126), .A2(n887), .ZN(n521) );
  AND2_X1 U575 ( .A1(G2104), .A2(G2105), .ZN(n888) );
  NAND2_X1 U576 ( .A1(G114), .A2(n888), .ZN(n520) );
  NAND2_X1 U577 ( .A1(n521), .A2(n520), .ZN(n527) );
  XOR2_X2 U578 ( .A(KEYINPUT17), .B(n522), .Z(n884) );
  NAND2_X1 U579 ( .A1(G138), .A2(n884), .ZN(n525) );
  AND2_X1 U580 ( .A1(n523), .A2(G2104), .ZN(n883) );
  NAND2_X1 U581 ( .A1(G102), .A2(n883), .ZN(n524) );
  NAND2_X1 U582 ( .A1(n525), .A2(n524), .ZN(n526) );
  NOR2_X1 U583 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U584 ( .A(KEYINPUT0), .B(G543), .Z(n535) );
  NAND2_X1 U585 ( .A1(n642), .A2(G51), .ZN(n529) );
  XNOR2_X1 U586 ( .A(KEYINPUT77), .B(n529), .ZN(n532) );
  XOR2_X1 U587 ( .A(G651), .B(KEYINPUT64), .Z(n534) );
  NOR2_X1 U588 ( .A1(G543), .A2(n534), .ZN(n530) );
  NAND2_X1 U589 ( .A1(n641), .A2(G63), .ZN(n531) );
  NOR2_X1 U590 ( .A1(n532), .A2(n519), .ZN(n533) );
  XNOR2_X1 U591 ( .A(KEYINPUT6), .B(n533), .ZN(n545) );
  OR2_X1 U592 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X2 U593 ( .A(KEYINPUT65), .B(n536), .ZN(n640) );
  NAND2_X1 U594 ( .A1(n640), .A2(G76), .ZN(n537) );
  XNOR2_X1 U595 ( .A(KEYINPUT74), .B(n537), .ZN(n541) );
  XOR2_X1 U596 ( .A(KEYINPUT73), .B(KEYINPUT4), .Z(n539) );
  NAND2_X1 U597 ( .A1(G89), .A2(n647), .ZN(n538) );
  XNOR2_X1 U598 ( .A(n539), .B(n538), .ZN(n540) );
  NAND2_X1 U599 ( .A1(n541), .A2(n540), .ZN(n543) );
  XOR2_X1 U600 ( .A(KEYINPUT75), .B(KEYINPUT5), .Z(n542) );
  XNOR2_X1 U601 ( .A(n543), .B(n542), .ZN(n544) );
  NAND2_X1 U602 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U603 ( .A(KEYINPUT67), .B(KEYINPUT9), .ZN(n550) );
  NAND2_X1 U604 ( .A1(G77), .A2(n640), .ZN(n548) );
  NAND2_X1 U605 ( .A1(G90), .A2(n647), .ZN(n547) );
  NAND2_X1 U606 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U607 ( .A(n550), .B(n549), .ZN(n555) );
  NAND2_X1 U608 ( .A1(n642), .A2(G52), .ZN(n551) );
  XNOR2_X1 U609 ( .A(n551), .B(KEYINPUT66), .ZN(n553) );
  NAND2_X1 U610 ( .A1(G64), .A2(n641), .ZN(n552) );
  NAND2_X1 U611 ( .A1(n553), .A2(n552), .ZN(n554) );
  NOR2_X1 U612 ( .A1(n555), .A2(n554), .ZN(G171) );
  INV_X1 U613 ( .A(G132), .ZN(G219) );
  INV_X1 U614 ( .A(G82), .ZN(G220) );
  INV_X1 U615 ( .A(G57), .ZN(G237) );
  XOR2_X1 U616 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U617 ( .A1(G94), .A2(G452), .ZN(n556) );
  XOR2_X1 U618 ( .A(KEYINPUT68), .B(n556), .Z(G173) );
  NAND2_X1 U619 ( .A1(G7), .A2(G661), .ZN(n557) );
  XNOR2_X1 U620 ( .A(n557), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U621 ( .A(G223), .B(KEYINPUT69), .ZN(n827) );
  NAND2_X1 U622 ( .A1(n827), .A2(G567), .ZN(n558) );
  XOR2_X1 U623 ( .A(KEYINPUT11), .B(n558), .Z(G234) );
  NAND2_X1 U624 ( .A1(n641), .A2(G56), .ZN(n559) );
  XOR2_X1 U625 ( .A(KEYINPUT14), .B(n559), .Z(n569) );
  NAND2_X1 U626 ( .A1(n647), .A2(G81), .ZN(n560) );
  XOR2_X1 U627 ( .A(KEYINPUT12), .B(n560), .Z(n564) );
  NAND2_X1 U628 ( .A1(n640), .A2(G68), .ZN(n562) );
  INV_X1 U629 ( .A(KEYINPUT70), .ZN(n561) );
  XNOR2_X1 U630 ( .A(n562), .B(n561), .ZN(n563) );
  NOR2_X1 U631 ( .A1(n564), .A2(n563), .ZN(n567) );
  NOR2_X1 U632 ( .A1(n569), .A2(n568), .ZN(n571) );
  NAND2_X1 U633 ( .A1(n642), .A2(G43), .ZN(n570) );
  INV_X1 U634 ( .A(G860), .ZN(n590) );
  OR2_X1 U635 ( .A1(n929), .A2(n590), .ZN(G153) );
  XOR2_X1 U636 ( .A(G171), .B(KEYINPUT72), .Z(G301) );
  NAND2_X1 U637 ( .A1(G868), .A2(G301), .ZN(n580) );
  NAND2_X1 U638 ( .A1(G92), .A2(n647), .ZN(n573) );
  NAND2_X1 U639 ( .A1(G54), .A2(n642), .ZN(n572) );
  NAND2_X1 U640 ( .A1(n573), .A2(n572), .ZN(n577) );
  NAND2_X1 U641 ( .A1(G66), .A2(n641), .ZN(n575) );
  NAND2_X1 U642 ( .A1(G79), .A2(n640), .ZN(n574) );
  NAND2_X1 U643 ( .A1(n575), .A2(n574), .ZN(n576) );
  NOR2_X1 U644 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n578), .B(KEYINPUT15), .ZN(n914) );
  INV_X1 U646 ( .A(G868), .ZN(n658) );
  NAND2_X1 U647 ( .A1(n914), .A2(n658), .ZN(n579) );
  NAND2_X1 U648 ( .A1(n580), .A2(n579), .ZN(G284) );
  NAND2_X1 U649 ( .A1(G78), .A2(n640), .ZN(n582) );
  NAND2_X1 U650 ( .A1(G53), .A2(n642), .ZN(n581) );
  NAND2_X1 U651 ( .A1(n582), .A2(n581), .ZN(n586) );
  NAND2_X1 U652 ( .A1(G65), .A2(n641), .ZN(n584) );
  NAND2_X1 U653 ( .A1(G91), .A2(n647), .ZN(n583) );
  NAND2_X1 U654 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X1 U655 ( .A1(n586), .A2(n585), .ZN(n918) );
  INV_X1 U656 ( .A(n918), .ZN(G299) );
  NOR2_X1 U657 ( .A1(G286), .A2(n658), .ZN(n587) );
  XNOR2_X1 U658 ( .A(n587), .B(KEYINPUT78), .ZN(n589) );
  NOR2_X1 U659 ( .A1(G299), .A2(G868), .ZN(n588) );
  NOR2_X1 U660 ( .A1(n589), .A2(n588), .ZN(G297) );
  NAND2_X1 U661 ( .A1(n590), .A2(G559), .ZN(n591) );
  INV_X1 U662 ( .A(n914), .ZN(n617) );
  NAND2_X1 U663 ( .A1(n591), .A2(n617), .ZN(n592) );
  XNOR2_X1 U664 ( .A(n592), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U665 ( .A1(G868), .A2(n929), .ZN(n593) );
  XOR2_X1 U666 ( .A(KEYINPUT79), .B(n593), .Z(n597) );
  NAND2_X1 U667 ( .A1(n617), .A2(G868), .ZN(n594) );
  NOR2_X1 U668 ( .A1(G559), .A2(n594), .ZN(n595) );
  XNOR2_X1 U669 ( .A(KEYINPUT80), .B(n595), .ZN(n596) );
  NOR2_X1 U670 ( .A1(n597), .A2(n596), .ZN(G282) );
  XNOR2_X1 U671 ( .A(G2096), .B(KEYINPUT82), .ZN(n606) );
  NAND2_X1 U672 ( .A1(G123), .A2(n887), .ZN(n598) );
  XNOR2_X1 U673 ( .A(n598), .B(KEYINPUT18), .ZN(n605) );
  NAND2_X1 U674 ( .A1(G111), .A2(n888), .ZN(n600) );
  NAND2_X1 U675 ( .A1(G99), .A2(n883), .ZN(n599) );
  NAND2_X1 U676 ( .A1(n600), .A2(n599), .ZN(n603) );
  NAND2_X1 U677 ( .A1(G135), .A2(n884), .ZN(n601) );
  XNOR2_X1 U678 ( .A(KEYINPUT81), .B(n601), .ZN(n602) );
  NOR2_X1 U679 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U680 ( .A1(n605), .A2(n604), .ZN(n970) );
  XNOR2_X1 U681 ( .A(n606), .B(n970), .ZN(n607) );
  NOR2_X1 U682 ( .A1(G2100), .A2(n607), .ZN(n608) );
  XNOR2_X1 U683 ( .A(KEYINPUT83), .B(n608), .ZN(G156) );
  NAND2_X1 U684 ( .A1(G80), .A2(n640), .ZN(n609) );
  XNOR2_X1 U685 ( .A(n609), .B(KEYINPUT84), .ZN(n616) );
  NAND2_X1 U686 ( .A1(G93), .A2(n647), .ZN(n611) );
  NAND2_X1 U687 ( .A1(G55), .A2(n642), .ZN(n610) );
  NAND2_X1 U688 ( .A1(n611), .A2(n610), .ZN(n614) );
  NAND2_X1 U689 ( .A1(G67), .A2(n641), .ZN(n612) );
  XNOR2_X1 U690 ( .A(KEYINPUT85), .B(n612), .ZN(n613) );
  NOR2_X1 U691 ( .A1(n614), .A2(n613), .ZN(n615) );
  NAND2_X1 U692 ( .A1(n616), .A2(n615), .ZN(n659) );
  NAND2_X1 U693 ( .A1(n617), .A2(G559), .ZN(n656) );
  XNOR2_X1 U694 ( .A(n929), .B(n656), .ZN(n618) );
  NOR2_X1 U695 ( .A1(G860), .A2(n618), .ZN(n619) );
  XOR2_X1 U696 ( .A(n659), .B(n619), .Z(G145) );
  NAND2_X1 U697 ( .A1(G86), .A2(n647), .ZN(n620) );
  XNOR2_X1 U698 ( .A(n620), .B(KEYINPUT86), .ZN(n627) );
  NAND2_X1 U699 ( .A1(G61), .A2(n641), .ZN(n622) );
  NAND2_X1 U700 ( .A1(G48), .A2(n642), .ZN(n621) );
  NAND2_X1 U701 ( .A1(n622), .A2(n621), .ZN(n625) );
  NAND2_X1 U702 ( .A1(n640), .A2(G73), .ZN(n623) );
  XOR2_X1 U703 ( .A(KEYINPUT2), .B(n623), .Z(n624) );
  NOR2_X1 U704 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U705 ( .A1(n627), .A2(n626), .ZN(G305) );
  NAND2_X1 U706 ( .A1(G87), .A2(n535), .ZN(n629) );
  NAND2_X1 U707 ( .A1(G74), .A2(G651), .ZN(n628) );
  NAND2_X1 U708 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U709 ( .A1(n641), .A2(n630), .ZN(n632) );
  NAND2_X1 U710 ( .A1(n642), .A2(G49), .ZN(n631) );
  NAND2_X1 U711 ( .A1(n632), .A2(n631), .ZN(G288) );
  NAND2_X1 U712 ( .A1(G62), .A2(n641), .ZN(n634) );
  NAND2_X1 U713 ( .A1(G75), .A2(n640), .ZN(n633) );
  NAND2_X1 U714 ( .A1(n634), .A2(n633), .ZN(n638) );
  NAND2_X1 U715 ( .A1(G88), .A2(n647), .ZN(n636) );
  NAND2_X1 U716 ( .A1(G50), .A2(n642), .ZN(n635) );
  NAND2_X1 U717 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U718 ( .A1(n638), .A2(n637), .ZN(n639) );
  XOR2_X1 U719 ( .A(KEYINPUT87), .B(n639), .Z(G166) );
  AND2_X1 U720 ( .A1(n640), .A2(G72), .ZN(n646) );
  NAND2_X1 U721 ( .A1(G60), .A2(n641), .ZN(n644) );
  NAND2_X1 U722 ( .A1(G47), .A2(n642), .ZN(n643) );
  NAND2_X1 U723 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U724 ( .A1(n646), .A2(n645), .ZN(n649) );
  NAND2_X1 U725 ( .A1(n647), .A2(G85), .ZN(n648) );
  NAND2_X1 U726 ( .A1(n649), .A2(n648), .ZN(G290) );
  XNOR2_X1 U727 ( .A(KEYINPUT19), .B(G305), .ZN(n650) );
  XNOR2_X1 U728 ( .A(n650), .B(G288), .ZN(n653) );
  XNOR2_X1 U729 ( .A(G166), .B(n929), .ZN(n651) );
  XNOR2_X1 U730 ( .A(n651), .B(n659), .ZN(n652) );
  XNOR2_X1 U731 ( .A(n653), .B(n652), .ZN(n655) );
  XNOR2_X1 U732 ( .A(G290), .B(n918), .ZN(n654) );
  XNOR2_X1 U733 ( .A(n655), .B(n654), .ZN(n900) );
  XOR2_X1 U734 ( .A(n900), .B(n656), .Z(n657) );
  NAND2_X1 U735 ( .A1(G868), .A2(n657), .ZN(n661) );
  NAND2_X1 U736 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U737 ( .A1(n661), .A2(n660), .ZN(G295) );
  NAND2_X1 U738 ( .A1(G2078), .A2(G2084), .ZN(n662) );
  XOR2_X1 U739 ( .A(KEYINPUT20), .B(n662), .Z(n663) );
  NAND2_X1 U740 ( .A1(G2090), .A2(n663), .ZN(n664) );
  XNOR2_X1 U741 ( .A(KEYINPUT21), .B(n664), .ZN(n665) );
  NAND2_X1 U742 ( .A1(n665), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U743 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U744 ( .A1(G69), .A2(G120), .ZN(n666) );
  NOR2_X1 U745 ( .A1(G237), .A2(n666), .ZN(n667) );
  NAND2_X1 U746 ( .A1(G108), .A2(n667), .ZN(n833) );
  NAND2_X1 U747 ( .A1(n833), .A2(G567), .ZN(n673) );
  NOR2_X1 U748 ( .A1(G220), .A2(G219), .ZN(n668) );
  XOR2_X1 U749 ( .A(KEYINPUT22), .B(n668), .Z(n669) );
  NOR2_X1 U750 ( .A1(G218), .A2(n669), .ZN(n670) );
  NAND2_X1 U751 ( .A1(G96), .A2(n670), .ZN(n832) );
  NAND2_X1 U752 ( .A1(G2106), .A2(n832), .ZN(n671) );
  XNOR2_X1 U753 ( .A(KEYINPUT88), .B(n671), .ZN(n672) );
  NAND2_X1 U754 ( .A1(n673), .A2(n672), .ZN(n834) );
  NAND2_X1 U755 ( .A1(G483), .A2(G661), .ZN(n674) );
  NOR2_X1 U756 ( .A1(n834), .A2(n674), .ZN(n675) );
  XOR2_X1 U757 ( .A(KEYINPUT89), .B(n675), .Z(n831) );
  NAND2_X1 U758 ( .A1(n831), .A2(G36), .ZN(G176) );
  NAND2_X1 U759 ( .A1(n888), .A2(G113), .ZN(n678) );
  NAND2_X1 U760 ( .A1(G101), .A2(n883), .ZN(n676) );
  XOR2_X1 U761 ( .A(KEYINPUT23), .B(n676), .Z(n677) );
  NAND2_X1 U762 ( .A1(n678), .A2(n677), .ZN(n682) );
  NAND2_X1 U763 ( .A1(G125), .A2(n887), .ZN(n680) );
  NAND2_X1 U764 ( .A1(G137), .A2(n884), .ZN(n679) );
  NAND2_X1 U765 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U766 ( .A1(n682), .A2(n681), .ZN(G160) );
  INV_X1 U767 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U768 ( .A(KEYINPUT104), .B(KEYINPUT40), .ZN(n817) );
  NAND2_X1 U769 ( .A1(G104), .A2(n883), .ZN(n684) );
  NAND2_X1 U770 ( .A1(G140), .A2(n884), .ZN(n683) );
  NAND2_X1 U771 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U772 ( .A(KEYINPUT34), .B(n685), .ZN(n691) );
  NAND2_X1 U773 ( .A1(n887), .A2(G128), .ZN(n686) );
  XOR2_X1 U774 ( .A(KEYINPUT91), .B(n686), .Z(n688) );
  NAND2_X1 U775 ( .A1(n888), .A2(G116), .ZN(n687) );
  NAND2_X1 U776 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U777 ( .A(n689), .B(KEYINPUT35), .Z(n690) );
  NOR2_X1 U778 ( .A1(n691), .A2(n690), .ZN(n692) );
  XOR2_X1 U779 ( .A(KEYINPUT36), .B(n692), .Z(n693) );
  XOR2_X1 U780 ( .A(KEYINPUT92), .B(n693), .Z(n898) );
  XNOR2_X1 U781 ( .A(G2067), .B(KEYINPUT37), .ZN(n810) );
  NOR2_X1 U782 ( .A1(n898), .A2(n810), .ZN(n964) );
  NAND2_X1 U783 ( .A1(G160), .A2(G40), .ZN(n695) );
  NOR2_X1 U784 ( .A1(n697), .A2(n695), .ZN(n812) );
  NAND2_X1 U785 ( .A1(n964), .A2(n812), .ZN(n694) );
  XOR2_X1 U786 ( .A(KEYINPUT93), .B(n694), .Z(n808) );
  INV_X1 U787 ( .A(n808), .ZN(n800) );
  INV_X1 U788 ( .A(n695), .ZN(n696) );
  INV_X1 U789 ( .A(n738), .ZN(n722) );
  NAND2_X1 U790 ( .A1(n722), .A2(G2072), .ZN(n698) );
  XNOR2_X1 U791 ( .A(n698), .B(KEYINPUT27), .ZN(n700) );
  XNOR2_X1 U792 ( .A(G1956), .B(KEYINPUT97), .ZN(n940) );
  NOR2_X1 U793 ( .A1(n940), .A2(n722), .ZN(n699) );
  NOR2_X1 U794 ( .A1(n700), .A2(n699), .ZN(n715) );
  NOR2_X1 U795 ( .A1(n715), .A2(n918), .ZN(n702) );
  XOR2_X1 U796 ( .A(KEYINPUT98), .B(KEYINPUT28), .Z(n701) );
  XNOR2_X1 U797 ( .A(n702), .B(n701), .ZN(n719) );
  INV_X1 U798 ( .A(G1996), .ZN(n995) );
  NOR2_X1 U799 ( .A1(n738), .A2(n995), .ZN(n704) );
  XNOR2_X1 U800 ( .A(n704), .B(n703), .ZN(n706) );
  NAND2_X1 U801 ( .A1(n738), .A2(G1341), .ZN(n705) );
  NAND2_X1 U802 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U803 ( .A1(n929), .A2(n707), .ZN(n711) );
  NAND2_X1 U804 ( .A1(G1348), .A2(n738), .ZN(n709) );
  NAND2_X1 U805 ( .A1(G2067), .A2(n722), .ZN(n708) );
  NAND2_X1 U806 ( .A1(n709), .A2(n708), .ZN(n712) );
  NOR2_X1 U807 ( .A1(n914), .A2(n712), .ZN(n710) );
  OR2_X1 U808 ( .A1(n711), .A2(n710), .ZN(n714) );
  NAND2_X1 U809 ( .A1(n914), .A2(n712), .ZN(n713) );
  NAND2_X1 U810 ( .A1(n714), .A2(n713), .ZN(n717) );
  NAND2_X1 U811 ( .A1(n715), .A2(n918), .ZN(n716) );
  NAND2_X1 U812 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U813 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U814 ( .A(KEYINPUT29), .B(n720), .ZN(n721) );
  INV_X1 U815 ( .A(n721), .ZN(n727) );
  OR2_X1 U816 ( .A1(n722), .A2(G1961), .ZN(n724) );
  XNOR2_X1 U817 ( .A(KEYINPUT25), .B(G2078), .ZN(n1000) );
  NAND2_X1 U818 ( .A1(n722), .A2(n1000), .ZN(n723) );
  NAND2_X1 U819 ( .A1(n724), .A2(n723), .ZN(n731) );
  NAND2_X1 U820 ( .A1(G171), .A2(n731), .ZN(n725) );
  XNOR2_X1 U821 ( .A(n725), .B(KEYINPUT96), .ZN(n726) );
  NAND2_X1 U822 ( .A1(n727), .A2(n726), .ZN(n737) );
  NOR2_X1 U823 ( .A1(G1966), .A2(n774), .ZN(n750) );
  NOR2_X1 U824 ( .A1(G2084), .A2(n738), .ZN(n747) );
  NOR2_X1 U825 ( .A1(n750), .A2(n747), .ZN(n728) );
  NAND2_X1 U826 ( .A1(G8), .A2(n728), .ZN(n729) );
  XNOR2_X1 U827 ( .A(KEYINPUT30), .B(n729), .ZN(n730) );
  NOR2_X1 U828 ( .A1(G168), .A2(n730), .ZN(n733) );
  NOR2_X1 U829 ( .A1(G171), .A2(n731), .ZN(n732) );
  NAND2_X1 U830 ( .A1(n737), .A2(n736), .ZN(n748) );
  NAND2_X1 U831 ( .A1(n748), .A2(G286), .ZN(n745) );
  INV_X1 U832 ( .A(G8), .ZN(n743) );
  NOR2_X1 U833 ( .A1(G1971), .A2(n774), .ZN(n740) );
  NOR2_X1 U834 ( .A1(G2090), .A2(n738), .ZN(n739) );
  NOR2_X1 U835 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U836 ( .A1(n741), .A2(G303), .ZN(n742) );
  OR2_X1 U837 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U838 ( .A(n746), .B(KEYINPUT32), .ZN(n754) );
  NAND2_X1 U839 ( .A1(G8), .A2(n747), .ZN(n752) );
  INV_X1 U840 ( .A(n748), .ZN(n749) );
  NOR2_X1 U841 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U842 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U843 ( .A1(n754), .A2(n753), .ZN(n768) );
  NOR2_X1 U844 ( .A1(G1976), .A2(G288), .ZN(n760) );
  NOR2_X1 U845 ( .A1(G1971), .A2(G303), .ZN(n755) );
  NOR2_X1 U846 ( .A1(n760), .A2(n755), .ZN(n932) );
  NAND2_X1 U847 ( .A1(n768), .A2(n932), .ZN(n756) );
  NAND2_X1 U848 ( .A1(G1976), .A2(G288), .ZN(n919) );
  NAND2_X1 U849 ( .A1(n756), .A2(n919), .ZN(n757) );
  XNOR2_X1 U850 ( .A(KEYINPUT100), .B(n757), .ZN(n758) );
  NOR2_X1 U851 ( .A1(n774), .A2(n758), .ZN(n759) );
  NOR2_X1 U852 ( .A1(KEYINPUT33), .A2(n759), .ZN(n763) );
  NAND2_X1 U853 ( .A1(n760), .A2(KEYINPUT33), .ZN(n761) );
  NOR2_X1 U854 ( .A1(n761), .A2(n774), .ZN(n762) );
  XOR2_X1 U855 ( .A(G1981), .B(G305), .Z(n915) );
  NAND2_X1 U856 ( .A1(n764), .A2(n915), .ZN(n778) );
  NOR2_X1 U857 ( .A1(G2090), .A2(G303), .ZN(n765) );
  XOR2_X1 U858 ( .A(KEYINPUT101), .B(n765), .Z(n766) );
  NAND2_X1 U859 ( .A1(G8), .A2(n766), .ZN(n767) );
  NAND2_X1 U860 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U861 ( .A(n769), .B(KEYINPUT102), .ZN(n770) );
  NAND2_X1 U862 ( .A1(n770), .A2(n774), .ZN(n771) );
  XNOR2_X1 U863 ( .A(n771), .B(KEYINPUT103), .ZN(n776) );
  NOR2_X1 U864 ( .A1(G1981), .A2(G305), .ZN(n772) );
  XOR2_X1 U865 ( .A(n772), .B(KEYINPUT24), .Z(n773) );
  NOR2_X1 U866 ( .A1(n774), .A2(n773), .ZN(n775) );
  NOR2_X1 U867 ( .A1(n776), .A2(n775), .ZN(n777) );
  NAND2_X1 U868 ( .A1(n778), .A2(n777), .ZN(n798) );
  NAND2_X1 U869 ( .A1(G107), .A2(n888), .ZN(n779) );
  XOR2_X1 U870 ( .A(KEYINPUT94), .B(n779), .Z(n784) );
  NAND2_X1 U871 ( .A1(G95), .A2(n883), .ZN(n781) );
  NAND2_X1 U872 ( .A1(G131), .A2(n884), .ZN(n780) );
  NAND2_X1 U873 ( .A1(n781), .A2(n780), .ZN(n782) );
  XOR2_X1 U874 ( .A(KEYINPUT95), .B(n782), .Z(n783) );
  NOR2_X1 U875 ( .A1(n784), .A2(n783), .ZN(n786) );
  NAND2_X1 U876 ( .A1(n887), .A2(G119), .ZN(n785) );
  NAND2_X1 U877 ( .A1(n786), .A2(n785), .ZN(n874) );
  AND2_X1 U878 ( .A1(n874), .A2(G1991), .ZN(n795) );
  NAND2_X1 U879 ( .A1(G129), .A2(n887), .ZN(n788) );
  NAND2_X1 U880 ( .A1(G117), .A2(n888), .ZN(n787) );
  NAND2_X1 U881 ( .A1(n788), .A2(n787), .ZN(n791) );
  NAND2_X1 U882 ( .A1(n883), .A2(G105), .ZN(n789) );
  XOR2_X1 U883 ( .A(KEYINPUT38), .B(n789), .Z(n790) );
  NOR2_X1 U884 ( .A1(n791), .A2(n790), .ZN(n793) );
  NAND2_X1 U885 ( .A1(n884), .A2(G141), .ZN(n792) );
  NAND2_X1 U886 ( .A1(n793), .A2(n792), .ZN(n876) );
  AND2_X1 U887 ( .A1(G1996), .A2(n876), .ZN(n794) );
  NOR2_X1 U888 ( .A1(n795), .A2(n794), .ZN(n975) );
  INV_X1 U889 ( .A(n812), .ZN(n796) );
  NOR2_X1 U890 ( .A1(n975), .A2(n796), .ZN(n805) );
  INV_X1 U891 ( .A(n805), .ZN(n797) );
  NAND2_X1 U892 ( .A1(n798), .A2(n797), .ZN(n799) );
  NOR2_X1 U893 ( .A1(n800), .A2(n799), .ZN(n802) );
  XNOR2_X1 U894 ( .A(G1986), .B(G290), .ZN(n926) );
  NAND2_X1 U895 ( .A1(n926), .A2(n812), .ZN(n801) );
  NAND2_X1 U896 ( .A1(n802), .A2(n801), .ZN(n815) );
  NOR2_X1 U897 ( .A1(G1996), .A2(n876), .ZN(n968) );
  NOR2_X1 U898 ( .A1(G1986), .A2(G290), .ZN(n803) );
  NOR2_X1 U899 ( .A1(G1991), .A2(n874), .ZN(n973) );
  NOR2_X1 U900 ( .A1(n803), .A2(n973), .ZN(n804) );
  NOR2_X1 U901 ( .A1(n805), .A2(n804), .ZN(n806) );
  NOR2_X1 U902 ( .A1(n968), .A2(n806), .ZN(n807) );
  XNOR2_X1 U903 ( .A(n807), .B(KEYINPUT39), .ZN(n809) );
  NAND2_X1 U904 ( .A1(n809), .A2(n808), .ZN(n811) );
  NAND2_X1 U905 ( .A1(n898), .A2(n810), .ZN(n966) );
  NAND2_X1 U906 ( .A1(n811), .A2(n966), .ZN(n813) );
  NAND2_X1 U907 ( .A1(n813), .A2(n812), .ZN(n814) );
  NAND2_X1 U908 ( .A1(n815), .A2(n814), .ZN(n816) );
  XNOR2_X1 U909 ( .A(n817), .B(n816), .ZN(G329) );
  XNOR2_X1 U910 ( .A(G1348), .B(G2454), .ZN(n818) );
  XNOR2_X1 U911 ( .A(n818), .B(G2430), .ZN(n819) );
  XNOR2_X1 U912 ( .A(n819), .B(G1341), .ZN(n825) );
  XOR2_X1 U913 ( .A(G2443), .B(G2427), .Z(n821) );
  XNOR2_X1 U914 ( .A(G2438), .B(G2446), .ZN(n820) );
  XNOR2_X1 U915 ( .A(n821), .B(n820), .ZN(n823) );
  XOR2_X1 U916 ( .A(G2451), .B(G2435), .Z(n822) );
  XNOR2_X1 U917 ( .A(n823), .B(n822), .ZN(n824) );
  XNOR2_X1 U918 ( .A(n825), .B(n824), .ZN(n826) );
  NAND2_X1 U919 ( .A1(n826), .A2(G14), .ZN(n905) );
  XNOR2_X1 U920 ( .A(KEYINPUT105), .B(n905), .ZN(G401) );
  NAND2_X1 U921 ( .A1(n827), .A2(G2106), .ZN(n828) );
  XNOR2_X1 U922 ( .A(n828), .B(KEYINPUT106), .ZN(G217) );
  AND2_X1 U923 ( .A1(G15), .A2(G2), .ZN(n829) );
  NAND2_X1 U924 ( .A1(G661), .A2(n829), .ZN(G259) );
  NAND2_X1 U925 ( .A1(G3), .A2(G1), .ZN(n830) );
  NAND2_X1 U926 ( .A1(n831), .A2(n830), .ZN(G188) );
  INV_X1 U928 ( .A(G120), .ZN(G236) );
  INV_X1 U929 ( .A(G96), .ZN(G221) );
  INV_X1 U930 ( .A(G69), .ZN(G235) );
  NOR2_X1 U931 ( .A1(n833), .A2(n832), .ZN(G325) );
  INV_X1 U932 ( .A(G325), .ZN(G261) );
  INV_X1 U933 ( .A(n834), .ZN(G319) );
  XNOR2_X1 U934 ( .A(G1991), .B(KEYINPUT41), .ZN(n844) );
  XOR2_X1 U935 ( .A(G1961), .B(G1956), .Z(n836) );
  XNOR2_X1 U936 ( .A(G1996), .B(G1986), .ZN(n835) );
  XNOR2_X1 U937 ( .A(n836), .B(n835), .ZN(n840) );
  XOR2_X1 U938 ( .A(G1966), .B(G1971), .Z(n838) );
  XNOR2_X1 U939 ( .A(G1981), .B(G1976), .ZN(n837) );
  XNOR2_X1 U940 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U941 ( .A(n840), .B(n839), .Z(n842) );
  XNOR2_X1 U942 ( .A(KEYINPUT108), .B(G2474), .ZN(n841) );
  XNOR2_X1 U943 ( .A(n842), .B(n841), .ZN(n843) );
  XNOR2_X1 U944 ( .A(n844), .B(n843), .ZN(G229) );
  XOR2_X1 U945 ( .A(KEYINPUT42), .B(G2090), .Z(n846) );
  XNOR2_X1 U946 ( .A(G2067), .B(G2084), .ZN(n845) );
  XNOR2_X1 U947 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U948 ( .A(n847), .B(G2100), .Z(n849) );
  XNOR2_X1 U949 ( .A(G2072), .B(G2078), .ZN(n848) );
  XNOR2_X1 U950 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U951 ( .A(G2096), .B(KEYINPUT43), .Z(n851) );
  XNOR2_X1 U952 ( .A(G2678), .B(KEYINPUT107), .ZN(n850) );
  XNOR2_X1 U953 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U954 ( .A(n853), .B(n852), .Z(G227) );
  NAND2_X1 U955 ( .A1(G112), .A2(n888), .ZN(n854) );
  XNOR2_X1 U956 ( .A(n854), .B(KEYINPUT110), .ZN(n860) );
  NAND2_X1 U957 ( .A1(G124), .A2(n887), .ZN(n855) );
  XOR2_X1 U958 ( .A(KEYINPUT44), .B(n855), .Z(n858) );
  NAND2_X1 U959 ( .A1(G100), .A2(n883), .ZN(n856) );
  XNOR2_X1 U960 ( .A(KEYINPUT111), .B(n856), .ZN(n857) );
  NOR2_X1 U961 ( .A1(n858), .A2(n857), .ZN(n859) );
  NAND2_X1 U962 ( .A1(n860), .A2(n859), .ZN(n863) );
  NAND2_X1 U963 ( .A1(G136), .A2(n884), .ZN(n861) );
  XNOR2_X1 U964 ( .A(KEYINPUT109), .B(n861), .ZN(n862) );
  NOR2_X1 U965 ( .A1(n863), .A2(n862), .ZN(G162) );
  NAND2_X1 U966 ( .A1(G106), .A2(n883), .ZN(n865) );
  NAND2_X1 U967 ( .A1(G142), .A2(n884), .ZN(n864) );
  NAND2_X1 U968 ( .A1(n865), .A2(n864), .ZN(n866) );
  XNOR2_X1 U969 ( .A(n866), .B(KEYINPUT45), .ZN(n868) );
  NAND2_X1 U970 ( .A1(G130), .A2(n887), .ZN(n867) );
  NAND2_X1 U971 ( .A1(n868), .A2(n867), .ZN(n871) );
  NAND2_X1 U972 ( .A1(n888), .A2(G118), .ZN(n869) );
  XOR2_X1 U973 ( .A(KEYINPUT112), .B(n869), .Z(n870) );
  NOR2_X1 U974 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U975 ( .A(n872), .B(G164), .ZN(n873) );
  XNOR2_X1 U976 ( .A(n873), .B(n970), .ZN(n875) );
  XNOR2_X1 U977 ( .A(n875), .B(n874), .ZN(n878) );
  XOR2_X1 U978 ( .A(G160), .B(n876), .Z(n877) );
  XNOR2_X1 U979 ( .A(n878), .B(n877), .ZN(n882) );
  XOR2_X1 U980 ( .A(KEYINPUT46), .B(KEYINPUT114), .Z(n880) );
  XNOR2_X1 U981 ( .A(KEYINPUT115), .B(KEYINPUT48), .ZN(n879) );
  XNOR2_X1 U982 ( .A(n880), .B(n879), .ZN(n881) );
  XOR2_X1 U983 ( .A(n882), .B(n881), .Z(n896) );
  NAND2_X1 U984 ( .A1(G103), .A2(n883), .ZN(n886) );
  NAND2_X1 U985 ( .A1(G139), .A2(n884), .ZN(n885) );
  NAND2_X1 U986 ( .A1(n886), .A2(n885), .ZN(n894) );
  NAND2_X1 U987 ( .A1(G127), .A2(n887), .ZN(n890) );
  NAND2_X1 U988 ( .A1(G115), .A2(n888), .ZN(n889) );
  NAND2_X1 U989 ( .A1(n890), .A2(n889), .ZN(n891) );
  XNOR2_X1 U990 ( .A(KEYINPUT47), .B(n891), .ZN(n892) );
  XNOR2_X1 U991 ( .A(KEYINPUT113), .B(n892), .ZN(n893) );
  NOR2_X1 U992 ( .A1(n894), .A2(n893), .ZN(n976) );
  XNOR2_X1 U993 ( .A(n976), .B(G162), .ZN(n895) );
  XNOR2_X1 U994 ( .A(n896), .B(n895), .ZN(n897) );
  XOR2_X1 U995 ( .A(n898), .B(n897), .Z(n899) );
  NOR2_X1 U996 ( .A1(G37), .A2(n899), .ZN(G395) );
  XOR2_X1 U997 ( .A(KEYINPUT116), .B(n900), .Z(n902) );
  XNOR2_X1 U998 ( .A(G171), .B(G286), .ZN(n901) );
  XNOR2_X1 U999 ( .A(n902), .B(n901), .ZN(n903) );
  XNOR2_X1 U1000 ( .A(n903), .B(n914), .ZN(n904) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n904), .ZN(G397) );
  NAND2_X1 U1002 ( .A1(n905), .A2(G319), .ZN(n906) );
  XNOR2_X1 U1003 ( .A(n906), .B(KEYINPUT117), .ZN(n909) );
  NOR2_X1 U1004 ( .A1(G229), .A2(G227), .ZN(n907) );
  XOR2_X1 U1005 ( .A(KEYINPUT49), .B(n907), .Z(n908) );
  NAND2_X1 U1006 ( .A1(n909), .A2(n908), .ZN(n912) );
  NOR2_X1 U1007 ( .A1(G395), .A2(G397), .ZN(n910) );
  XOR2_X1 U1008 ( .A(KEYINPUT118), .B(n910), .Z(n911) );
  NOR2_X1 U1009 ( .A1(n912), .A2(n911), .ZN(n913) );
  XNOR2_X1 U1010 ( .A(KEYINPUT119), .B(n913), .ZN(G225) );
  INV_X1 U1011 ( .A(G225), .ZN(G308) );
  INV_X1 U1012 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1013 ( .A(KEYINPUT56), .B(G16), .Z(n937) );
  XNOR2_X1 U1014 ( .A(G1348), .B(n914), .ZN(n935) );
  XNOR2_X1 U1015 ( .A(G1966), .B(G168), .ZN(n916) );
  NAND2_X1 U1016 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1017 ( .A(n917), .B(KEYINPUT57), .ZN(n928) );
  XNOR2_X1 U1018 ( .A(G1956), .B(n918), .ZN(n920) );
  NAND2_X1 U1019 ( .A1(n920), .A2(n919), .ZN(n922) );
  XOR2_X1 U1020 ( .A(G171), .B(G1961), .Z(n921) );
  NOR2_X1 U1021 ( .A1(n922), .A2(n921), .ZN(n924) );
  NAND2_X1 U1022 ( .A1(G1971), .A2(G303), .ZN(n923) );
  NAND2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n925) );
  NOR2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n931) );
  XNOR2_X1 U1026 ( .A(G1341), .B(n929), .ZN(n930) );
  NOR2_X1 U1027 ( .A1(n931), .A2(n930), .ZN(n933) );
  NAND2_X1 U1028 ( .A1(n933), .A2(n932), .ZN(n934) );
  NOR2_X1 U1029 ( .A1(n935), .A2(n934), .ZN(n936) );
  NOR2_X1 U1030 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1031 ( .A(KEYINPUT125), .B(n938), .ZN(n994) );
  XOR2_X1 U1032 ( .A(G16), .B(KEYINPUT126), .Z(n962) );
  XNOR2_X1 U1033 ( .A(KEYINPUT127), .B(G1966), .ZN(n939) );
  XNOR2_X1 U1034 ( .A(n939), .B(G21), .ZN(n952) );
  XNOR2_X1 U1035 ( .A(G20), .B(n940), .ZN(n944) );
  XNOR2_X1 U1036 ( .A(G1981), .B(G6), .ZN(n942) );
  XNOR2_X1 U1037 ( .A(G1341), .B(G19), .ZN(n941) );
  NOR2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1039 ( .A1(n944), .A2(n943), .ZN(n947) );
  XOR2_X1 U1040 ( .A(KEYINPUT59), .B(G1348), .Z(n945) );
  XNOR2_X1 U1041 ( .A(G4), .B(n945), .ZN(n946) );
  NOR2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1043 ( .A(KEYINPUT60), .B(n948), .Z(n950) );
  XNOR2_X1 U1044 ( .A(G1961), .B(G5), .ZN(n949) );
  NOR2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n959) );
  XNOR2_X1 U1047 ( .A(G1976), .B(G23), .ZN(n954) );
  XNOR2_X1 U1048 ( .A(G1971), .B(G22), .ZN(n953) );
  NOR2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n956) );
  XOR2_X1 U1050 ( .A(G1986), .B(G24), .Z(n955) );
  NAND2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1052 ( .A(KEYINPUT58), .B(n957), .ZN(n958) );
  NOR2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1054 ( .A(n960), .B(KEYINPUT61), .ZN(n961) );
  NAND2_X1 U1055 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1056 ( .A1(G11), .A2(n963), .ZN(n992) );
  INV_X1 U1057 ( .A(n964), .ZN(n965) );
  NAND2_X1 U1058 ( .A1(n966), .A2(n965), .ZN(n985) );
  XOR2_X1 U1059 ( .A(G2090), .B(G162), .Z(n967) );
  NOR2_X1 U1060 ( .A1(n968), .A2(n967), .ZN(n969) );
  XOR2_X1 U1061 ( .A(KEYINPUT51), .B(n969), .Z(n983) );
  XNOR2_X1 U1062 ( .A(G160), .B(G2084), .ZN(n971) );
  NAND2_X1 U1063 ( .A1(n971), .A2(n970), .ZN(n972) );
  NOR2_X1 U1064 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1065 ( .A1(n975), .A2(n974), .ZN(n981) );
  XOR2_X1 U1066 ( .A(G2072), .B(n976), .Z(n978) );
  XOR2_X1 U1067 ( .A(G164), .B(G2078), .Z(n977) );
  NOR2_X1 U1068 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1069 ( .A(KEYINPUT50), .B(n979), .Z(n980) );
  NOR2_X1 U1070 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1071 ( .A1(n983), .A2(n982), .ZN(n984) );
  NOR2_X1 U1072 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1073 ( .A(KEYINPUT52), .B(n986), .ZN(n988) );
  INV_X1 U1074 ( .A(KEYINPUT55), .ZN(n987) );
  NAND2_X1 U1075 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1076 ( .A1(n989), .A2(G29), .ZN(n990) );
  XOR2_X1 U1077 ( .A(KEYINPUT120), .B(n990), .Z(n991) );
  NOR2_X1 U1078 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1079 ( .A1(n994), .A2(n993), .ZN(n1019) );
  XNOR2_X1 U1080 ( .A(G32), .B(n995), .ZN(n999) );
  XNOR2_X1 U1081 ( .A(G2067), .B(G26), .ZN(n997) );
  XNOR2_X1 U1082 ( .A(G33), .B(G2072), .ZN(n996) );
  NOR2_X1 U1083 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1084 ( .A1(n999), .A2(n998), .ZN(n1003) );
  XNOR2_X1 U1085 ( .A(G27), .B(n1000), .ZN(n1001) );
  XNOR2_X1 U1086 ( .A(KEYINPUT121), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1087 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1088 ( .A(KEYINPUT122), .B(n1004), .ZN(n1005) );
  NAND2_X1 U1089 ( .A1(n1005), .A2(G28), .ZN(n1007) );
  XNOR2_X1 U1090 ( .A(G25), .B(G1991), .ZN(n1006) );
  NOR2_X1 U1091 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XOR2_X1 U1092 ( .A(KEYINPUT53), .B(n1008), .Z(n1012) );
  XNOR2_X1 U1093 ( .A(KEYINPUT54), .B(G34), .ZN(n1009) );
  XNOR2_X1 U1094 ( .A(n1009), .B(KEYINPUT123), .ZN(n1010) );
  XNOR2_X1 U1095 ( .A(G2084), .B(n1010), .ZN(n1011) );
  NAND2_X1 U1096 ( .A1(n1012), .A2(n1011), .ZN(n1014) );
  XNOR2_X1 U1097 ( .A(G35), .B(G2090), .ZN(n1013) );
  NOR2_X1 U1098 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1099 ( .A(KEYINPUT55), .B(n1015), .Z(n1017) );
  XNOR2_X1 U1100 ( .A(G29), .B(KEYINPUT124), .ZN(n1016) );
  NOR2_X1 U1101 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NOR2_X1 U1102 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1103 ( .A(n1020), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1104 ( .A(G311), .ZN(G150) );
endmodule

