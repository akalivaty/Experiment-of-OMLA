//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 0 1 0 0 0 0 0 0 0 1 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 0 1 1 0 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 1 1 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:12 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n555, new_n557, new_n558,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n621, new_n624, new_n625,
    new_n626, new_n628, new_n629, new_n630, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n866, new_n867, new_n868, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1246;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT64), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n454));
  XNOR2_X1  g029(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT66), .ZN(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  INV_X1    g034(.A(G2106), .ZN(new_n460));
  OR2_X1    g035(.A1(new_n455), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n456), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G567), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(G319));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(G101), .ZN(new_n474));
  OAI21_X1  g049(.A(KEYINPUT67), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n466), .A2(G2105), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT67), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n476), .A2(new_n477), .A3(G101), .ZN(new_n478));
  AOI22_X1  g053(.A1(new_n471), .A2(G137), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(G113), .A2(G2104), .ZN(new_n480));
  INV_X1    g055(.A(G125), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n480), .B1(new_n470), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  AND2_X1   g058(.A1(new_n479), .A2(new_n483), .ZN(G160));
  NOR2_X1   g059(.A1(new_n470), .A2(new_n472), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n471), .A2(G136), .ZN(new_n487));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G112), .C2(new_n472), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n486), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  OR2_X1    g066(.A1(G102), .A2(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n492), .B(G2104), .C1(G114), .C2(new_n472), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n467), .A2(new_n469), .A3(G126), .A4(G2105), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n467), .A2(new_n469), .A3(G138), .A4(new_n472), .ZN(new_n496));
  OR2_X1    g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n495), .B1(new_n497), .B2(new_n498), .ZN(G164));
  NAND2_X1  g074(.A1(G75), .A2(G543), .ZN(new_n500));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G62), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n500), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(G50), .A2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G88), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n508), .B1(new_n505), .B2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT68), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n511), .B1(new_n512), .B2(G651), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n514), .A2(KEYINPUT68), .A3(KEYINPUT6), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n513), .A2(new_n515), .B1(new_n512), .B2(G651), .ZN(new_n516));
  AOI22_X1  g091(.A1(G651), .A2(new_n507), .B1(new_n510), .B2(new_n516), .ZN(G166));
  INV_X1    g092(.A(KEYINPUT69), .ZN(new_n518));
  OAI21_X1  g093(.A(G543), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n513), .A2(new_n515), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n512), .A2(G651), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n520), .A2(new_n518), .A3(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G51), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT70), .B(KEYINPUT7), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n526), .B(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(G63), .A2(G651), .ZN(new_n529));
  AND3_X1   g104(.A1(new_n514), .A2(KEYINPUT68), .A3(KEYINPUT6), .ZN(new_n530));
  AOI21_X1  g105(.A(KEYINPUT68), .B1(new_n514), .B2(KEYINPUT6), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n521), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(G89), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n529), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(new_n505), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n528), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  AND2_X1   g111(.A1(new_n525), .A2(new_n536), .ZN(G168));
  NAND2_X1  g112(.A1(new_n524), .A2(G52), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n532), .A2(new_n505), .ZN(new_n539));
  NAND2_X1  g114(.A1(G77), .A2(G543), .ZN(new_n540));
  INV_X1    g115(.A(G64), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n505), .B2(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n539), .A2(G90), .B1(G651), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n538), .A2(new_n543), .ZN(G301));
  INV_X1    g119(.A(G301), .ZN(G171));
  NAND2_X1  g120(.A1(G68), .A2(G543), .ZN(new_n546));
  INV_X1    g121(.A(G56), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n505), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G651), .ZN(new_n549));
  INV_X1    g124(.A(G81), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n516), .A2(new_n535), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n552), .B1(G43), .B2(new_n524), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  AND3_X1   g129(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G36), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n555), .A2(new_n558), .ZN(G188));
  NAND2_X1  g134(.A1(new_n532), .A2(KEYINPUT69), .ZN(new_n560));
  NAND4_X1  g135(.A1(new_n560), .A2(G53), .A3(G543), .A4(new_n522), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(KEYINPUT9), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n501), .B1(new_n532), .B2(KEYINPUT69), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n563), .A2(new_n564), .A3(G53), .A4(new_n522), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  INV_X1    g142(.A(G65), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n505), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G651), .ZN(new_n570));
  INV_X1    g145(.A(G91), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n571), .B2(new_n551), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n566), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(KEYINPUT71), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT71), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n566), .A2(new_n576), .A3(new_n573), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n575), .A2(new_n577), .ZN(G299));
  NAND2_X1  g153(.A1(new_n525), .A2(new_n536), .ZN(G286));
  INV_X1    g154(.A(G166), .ZN(G303));
  NAND3_X1  g155(.A1(new_n563), .A2(G49), .A3(new_n522), .ZN(new_n581));
  INV_X1    g156(.A(G74), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n514), .B1(new_n505), .B2(new_n582), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n583), .B1(new_n539), .B2(G87), .ZN(new_n584));
  AND2_X1   g159(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(G288));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G61), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n505), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(G651), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(KEYINPUT72), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT72), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n589), .A2(new_n592), .A3(G651), .ZN(new_n593));
  NAND2_X1  g168(.A1(G48), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G86), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n505), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(new_n516), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n591), .A2(new_n593), .A3(new_n597), .ZN(G305));
  NAND2_X1  g173(.A1(G72), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G60), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n505), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(G651), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT73), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n603), .B1(G85), .B2(new_n539), .ZN(new_n604));
  XOR2_X1   g179(.A(KEYINPUT74), .B(G47), .Z(new_n605));
  NAND2_X1  g180(.A1(new_n524), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n604), .A2(new_n606), .ZN(G290));
  NAND2_X1  g182(.A1(G301), .A2(G868), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n516), .A2(G92), .A3(new_n535), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT10), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n609), .B(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n524), .A2(G54), .ZN(new_n612));
  AND2_X1   g187(.A1(new_n535), .A2(G66), .ZN(new_n613));
  NAND2_X1  g188(.A1(G79), .A2(G543), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT75), .ZN(new_n615));
  OAI21_X1  g190(.A(G651), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  AND3_X1   g191(.A1(new_n611), .A2(new_n612), .A3(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n608), .B1(new_n617), .B2(G868), .ZN(G284));
  OAI21_X1  g193(.A(new_n608), .B1(new_n617), .B2(G868), .ZN(G321));
  INV_X1    g194(.A(G868), .ZN(new_n620));
  NAND2_X1  g195(.A1(G299), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(new_n620), .B2(G168), .ZN(G297));
  OAI21_X1  g197(.A(new_n621), .B1(new_n620), .B2(G168), .ZN(G280));
  INV_X1    g198(.A(new_n617), .ZN(new_n624));
  INV_X1    g199(.A(G860), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n624), .B1(G559), .B2(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT76), .ZN(G148));
  INV_X1    g202(.A(new_n553), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(new_n620), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n624), .A2(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n629), .B1(new_n630), .B2(new_n620), .ZN(G323));
  XNOR2_X1  g206(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g207(.A1(new_n485), .A2(G123), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n471), .A2(G135), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n472), .A2(G111), .ZN(new_n635));
  OAI21_X1  g210(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n633), .B(new_n634), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(G2096), .Z(new_n638));
  NOR2_X1   g213(.A1(new_n470), .A2(new_n473), .ZN(new_n639));
  XOR2_X1   g214(.A(KEYINPUT77), .B(KEYINPUT12), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(KEYINPUT13), .B(G2100), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n638), .A2(new_n643), .ZN(G156));
  XNOR2_X1  g219(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n645));
  INV_X1    g220(.A(G1348), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2451), .B(G2454), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(G1341), .ZN(new_n650));
  INV_X1    g225(.A(KEYINPUT14), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT15), .B(G2435), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2438), .ZN(new_n653));
  XOR2_X1   g228(.A(G2427), .B(G2430), .Z(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n651), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n656), .A2(KEYINPUT79), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(KEYINPUT79), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n653), .A2(new_n655), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n650), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  AOI211_X1 g237(.A(G1341), .B(new_n660), .C1(new_n657), .C2(new_n658), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n649), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(new_n658), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n656), .A2(KEYINPUT79), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n661), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n667), .A2(G1341), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n659), .A2(new_n650), .A3(new_n661), .ZN(new_n669));
  INV_X1    g244(.A(new_n649), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n668), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2443), .B(G2446), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n664), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n673), .A2(G14), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n672), .B1(new_n664), .B2(new_n671), .ZN(new_n675));
  OAI21_X1  g250(.A(KEYINPUT80), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n675), .ZN(new_n677));
  INV_X1    g252(.A(KEYINPUT80), .ZN(new_n678));
  NAND4_X1  g253(.A1(new_n677), .A2(new_n678), .A3(G14), .A4(new_n673), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(G401));
  XOR2_X1   g256(.A(G2084), .B(G2090), .Z(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G2067), .B(G2678), .Z(new_n684));
  NOR2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G2072), .B(G2078), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT18), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n683), .A2(new_n684), .ZN(new_n689));
  AND3_X1   g264(.A1(new_n689), .A2(KEYINPUT17), .A3(new_n686), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n686), .B1(new_n689), .B2(KEYINPUT17), .ZN(new_n691));
  NOR3_X1   g266(.A1(new_n690), .A2(new_n691), .A3(new_n685), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G2096), .B(G2100), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(G227));
  XNOR2_X1  g270(.A(G1971), .B(G1976), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT81), .B(KEYINPUT19), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1956), .B(G2474), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1961), .B(G1966), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n698), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n699), .B(new_n700), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n699), .A2(new_n700), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n698), .A2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT20), .ZN(new_n705));
  OAI221_X1 g280(.A(new_n701), .B1(new_n698), .B2(new_n702), .C1(new_n704), .C2(new_n705), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(new_n705), .B2(new_n704), .ZN(new_n707));
  INV_X1    g282(.A(G1991), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n707), .A2(new_n708), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(G1996), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  AOI21_X1  g289(.A(G1996), .B1(new_n709), .B2(new_n710), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(G1981), .B(G1986), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n714), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n717), .B1(new_n713), .B2(new_n715), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n721));
  AND3_X1   g296(.A1(new_n719), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n721), .B1(new_n719), .B2(new_n720), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(G229));
  INV_X1    g300(.A(G16), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G24), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT83), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(G290), .B2(G16), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(G1986), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n485), .A2(G119), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n471), .A2(G131), .ZN(new_n732));
  OR2_X1    g307(.A1(G95), .A2(G2105), .ZN(new_n733));
  OAI211_X1 g308(.A(new_n733), .B(G2104), .C1(G107), .C2(new_n472), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n731), .A2(new_n732), .A3(new_n734), .ZN(new_n735));
  MUX2_X1   g310(.A(G25), .B(new_n735), .S(G29), .Z(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT82), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT35), .B(G1991), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n730), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n726), .A2(G6), .ZN(new_n741));
  INV_X1    g316(.A(G305), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n741), .B1(new_n742), .B2(new_n726), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT32), .B(G1981), .ZN(new_n744));
  AND2_X1   g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n743), .A2(new_n744), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n726), .A2(G22), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G166), .B2(new_n726), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G1971), .ZN(new_n749));
  OR3_X1    g324(.A1(new_n745), .A2(new_n746), .A3(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT34), .ZN(new_n751));
  NOR2_X1   g326(.A1(G16), .A2(G23), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(new_n585), .B2(G16), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT33), .B(G1976), .Z(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  OR3_X1    g330(.A1(new_n750), .A2(new_n751), .A3(new_n755), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n751), .B1(new_n750), .B2(new_n755), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n740), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT84), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(KEYINPUT36), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT85), .Z(new_n761));
  NAND2_X1  g336(.A1(new_n758), .A2(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(G28), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n763), .A2(KEYINPUT30), .ZN(new_n764));
  AOI21_X1  g339(.A(G29), .B1(new_n763), .B2(KEYINPUT30), .ZN(new_n765));
  OR2_X1    g340(.A1(KEYINPUT31), .A2(G11), .ZN(new_n766));
  NAND2_X1  g341(.A1(KEYINPUT31), .A2(G11), .ZN(new_n767));
  AOI22_X1  g342(.A1(new_n764), .A2(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(G29), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n768), .B1(new_n637), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n485), .A2(G129), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n471), .A2(G141), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n476), .A2(G105), .ZN(new_n773));
  NAND3_X1  g348(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT26), .Z(new_n775));
  NAND4_X1  g350(.A1(new_n771), .A2(new_n772), .A3(new_n773), .A4(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n777), .A2(G29), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G29), .B2(G32), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT27), .B(G1996), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n770), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(G2084), .ZN(new_n782));
  NOR2_X1   g357(.A1(G160), .A2(new_n769), .ZN(new_n783));
  NAND2_X1  g358(.A1(KEYINPUT24), .A2(G34), .ZN(new_n784));
  NOR2_X1   g359(.A1(KEYINPUT24), .A2(G34), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n785), .A2(G29), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n783), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  OAI221_X1 g362(.A(new_n781), .B1(new_n782), .B2(new_n787), .C1(new_n779), .C2(new_n780), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n769), .A2(G35), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G162), .B2(new_n769), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT29), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n788), .B1(G2090), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n787), .A2(new_n782), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT93), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n791), .A2(G2090), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n476), .A2(G103), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n797), .A2(KEYINPUT88), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(KEYINPUT88), .ZN(new_n799));
  AND3_X1   g374(.A1(new_n798), .A2(KEYINPUT25), .A3(new_n799), .ZN(new_n800));
  AOI21_X1  g375(.A(KEYINPUT25), .B1(new_n798), .B2(new_n799), .ZN(new_n801));
  AND2_X1   g376(.A1(new_n471), .A2(G139), .ZN(new_n802));
  NOR3_X1   g377(.A1(new_n800), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(G115), .A2(G2104), .ZN(new_n804));
  INV_X1    g379(.A(G127), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n804), .B1(new_n470), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n806), .A2(G2105), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT89), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n803), .A2(new_n809), .ZN(new_n810));
  MUX2_X1   g385(.A(G33), .B(new_n810), .S(G29), .Z(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(G2072), .Z(new_n812));
  NOR2_X1   g387(.A1(G27), .A2(G29), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(G164), .B2(G29), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT94), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(G2078), .ZN(new_n816));
  NAND4_X1  g391(.A1(new_n792), .A2(new_n796), .A3(new_n812), .A4(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n769), .A2(G26), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT28), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n485), .A2(G128), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n471), .A2(G140), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n472), .A2(G116), .ZN(new_n822));
  OAI21_X1  g397(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n823));
  OAI211_X1 g398(.A(new_n820), .B(new_n821), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(G29), .ZN(new_n825));
  AND2_X1   g400(.A1(new_n825), .A2(KEYINPUT87), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n825), .A2(KEYINPUT87), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n819), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(G2067), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n726), .A2(G21), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(G168), .B2(new_n726), .ZN(new_n832));
  INV_X1    g407(.A(G1966), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  OAI211_X1 g409(.A(new_n830), .B(new_n834), .C1(G2078), .C2(new_n815), .ZN(new_n835));
  NOR2_X1   g410(.A1(G5), .A2(G16), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT90), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(G301), .B2(new_n726), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT91), .ZN(new_n839));
  INV_X1    g414(.A(G1961), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n726), .A2(G4), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n842), .B1(new_n617), .B2(new_n726), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(new_n646), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  NOR3_X1   g420(.A1(new_n817), .A2(new_n835), .A3(new_n845), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n839), .A2(new_n840), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT92), .ZN(new_n848));
  OR2_X1    g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n726), .A2(G19), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n850), .B1(new_n553), .B2(new_n726), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT86), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(G1341), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n847), .A2(new_n848), .ZN(new_n854));
  AND3_X1   g429(.A1(new_n849), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n762), .A2(new_n846), .A3(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT23), .ZN(new_n857));
  AND3_X1   g432(.A1(new_n857), .A2(new_n726), .A3(G20), .ZN(new_n858));
  NAND2_X1  g433(.A1(G299), .A2(G16), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n857), .B1(new_n726), .B2(G20), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n858), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(G1956), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n863), .B1(new_n758), .B2(new_n761), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n856), .A2(new_n864), .ZN(G311));
  NAND2_X1  g440(.A1(G311), .A2(KEYINPUT95), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT95), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n867), .B1(new_n856), .B2(new_n864), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n866), .A2(new_n868), .ZN(G150));
  AND2_X1   g444(.A1(new_n524), .A2(G55), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n539), .A2(G93), .ZN(new_n871));
  NAND2_X1  g446(.A1(G80), .A2(G543), .ZN(new_n872));
  INV_X1    g447(.A(G67), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n872), .B1(new_n505), .B2(new_n873), .ZN(new_n874));
  AND2_X1   g449(.A1(new_n874), .A2(KEYINPUT97), .ZN(new_n875));
  OAI21_X1  g450(.A(G651), .B1(new_n874), .B2(KEYINPUT97), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n871), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n870), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(new_n628), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n553), .B1(new_n870), .B2(new_n877), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  XOR2_X1   g456(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n882));
  XNOR2_X1  g457(.A(new_n881), .B(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n617), .A2(G559), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n885), .B(KEYINPUT39), .Z(new_n886));
  AOI21_X1  g461(.A(G860), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n887), .B1(new_n886), .B2(new_n884), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n878), .A2(new_n625), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(KEYINPUT37), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n888), .A2(new_n890), .ZN(G145));
  INV_X1    g466(.A(KEYINPUT98), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n824), .B(new_n735), .ZN(new_n893));
  XOR2_X1   g468(.A(new_n893), .B(new_n641), .Z(new_n894));
  NAND3_X1  g469(.A1(new_n803), .A2(new_n809), .A3(new_n776), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n776), .B1(new_n803), .B2(new_n809), .ZN(new_n897));
  OAI21_X1  g472(.A(G162), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n810), .A2(new_n777), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n899), .A2(new_n490), .A3(new_n895), .ZN(new_n900));
  XOR2_X1   g475(.A(G160), .B(new_n637), .Z(new_n901));
  AND3_X1   g476(.A1(new_n898), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n901), .B1(new_n898), .B2(new_n900), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n894), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n898), .A2(new_n900), .ZN(new_n905));
  INV_X1    g480(.A(new_n901), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n898), .A2(new_n900), .A3(new_n901), .ZN(new_n908));
  INV_X1    g483(.A(new_n894), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n496), .B(KEYINPUT4), .ZN(new_n911));
  INV_X1    g486(.A(new_n495), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n485), .A2(G130), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n471), .A2(G142), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n472), .A2(G118), .ZN(new_n916));
  OAI21_X1  g491(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n917));
  OAI211_X1 g492(.A(new_n914), .B(new_n915), .C1(new_n916), .C2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n913), .B(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n904), .A2(new_n910), .A3(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(G37), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n919), .B1(new_n904), .B2(new_n910), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n892), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n904), .A2(new_n910), .ZN(new_n925));
  INV_X1    g500(.A(new_n919), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n927), .A2(KEYINPUT98), .A3(new_n921), .A4(new_n920), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n924), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n929), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g505(.A1(G290), .A2(new_n585), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n604), .A2(G288), .A3(new_n606), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(G305), .B(G303), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n931), .A2(new_n934), .A3(new_n932), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT42), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n939), .A2(KEYINPUT100), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(KEYINPUT100), .ZN(new_n941));
  XOR2_X1   g516(.A(new_n941), .B(KEYINPUT101), .Z(new_n942));
  OR3_X1    g517(.A1(new_n938), .A2(new_n940), .A3(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n942), .B1(new_n938), .B2(new_n940), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n624), .B1(new_n575), .B2(new_n577), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n576), .B1(new_n566), .B2(new_n573), .ZN(new_n947));
  AOI211_X1 g522(.A(KEYINPUT71), .B(new_n572), .C1(new_n562), .C2(new_n565), .ZN(new_n948));
  NOR3_X1   g523(.A1(new_n947), .A2(new_n948), .A3(new_n617), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT99), .B1(new_n946), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n617), .B1(new_n947), .B2(new_n948), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT99), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n950), .A2(new_n953), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n630), .B(new_n881), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n575), .A2(new_n624), .A3(new_n577), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(new_n951), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n958), .A2(KEYINPUT41), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n959), .B1(new_n954), .B2(KEYINPUT41), .ZN(new_n960));
  INV_X1    g535(.A(new_n955), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n945), .A2(new_n956), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n945), .B1(new_n962), .B2(new_n956), .ZN(new_n964));
  OAI21_X1  g539(.A(G868), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n965), .B1(G868), .B2(new_n878), .ZN(G295));
  OAI21_X1  g541(.A(new_n965), .B1(G868), .B2(new_n878), .ZN(G331));
  NAND2_X1  g542(.A1(G286), .A2(G301), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT102), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n525), .A2(new_n538), .A3(new_n536), .A4(new_n543), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n969), .B1(new_n968), .B2(new_n970), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n881), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n968), .A2(new_n970), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(KEYINPUT102), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n976), .A2(new_n880), .A3(new_n879), .A4(new_n971), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n978), .A2(new_n950), .A3(new_n953), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n979), .B1(new_n960), .B2(new_n978), .ZN(new_n980));
  AOI21_X1  g555(.A(G37), .B1(new_n980), .B2(new_n938), .ZN(new_n981));
  INV_X1    g556(.A(new_n953), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n952), .B1(new_n957), .B2(new_n951), .ZN(new_n983));
  OAI21_X1  g558(.A(KEYINPUT41), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n959), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n978), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  AND4_X1   g561(.A1(new_n950), .A2(new_n974), .A3(new_n953), .A4(new_n977), .ZN(new_n987));
  OR3_X1    g562(.A1(new_n986), .A2(new_n938), .A3(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT43), .B1(new_n981), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n938), .B1(new_n986), .B2(new_n987), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT41), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n991), .B1(new_n974), .B2(new_n977), .ZN(new_n992));
  OR2_X1    g567(.A1(new_n992), .A2(new_n954), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n938), .B1(new_n992), .B2(new_n958), .ZN(new_n994));
  AOI21_X1  g569(.A(G37), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  AND3_X1   g570(.A1(new_n990), .A2(new_n995), .A3(KEYINPUT43), .ZN(new_n996));
  OAI21_X1  g571(.A(KEYINPUT44), .B1(new_n989), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT44), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT43), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n999), .B1(new_n981), .B2(new_n988), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n990), .A2(new_n995), .A3(new_n999), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n998), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n997), .A2(new_n1002), .ZN(G397));
  INV_X1    g578(.A(G1384), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n913), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT45), .ZN(new_n1006));
  AND3_X1   g581(.A1(new_n479), .A2(G40), .A3(new_n483), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n824), .B(new_n829), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n776), .B(new_n712), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1008), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  OR2_X1    g586(.A1(new_n1011), .A2(KEYINPUT105), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(KEYINPUT105), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n735), .A2(new_n738), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1015), .B1(G2067), .B2(new_n824), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1008), .ZN(new_n1017));
  AND3_X1   g592(.A1(new_n1016), .A2(KEYINPUT124), .A3(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT124), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  OR3_X1    g595(.A1(G290), .A2(KEYINPUT103), .A3(G1986), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT103), .B1(G290), .B2(G1986), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1021), .A2(new_n1017), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT48), .ZN(new_n1024));
  OR2_X1    g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  AND2_X1   g600(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1026));
  XNOR2_X1  g601(.A(new_n735), .B(new_n738), .ZN(new_n1027));
  XNOR2_X1  g602(.A(new_n1027), .B(KEYINPUT106), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n1017), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1025), .A2(new_n1026), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(KEYINPUT46), .B1(new_n1017), .B2(new_n712), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1008), .B1(new_n1009), .B2(new_n777), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1017), .A2(KEYINPUT46), .A3(new_n712), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g611(.A(new_n1036), .B(KEYINPUT47), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1031), .A2(new_n1037), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1020), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT125), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(KEYINPUT125), .B1(new_n1020), .B2(new_n1038), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g618(.A(KEYINPUT108), .B(G8), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(G1384), .B1(new_n911), .B2(new_n912), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1045), .B1(new_n1007), .B2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n581), .A2(new_n584), .A3(G1976), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n1047), .A2(KEYINPUT109), .A3(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1007), .A2(new_n1046), .ZN(new_n1050));
  AOI21_X1  g625(.A(G1976), .B1(new_n581), .B2(new_n584), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1050), .A2(new_n1051), .A3(new_n1044), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT52), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1049), .A2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1047), .A2(KEYINPUT109), .A3(new_n1048), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1056), .A2(new_n1053), .A3(new_n1052), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  XOR2_X1   g633(.A(KEYINPUT110), .B(G1981), .Z(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n591), .A2(new_n593), .A3(new_n597), .A4(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(G1981), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1061), .B1(new_n742), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT49), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  OAI211_X1 g640(.A(KEYINPUT49), .B(new_n1061), .C1(new_n742), .C2(new_n1062), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1065), .A2(new_n1066), .A3(new_n1047), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1058), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT50), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n913), .A2(new_n1069), .A3(new_n1004), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(KEYINPUT112), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT112), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1046), .A2(new_n1072), .A3(new_n1069), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1007), .B1(new_n1046), .B2(new_n1069), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(KEYINPUT111), .ZN(new_n1076));
  INV_X1    g651(.A(G2090), .ZN(new_n1077));
  OAI21_X1  g652(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT111), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1078), .A2(new_n1079), .A3(new_n1007), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1074), .A2(new_n1076), .A3(new_n1077), .A4(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n913), .A2(KEYINPUT45), .A3(new_n1004), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1006), .B1(G164), .B2(G1384), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1082), .A2(new_n1083), .A3(new_n1007), .ZN(new_n1084));
  INV_X1    g659(.A(G1971), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1081), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(new_n1044), .ZN(new_n1088));
  NAND3_X1  g663(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT55), .ZN(new_n1090));
  INV_X1    g665(.A(G8), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1090), .B1(G166), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1089), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1088), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1084), .A2(new_n833), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1070), .A2(new_n1078), .A3(new_n782), .A4(new_n1007), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1045), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(G168), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1099), .A2(KEYINPUT63), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1095), .A2(new_n1100), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1070), .A2(new_n1078), .A3(new_n1077), .A4(new_n1007), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1086), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT107), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1093), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1089), .A2(KEYINPUT107), .A3(new_n1092), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1103), .A2(new_n1107), .A3(G8), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1068), .B1(new_n1101), .B2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g684(.A1(G288), .A2(G1976), .ZN(new_n1110));
  AND2_X1   g685(.A1(new_n1067), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1061), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1047), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1093), .B1(new_n1103), .B2(G8), .ZN(new_n1114));
  NOR3_X1   g689(.A1(new_n1068), .A2(new_n1099), .A3(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT63), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1113), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1109), .A2(new_n1117), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1058), .A2(new_n1108), .A3(new_n1067), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1119), .A2(new_n1095), .A3(KEYINPUT122), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT122), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1058), .A2(new_n1108), .A3(new_n1067), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1093), .B1(new_n1087), .B2(new_n1044), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1121), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1120), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT113), .ZN(new_n1126));
  NOR3_X1   g701(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1126), .B1(new_n1075), .B2(new_n1127), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1070), .A2(new_n1078), .A3(KEYINPUT113), .A4(new_n1007), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(new_n840), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT120), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT53), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n1084), .A2(new_n1133), .A3(G2078), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1131), .A2(new_n1132), .A3(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1133), .B1(new_n1084), .B2(G2078), .ZN(new_n1137));
  AOI21_X1  g712(.A(G1961), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1138));
  OAI21_X1  g713(.A(KEYINPUT120), .B1(new_n1138), .B2(new_n1134), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1136), .A2(new_n1137), .A3(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1125), .A2(G171), .A3(new_n1140), .ZN(new_n1141));
  NOR2_X1   g716(.A1(G168), .A2(new_n1045), .ZN(new_n1142));
  OR2_X1    g717(.A1(new_n1142), .A2(KEYINPUT51), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1143), .B1(new_n1098), .B2(KEYINPUT119), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(new_n1044), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT119), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1142), .ZN(new_n1149));
  AND2_X1   g724(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1149), .B1(new_n1150), .B2(new_n1091), .ZN(new_n1151));
  AOI22_X1  g726(.A1(new_n1144), .A2(new_n1148), .B1(new_n1151), .B2(KEYINPUT51), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1150), .A2(new_n1149), .ZN(new_n1153));
  OAI21_X1  g728(.A(KEYINPUT62), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1091), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1155));
  OAI21_X1  g730(.A(KEYINPUT51), .B1(new_n1155), .B2(new_n1142), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1142), .A2(KEYINPUT51), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1157), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1098), .A2(KEYINPUT119), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1156), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT62), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1153), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1154), .A2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1118), .B1(new_n1141), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1166));
  XOR2_X1   g741(.A(G301), .B(KEYINPUT54), .Z(new_n1167));
  AND2_X1   g742(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1168));
  INV_X1    g743(.A(G2078), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n479), .A2(KEYINPUT53), .A3(G40), .A4(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT121), .ZN(new_n1171));
  OR2_X1    g746(.A1(new_n482), .A2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n472), .B1(new_n482), .B2(new_n1171), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1170), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1168), .A2(new_n1174), .ZN(new_n1175));
  AND4_X1   g750(.A1(new_n1131), .A2(new_n1137), .A3(new_n1167), .A4(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1167), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1176), .B1(new_n1140), .B2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g753(.A(KEYINPUT122), .B1(new_n1119), .B2(new_n1095), .ZN(new_n1179));
  NOR3_X1   g754(.A1(new_n1122), .A2(new_n1123), .A3(new_n1121), .ZN(new_n1180));
  OAI211_X1 g755(.A(new_n1166), .B(new_n1178), .C1(new_n1179), .C2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT123), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND4_X1  g758(.A1(new_n1125), .A2(KEYINPUT123), .A3(new_n1166), .A4(new_n1178), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1050), .A2(G2067), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1186), .B1(new_n1130), .B2(new_n646), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1187), .A2(KEYINPUT60), .A3(new_n624), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT118), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1187), .A2(KEYINPUT60), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1191), .A2(new_n617), .ZN(new_n1192));
  NAND4_X1  g767(.A1(new_n1187), .A2(KEYINPUT118), .A3(KEYINPUT60), .A4(new_n624), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1190), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  OR2_X1    g769(.A1(new_n1187), .A2(KEYINPUT60), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1074), .A2(new_n1076), .A3(new_n1080), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1197), .A2(new_n862), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT57), .ZN(new_n1199));
  XNOR2_X1  g774(.A(new_n574), .B(new_n1199), .ZN(new_n1200));
  XNOR2_X1  g775(.A(KEYINPUT56), .B(G2072), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1168), .A2(new_n1007), .A3(new_n1201), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1198), .A2(new_n1200), .A3(new_n1202), .ZN(new_n1203));
  INV_X1    g778(.A(new_n1203), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1200), .B1(new_n1198), .B2(new_n1202), .ZN(new_n1205));
  OAI21_X1  g780(.A(KEYINPUT61), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1198), .A2(new_n1202), .ZN(new_n1207));
  INV_X1    g782(.A(new_n1200), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NOR2_X1   g784(.A1(KEYINPUT117), .A2(KEYINPUT61), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1209), .A2(new_n1203), .A3(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1205), .A2(KEYINPUT117), .ZN(new_n1212));
  NAND3_X1  g787(.A1(new_n1206), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  XOR2_X1   g788(.A(KEYINPUT58), .B(G1341), .Z(new_n1214));
  NAND2_X1  g789(.A1(new_n1050), .A2(new_n1214), .ZN(new_n1215));
  XNOR2_X1  g790(.A(new_n1215), .B(KEYINPUT116), .ZN(new_n1216));
  NOR2_X1   g791(.A1(new_n1084), .A2(G1996), .ZN(new_n1217));
  OAI21_X1  g792(.A(new_n553), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  XNOR2_X1  g793(.A(new_n1218), .B(KEYINPUT59), .ZN(new_n1219));
  NAND3_X1  g794(.A1(new_n1196), .A2(new_n1213), .A3(new_n1219), .ZN(new_n1220));
  INV_X1    g795(.A(KEYINPUT114), .ZN(new_n1221));
  OR3_X1    g796(.A1(new_n1187), .A2(new_n1221), .A3(new_n624), .ZN(new_n1222));
  OAI21_X1  g797(.A(new_n1221), .B1(new_n1187), .B2(new_n624), .ZN(new_n1223));
  NAND3_X1  g798(.A1(new_n1222), .A2(new_n1209), .A3(new_n1223), .ZN(new_n1224));
  NAND3_X1  g799(.A1(new_n1224), .A2(KEYINPUT115), .A3(new_n1203), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1224), .A2(new_n1203), .ZN(new_n1226));
  INV_X1    g801(.A(KEYINPUT115), .ZN(new_n1227));
  NAND2_X1  g802(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  NAND3_X1  g803(.A1(new_n1220), .A2(new_n1225), .A3(new_n1228), .ZN(new_n1229));
  AOI21_X1  g804(.A(new_n1165), .B1(new_n1185), .B2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g805(.A1(G290), .A2(G1986), .A3(new_n1017), .ZN(new_n1231));
  NAND2_X1  g806(.A1(new_n1023), .A2(new_n1231), .ZN(new_n1232));
  XNOR2_X1  g807(.A(new_n1232), .B(KEYINPUT104), .ZN(new_n1233));
  NAND3_X1  g808(.A1(new_n1233), .A2(new_n1026), .A3(new_n1029), .ZN(new_n1234));
  OAI21_X1  g809(.A(new_n1043), .B1(new_n1230), .B2(new_n1234), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g810(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1237));
  NOR2_X1   g811(.A1(G227), .A2(new_n464), .ZN(new_n1238));
  NAND2_X1  g812(.A1(new_n680), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g813(.A(KEYINPUT126), .ZN(new_n1240));
  NAND2_X1  g814(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  NAND3_X1  g815(.A1(new_n680), .A2(KEYINPUT126), .A3(new_n1238), .ZN(new_n1242));
  NAND2_X1  g816(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  NAND3_X1  g817(.A1(new_n1243), .A2(new_n724), .A3(new_n929), .ZN(new_n1244));
  NOR2_X1   g818(.A1(new_n1237), .A2(new_n1244), .ZN(G308));
  AND2_X1   g819(.A1(new_n929), .A2(new_n724), .ZN(new_n1246));
  OAI211_X1 g820(.A(new_n1246), .B(new_n1243), .C1(new_n1000), .C2(new_n1001), .ZN(G225));
endmodule


