

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591;

  XNOR2_X1 U323 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U324 ( .A(n346), .B(n345), .ZN(n348) );
  XOR2_X1 U325 ( .A(n343), .B(n342), .Z(n291) );
  XOR2_X1 U326 ( .A(n380), .B(n408), .Z(n292) );
  OR2_X1 U327 ( .A1(n554), .A2(n532), .ZN(n390) );
  XNOR2_X1 U328 ( .A(n344), .B(n291), .ZN(n345) );
  XNOR2_X1 U329 ( .A(n409), .B(G64GAT), .ZN(n410) );
  INV_X1 U330 ( .A(KEYINPUT37), .ZN(n416) );
  NOR2_X1 U331 ( .A1(n535), .A2(n472), .ZN(n576) );
  XNOR2_X1 U332 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U333 ( .A(n419), .B(n418), .ZN(n521) );
  NOR2_X1 U334 ( .A1(n476), .A2(n384), .ZN(n571) );
  XOR2_X1 U335 ( .A(n473), .B(KEYINPUT28), .Z(n538) );
  XNOR2_X1 U336 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U337 ( .A(n455), .B(G29GAT), .ZN(n456) );
  XNOR2_X1 U338 ( .A(n480), .B(n479), .ZN(G1351GAT) );
  XNOR2_X1 U339 ( .A(n457), .B(n456), .ZN(G1328GAT) );
  XOR2_X1 U340 ( .A(KEYINPUT0), .B(G134GAT), .Z(n294) );
  XNOR2_X1 U341 ( .A(KEYINPUT80), .B(G120GAT), .ZN(n293) );
  XNOR2_X1 U342 ( .A(n294), .B(n293), .ZN(n295) );
  XNOR2_X1 U343 ( .A(G113GAT), .B(n295), .ZN(n347) );
  XOR2_X1 U344 ( .A(KEYINPUT88), .B(KEYINPUT87), .Z(n297) );
  XNOR2_X1 U345 ( .A(KEYINPUT1), .B(KEYINPUT4), .ZN(n296) );
  XNOR2_X1 U346 ( .A(n297), .B(n296), .ZN(n311) );
  XOR2_X1 U347 ( .A(G155GAT), .B(G148GAT), .Z(n299) );
  XNOR2_X1 U348 ( .A(G29GAT), .B(G127GAT), .ZN(n298) );
  XNOR2_X1 U349 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U350 ( .A(KEYINPUT6), .B(KEYINPUT5), .Z(n301) );
  XNOR2_X1 U351 ( .A(G1GAT), .B(G57GAT), .ZN(n300) );
  XNOR2_X1 U352 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U353 ( .A(n303), .B(n302), .Z(n309) );
  XNOR2_X1 U354 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n304) );
  XNOR2_X1 U355 ( .A(n304), .B(KEYINPUT2), .ZN(n354) );
  XOR2_X1 U356 ( .A(G85GAT), .B(G162GAT), .Z(n306) );
  NAND2_X1 U357 ( .A1(G225GAT), .A2(G233GAT), .ZN(n305) );
  XNOR2_X1 U358 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U359 ( .A(n354), .B(n307), .ZN(n308) );
  XNOR2_X1 U360 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U361 ( .A(n311), .B(n310), .Z(n312) );
  XNOR2_X1 U362 ( .A(n347), .B(n312), .ZN(n535) );
  XOR2_X1 U363 ( .A(KEYINPUT9), .B(KEYINPUT74), .Z(n314) );
  XNOR2_X1 U364 ( .A(G106GAT), .B(KEYINPUT10), .ZN(n313) );
  XNOR2_X1 U365 ( .A(n314), .B(n313), .ZN(n331) );
  XOR2_X1 U366 ( .A(G92GAT), .B(KEYINPUT64), .Z(n316) );
  XNOR2_X1 U367 ( .A(KEYINPUT75), .B(KEYINPUT76), .ZN(n315) );
  XNOR2_X1 U368 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U369 ( .A(G36GAT), .B(G190GAT), .Z(n374) );
  XOR2_X1 U370 ( .A(n317), .B(n374), .Z(n319) );
  XNOR2_X1 U371 ( .A(G134GAT), .B(G218GAT), .ZN(n318) );
  XNOR2_X1 U372 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U373 ( .A(G99GAT), .B(G85GAT), .Z(n437) );
  XOR2_X1 U374 ( .A(n437), .B(KEYINPUT11), .Z(n321) );
  NAND2_X1 U375 ( .A1(G232GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U376 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U377 ( .A(n323), .B(n322), .Z(n329) );
  XOR2_X1 U378 ( .A(KEYINPUT67), .B(KEYINPUT8), .Z(n325) );
  XNOR2_X1 U379 ( .A(G43GAT), .B(G29GAT), .ZN(n324) );
  XNOR2_X1 U380 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U381 ( .A(KEYINPUT7), .B(n326), .ZN(n436) );
  INV_X1 U382 ( .A(n436), .ZN(n327) );
  XOR2_X1 U383 ( .A(G50GAT), .B(G162GAT), .Z(n349) );
  XNOR2_X1 U384 ( .A(n327), .B(n349), .ZN(n328) );
  XNOR2_X1 U385 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U386 ( .A(n331), .B(n330), .ZN(n563) );
  INV_X1 U387 ( .A(n563), .ZN(n548) );
  XNOR2_X1 U388 ( .A(n548), .B(KEYINPUT36), .ZN(n589) );
  INV_X1 U389 ( .A(KEYINPUT92), .ZN(n397) );
  INV_X1 U390 ( .A(KEYINPUT17), .ZN(n332) );
  NAND2_X1 U391 ( .A1(n332), .A2(KEYINPUT18), .ZN(n335) );
  INV_X1 U392 ( .A(KEYINPUT18), .ZN(n333) );
  NAND2_X1 U393 ( .A1(n333), .A2(KEYINPUT17), .ZN(n334) );
  NAND2_X1 U394 ( .A1(n335), .A2(n334), .ZN(n337) );
  XNOR2_X1 U395 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n336) );
  XNOR2_X1 U396 ( .A(n337), .B(n336), .ZN(n380) );
  XOR2_X1 U397 ( .A(G15GAT), .B(G127GAT), .Z(n408) );
  XNOR2_X1 U398 ( .A(G99GAT), .B(G190GAT), .ZN(n338) );
  XNOR2_X1 U399 ( .A(n292), .B(n338), .ZN(n346) );
  XOR2_X1 U400 ( .A(KEYINPUT20), .B(KEYINPUT81), .Z(n340) );
  XNOR2_X1 U401 ( .A(G43GAT), .B(G71GAT), .ZN(n339) );
  XNOR2_X1 U402 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U403 ( .A(n341), .B(KEYINPUT82), .ZN(n344) );
  XOR2_X1 U404 ( .A(G176GAT), .B(G183GAT), .Z(n343) );
  NAND2_X1 U405 ( .A1(G227GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U406 ( .A(n348), .B(n347), .ZN(n384) );
  INV_X1 U407 ( .A(n384), .ZN(n391) );
  XOR2_X1 U408 ( .A(KEYINPUT83), .B(KEYINPUT23), .Z(n351) );
  XOR2_X1 U409 ( .A(G22GAT), .B(G155GAT), .Z(n400) );
  XNOR2_X1 U410 ( .A(n349), .B(n400), .ZN(n350) );
  XNOR2_X1 U411 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U412 ( .A(n352), .B(G204GAT), .Z(n359) );
  INV_X1 U413 ( .A(KEYINPUT84), .ZN(n353) );
  XNOR2_X1 U414 ( .A(n354), .B(n353), .ZN(n356) );
  NAND2_X1 U415 ( .A1(G228GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U416 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U417 ( .A(n357), .B(KEYINPUT85), .ZN(n358) );
  XNOR2_X1 U418 ( .A(n359), .B(n358), .ZN(n363) );
  XOR2_X1 U419 ( .A(KEYINPUT22), .B(G211GAT), .Z(n361) );
  XNOR2_X1 U420 ( .A(KEYINPUT86), .B(KEYINPUT24), .ZN(n360) );
  XNOR2_X1 U421 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U422 ( .A(n363), .B(n362), .ZN(n368) );
  XOR2_X1 U423 ( .A(G78GAT), .B(G148GAT), .Z(n365) );
  XNOR2_X1 U424 ( .A(G106GAT), .B(KEYINPUT71), .ZN(n364) );
  XNOR2_X1 U425 ( .A(n365), .B(n364), .ZN(n448) );
  XNOR2_X1 U426 ( .A(G197GAT), .B(G218GAT), .ZN(n366) );
  XNOR2_X1 U427 ( .A(n366), .B(KEYINPUT21), .ZN(n371) );
  XOR2_X1 U428 ( .A(n448), .B(n371), .Z(n367) );
  XNOR2_X1 U429 ( .A(n368), .B(n367), .ZN(n473) );
  NOR2_X1 U430 ( .A1(n391), .A2(n473), .ZN(n369) );
  XNOR2_X1 U431 ( .A(n369), .B(KEYINPUT26), .ZN(n575) );
  INV_X1 U432 ( .A(n575), .ZN(n554) );
  XNOR2_X1 U433 ( .A(G8GAT), .B(G183GAT), .ZN(n370) );
  XNOR2_X1 U434 ( .A(n370), .B(G211GAT), .ZN(n401) );
  XOR2_X1 U435 ( .A(n371), .B(KEYINPUT89), .Z(n373) );
  NAND2_X1 U436 ( .A1(G226GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U437 ( .A(n373), .B(n372), .ZN(n377) );
  XNOR2_X1 U438 ( .A(n374), .B(KEYINPUT90), .ZN(n375) );
  XNOR2_X1 U439 ( .A(n375), .B(KEYINPUT91), .ZN(n376) );
  XOR2_X1 U440 ( .A(n377), .B(n376), .Z(n382) );
  XOR2_X1 U441 ( .A(G64GAT), .B(G92GAT), .Z(n379) );
  XNOR2_X1 U442 ( .A(G176GAT), .B(G204GAT), .ZN(n378) );
  XNOR2_X1 U443 ( .A(n379), .B(n378), .ZN(n447) );
  XNOR2_X1 U444 ( .A(n380), .B(n447), .ZN(n381) );
  XNOR2_X1 U445 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U446 ( .A(n401), .B(n383), .ZN(n493) );
  XNOR2_X1 U447 ( .A(KEYINPUT27), .B(n493), .ZN(n532) );
  INV_X1 U448 ( .A(n473), .ZN(n386) );
  NOR2_X1 U449 ( .A1(n384), .A2(n493), .ZN(n385) );
  NOR2_X1 U450 ( .A1(n386), .A2(n385), .ZN(n387) );
  XOR2_X1 U451 ( .A(KEYINPUT25), .B(n387), .Z(n388) );
  NOR2_X1 U452 ( .A1(n535), .A2(n388), .ZN(n389) );
  NAND2_X1 U453 ( .A1(n390), .A2(n389), .ZN(n395) );
  NOR2_X1 U454 ( .A1(n532), .A2(n538), .ZN(n392) );
  NAND2_X1 U455 ( .A1(n384), .A2(n392), .ZN(n393) );
  NAND2_X1 U456 ( .A1(n393), .A2(n535), .ZN(n394) );
  NAND2_X1 U457 ( .A1(n395), .A2(n394), .ZN(n396) );
  XNOR2_X1 U458 ( .A(n397), .B(n396), .ZN(n486) );
  XOR2_X1 U459 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n399) );
  XNOR2_X1 U460 ( .A(G1GAT), .B(KEYINPUT14), .ZN(n398) );
  XNOR2_X1 U461 ( .A(n399), .B(n398), .ZN(n413) );
  XNOR2_X1 U462 ( .A(n401), .B(n400), .ZN(n403) );
  AND2_X1 U463 ( .A1(G231GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U464 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U465 ( .A(n404), .B(KEYINPUT77), .Z(n407) );
  XNOR2_X1 U466 ( .A(G71GAT), .B(G57GAT), .ZN(n405) );
  XNOR2_X1 U467 ( .A(n405), .B(KEYINPUT13), .ZN(n438) );
  XNOR2_X1 U468 ( .A(n438), .B(KEYINPUT78), .ZN(n406) );
  XNOR2_X1 U469 ( .A(n407), .B(n406), .ZN(n411) );
  XOR2_X1 U470 ( .A(n408), .B(G78GAT), .Z(n409) );
  XOR2_X1 U471 ( .A(n413), .B(n412), .Z(n585) );
  NAND2_X1 U472 ( .A1(n486), .A2(n585), .ZN(n414) );
  XNOR2_X1 U473 ( .A(n414), .B(KEYINPUT96), .ZN(n415) );
  NOR2_X1 U474 ( .A1(n589), .A2(n415), .ZN(n419) );
  XNOR2_X1 U475 ( .A(KEYINPUT97), .B(KEYINPUT98), .ZN(n417) );
  XOR2_X1 U476 ( .A(G8GAT), .B(KEYINPUT68), .Z(n421) );
  XNOR2_X1 U477 ( .A(KEYINPUT29), .B(KEYINPUT65), .ZN(n420) );
  XNOR2_X1 U478 ( .A(n421), .B(n420), .ZN(n434) );
  XOR2_X1 U479 ( .A(G22GAT), .B(G141GAT), .Z(n423) );
  XNOR2_X1 U480 ( .A(G50GAT), .B(G36GAT), .ZN(n422) );
  XNOR2_X1 U481 ( .A(n423), .B(n422), .ZN(n427) );
  XOR2_X1 U482 ( .A(G113GAT), .B(G15GAT), .Z(n425) );
  XNOR2_X1 U483 ( .A(G169GAT), .B(G197GAT), .ZN(n424) );
  XNOR2_X1 U484 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U485 ( .A(n427), .B(n426), .Z(n432) );
  XOR2_X1 U486 ( .A(KEYINPUT66), .B(G1GAT), .Z(n429) );
  NAND2_X1 U487 ( .A1(G229GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U488 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U489 ( .A(KEYINPUT30), .B(n430), .ZN(n431) );
  XNOR2_X1 U490 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U491 ( .A(n434), .B(n433), .Z(n435) );
  XOR2_X1 U492 ( .A(n436), .B(n435), .Z(n577) );
  INV_X1 U493 ( .A(n577), .ZN(n568) );
  XOR2_X1 U494 ( .A(n438), .B(n437), .Z(n440) );
  NAND2_X1 U495 ( .A1(G230GAT), .A2(G233GAT), .ZN(n439) );
  XNOR2_X1 U496 ( .A(n440), .B(n439), .ZN(n452) );
  XOR2_X1 U497 ( .A(KEYINPUT73), .B(KEYINPUT70), .Z(n442) );
  XNOR2_X1 U498 ( .A(KEYINPUT69), .B(KEYINPUT33), .ZN(n441) );
  XNOR2_X1 U499 ( .A(n442), .B(n441), .ZN(n446) );
  XOR2_X1 U500 ( .A(KEYINPUT72), .B(KEYINPUT31), .Z(n444) );
  XNOR2_X1 U501 ( .A(G120GAT), .B(KEYINPUT32), .ZN(n443) );
  XNOR2_X1 U502 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U503 ( .A(n446), .B(n445), .Z(n450) );
  XNOR2_X1 U504 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U505 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U506 ( .A(n452), .B(n451), .Z(n581) );
  NAND2_X1 U507 ( .A1(n568), .A2(n581), .ZN(n488) );
  OR2_X1 U508 ( .A1(n521), .A2(n488), .ZN(n453) );
  XNOR2_X1 U509 ( .A(n453), .B(KEYINPUT38), .ZN(n454) );
  XNOR2_X1 U510 ( .A(KEYINPUT99), .B(n454), .ZN(n504) );
  NAND2_X1 U511 ( .A1(n535), .A2(n504), .ZN(n457) );
  XOR2_X1 U512 ( .A(KEYINPUT100), .B(KEYINPUT39), .Z(n455) );
  XOR2_X1 U513 ( .A(KEYINPUT122), .B(KEYINPUT55), .Z(n475) );
  XOR2_X1 U514 ( .A(KEYINPUT54), .B(KEYINPUT121), .Z(n471) );
  XNOR2_X1 U515 ( .A(n585), .B(KEYINPUT110), .ZN(n573) );
  XNOR2_X1 U516 ( .A(KEYINPUT41), .B(n581), .ZN(n557) );
  INV_X1 U517 ( .A(n557), .ZN(n507) );
  NOR2_X1 U518 ( .A1(n507), .A2(n577), .ZN(n459) );
  XNOR2_X1 U519 ( .A(KEYINPUT46), .B(KEYINPUT111), .ZN(n458) );
  XNOR2_X1 U520 ( .A(n459), .B(n458), .ZN(n460) );
  NAND2_X1 U521 ( .A1(n573), .A2(n460), .ZN(n461) );
  NOR2_X1 U522 ( .A1(n563), .A2(n461), .ZN(n462) );
  XOR2_X1 U523 ( .A(KEYINPUT47), .B(n462), .Z(n468) );
  NOR2_X1 U524 ( .A1(n585), .A2(n589), .ZN(n463) );
  XNOR2_X1 U525 ( .A(KEYINPUT45), .B(n463), .ZN(n464) );
  NAND2_X1 U526 ( .A1(n464), .A2(n581), .ZN(n465) );
  NOR2_X1 U527 ( .A1(n568), .A2(n465), .ZN(n466) );
  XNOR2_X1 U528 ( .A(KEYINPUT112), .B(n466), .ZN(n467) );
  NOR2_X1 U529 ( .A1(n468), .A2(n467), .ZN(n469) );
  XNOR2_X1 U530 ( .A(n469), .B(KEYINPUT48), .ZN(n533) );
  NOR2_X1 U531 ( .A1(n533), .A2(n493), .ZN(n470) );
  XOR2_X1 U532 ( .A(n471), .B(n470), .Z(n472) );
  NAND2_X1 U533 ( .A1(n576), .A2(n473), .ZN(n474) );
  XNOR2_X1 U534 ( .A(n475), .B(n474), .ZN(n476) );
  NAND2_X1 U535 ( .A1(n571), .A2(n563), .ZN(n480) );
  XOR2_X1 U536 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n478) );
  INV_X1 U537 ( .A(G190GAT), .ZN(n477) );
  NAND2_X1 U538 ( .A1(n571), .A2(n557), .ZN(n483) );
  XOR2_X1 U539 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n481) );
  XNOR2_X1 U540 ( .A(n481), .B(G176GAT), .ZN(n482) );
  XNOR2_X1 U541 ( .A(n483), .B(n482), .ZN(G1349GAT) );
  INV_X1 U542 ( .A(n585), .ZN(n561) );
  NAND2_X1 U543 ( .A1(n561), .A2(n548), .ZN(n484) );
  XNOR2_X1 U544 ( .A(n484), .B(KEYINPUT16), .ZN(n485) );
  XNOR2_X1 U545 ( .A(n485), .B(KEYINPUT79), .ZN(n487) );
  NAND2_X1 U546 ( .A1(n487), .A2(n486), .ZN(n509) );
  NOR2_X1 U547 ( .A1(n488), .A2(n509), .ZN(n498) );
  NAND2_X1 U548 ( .A1(n498), .A2(n535), .ZN(n492) );
  XOR2_X1 U549 ( .A(KEYINPUT93), .B(KEYINPUT34), .Z(n490) );
  XNOR2_X1 U550 ( .A(G1GAT), .B(KEYINPUT94), .ZN(n489) );
  XNOR2_X1 U551 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n492), .B(n491), .ZN(G1324GAT) );
  INV_X1 U553 ( .A(n493), .ZN(n523) );
  NAND2_X1 U554 ( .A1(n498), .A2(n523), .ZN(n494) );
  XNOR2_X1 U555 ( .A(n494), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U556 ( .A(KEYINPUT95), .B(KEYINPUT35), .Z(n496) );
  NAND2_X1 U557 ( .A1(n498), .A2(n391), .ZN(n495) );
  XNOR2_X1 U558 ( .A(n496), .B(n495), .ZN(n497) );
  XOR2_X1 U559 ( .A(G15GAT), .B(n497), .Z(G1326GAT) );
  NAND2_X1 U560 ( .A1(n498), .A2(n538), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n499), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U562 ( .A(G36GAT), .B(KEYINPUT101), .Z(n501) );
  NAND2_X1 U563 ( .A1(n523), .A2(n504), .ZN(n500) );
  XNOR2_X1 U564 ( .A(n501), .B(n500), .ZN(G1329GAT) );
  NAND2_X1 U565 ( .A1(n504), .A2(n391), .ZN(n502) );
  XNOR2_X1 U566 ( .A(n502), .B(KEYINPUT40), .ZN(n503) );
  XNOR2_X1 U567 ( .A(G43GAT), .B(n503), .ZN(G1330GAT) );
  NAND2_X1 U568 ( .A1(n504), .A2(n538), .ZN(n505) );
  XNOR2_X1 U569 ( .A(n505), .B(KEYINPUT102), .ZN(n506) );
  XNOR2_X1 U570 ( .A(G50GAT), .B(n506), .ZN(G1331GAT) );
  XOR2_X1 U571 ( .A(KEYINPUT103), .B(KEYINPUT42), .Z(n511) );
  NOR2_X1 U572 ( .A1(n507), .A2(n568), .ZN(n508) );
  XOR2_X1 U573 ( .A(n508), .B(KEYINPUT104), .Z(n520) );
  NOR2_X1 U574 ( .A1(n520), .A2(n509), .ZN(n517) );
  NAND2_X1 U575 ( .A1(n517), .A2(n535), .ZN(n510) );
  XNOR2_X1 U576 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U577 ( .A(G57GAT), .B(n512), .ZN(G1332GAT) );
  XOR2_X1 U578 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n514) );
  NAND2_X1 U579 ( .A1(n517), .A2(n523), .ZN(n513) );
  XNOR2_X1 U580 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U581 ( .A(G64GAT), .B(n515), .ZN(G1333GAT) );
  NAND2_X1 U582 ( .A1(n391), .A2(n517), .ZN(n516) );
  XNOR2_X1 U583 ( .A(n516), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U584 ( .A(G78GAT), .B(KEYINPUT43), .Z(n519) );
  NAND2_X1 U585 ( .A1(n517), .A2(n538), .ZN(n518) );
  XNOR2_X1 U586 ( .A(n519), .B(n518), .ZN(G1335GAT) );
  NOR2_X1 U587 ( .A1(n521), .A2(n520), .ZN(n528) );
  NAND2_X1 U588 ( .A1(n528), .A2(n535), .ZN(n522) );
  XNOR2_X1 U589 ( .A(n522), .B(G85GAT), .ZN(G1336GAT) );
  XOR2_X1 U590 ( .A(G92GAT), .B(KEYINPUT107), .Z(n525) );
  NAND2_X1 U591 ( .A1(n528), .A2(n523), .ZN(n524) );
  XNOR2_X1 U592 ( .A(n525), .B(n524), .ZN(G1337GAT) );
  NAND2_X1 U593 ( .A1(n391), .A2(n528), .ZN(n526) );
  XNOR2_X1 U594 ( .A(n526), .B(KEYINPUT108), .ZN(n527) );
  XNOR2_X1 U595 ( .A(G99GAT), .B(n527), .ZN(G1338GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT44), .B(KEYINPUT109), .Z(n530) );
  NAND2_X1 U597 ( .A1(n528), .A2(n538), .ZN(n529) );
  XNOR2_X1 U598 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U599 ( .A(G106GAT), .B(n531), .ZN(G1339GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n540) );
  NOR2_X1 U601 ( .A1(n533), .A2(n532), .ZN(n534) );
  NAND2_X1 U602 ( .A1(n535), .A2(n534), .ZN(n555) );
  NOR2_X1 U603 ( .A1(n384), .A2(n555), .ZN(n536) );
  XNOR2_X1 U604 ( .A(n536), .B(KEYINPUT113), .ZN(n537) );
  NOR2_X1 U605 ( .A1(n538), .A2(n537), .ZN(n545) );
  NAND2_X1 U606 ( .A1(n545), .A2(n568), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U608 ( .A(G113GAT), .B(n541), .ZN(G1340GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n543) );
  NAND2_X1 U610 ( .A1(n545), .A2(n557), .ZN(n542) );
  XNOR2_X1 U611 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U612 ( .A(G120GAT), .B(n544), .ZN(G1341GAT) );
  INV_X1 U613 ( .A(n545), .ZN(n549) );
  NOR2_X1 U614 ( .A1(n573), .A2(n549), .ZN(n546) );
  XOR2_X1 U615 ( .A(KEYINPUT50), .B(n546), .Z(n547) );
  XNOR2_X1 U616 ( .A(G127GAT), .B(n547), .ZN(G1342GAT) );
  NOR2_X1 U617 ( .A1(n549), .A2(n548), .ZN(n553) );
  XOR2_X1 U618 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n551) );
  XNOR2_X1 U619 ( .A(G134GAT), .B(KEYINPUT118), .ZN(n550) );
  XNOR2_X1 U620 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U621 ( .A(n553), .B(n552), .ZN(G1343GAT) );
  NOR2_X1 U622 ( .A1(n554), .A2(n555), .ZN(n564) );
  NAND2_X1 U623 ( .A1(n568), .A2(n564), .ZN(n556) );
  XNOR2_X1 U624 ( .A(G141GAT), .B(n556), .ZN(G1344GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n559) );
  NAND2_X1 U626 ( .A1(n564), .A2(n557), .ZN(n558) );
  XNOR2_X1 U627 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U628 ( .A(G148GAT), .B(n560), .ZN(G1345GAT) );
  NAND2_X1 U629 ( .A1(n564), .A2(n561), .ZN(n562) );
  XNOR2_X1 U630 ( .A(G155GAT), .B(n562), .ZN(G1346GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n566) );
  NAND2_X1 U632 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U634 ( .A(G162GAT), .B(n567), .ZN(G1347GAT) );
  XOR2_X1 U635 ( .A(G169GAT), .B(KEYINPUT123), .Z(n570) );
  NAND2_X1 U636 ( .A1(n571), .A2(n568), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n570), .B(n569), .ZN(G1348GAT) );
  INV_X1 U638 ( .A(n571), .ZN(n572) );
  NOR2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U640 ( .A(G183GAT), .B(n574), .Z(G1350GAT) );
  NAND2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n588) );
  NOR2_X1 U642 ( .A1(n577), .A2(n588), .ZN(n579) );
  XNOR2_X1 U643 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(G197GAT), .B(n580), .ZN(G1352GAT) );
  NOR2_X1 U646 ( .A1(n581), .A2(n588), .ZN(n583) );
  XNOR2_X1 U647 ( .A(KEYINPUT125), .B(KEYINPUT61), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(n584) );
  XOR2_X1 U649 ( .A(G204GAT), .B(n584), .Z(G1353GAT) );
  NOR2_X1 U650 ( .A1(n585), .A2(n588), .ZN(n586) );
  XOR2_X1 U651 ( .A(KEYINPUT126), .B(n586), .Z(n587) );
  XNOR2_X1 U652 ( .A(G211GAT), .B(n587), .ZN(G1354GAT) );
  NOR2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U654 ( .A(KEYINPUT62), .B(n590), .Z(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

