//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 0 0 0 1 1 0 1 1 0 0 0 0 1 0 1 0 1 0 0 1 1 0 0 0 0 0 0 0 0 1 1 1 0 0 1 0 0 0 0 1 1 0 0 0 1 0 1 1 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:43 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  OR3_X1    g0003(.A1(new_n203), .A2(KEYINPUT64), .A3(G13), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(new_n203), .B2(G13), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT0), .Z(new_n208));
  INV_X1    g0008(.A(G87), .ZN(new_n209));
  INV_X1    g0009(.A(G250), .ZN(new_n210));
  INV_X1    g0010(.A(G97), .ZN(new_n211));
  INV_X1    g0011(.A(G257), .ZN(new_n212));
  OAI22_X1  g0012(.A1(new_n209), .A2(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AOI21_X1  g0013(.A(new_n213), .B1(G68), .B2(G238), .ZN(new_n214));
  INV_X1    g0014(.A(G107), .ZN(new_n215));
  INV_X1    g0015(.A(G264), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  AOI21_X1  g0017(.A(new_n217), .B1(G116), .B2(G270), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G50), .A2(G226), .ZN(new_n219));
  INV_X1    g0019(.A(G77), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n218), .B(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G58), .ZN(new_n223));
  INV_X1    g0023(.A(G232), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n203), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT1), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g0030(.A(G68), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n223), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(G50), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT65), .ZN(new_n234));
  AOI211_X1 g0034(.A(new_n208), .B(new_n227), .C1(new_n230), .C2(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(new_n224), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G264), .ZN(new_n241));
  INV_X1    g0041(.A(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n239), .B(new_n243), .Z(G358));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G97), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  XNOR2_X1  g0051(.A(KEYINPUT8), .B(G58), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G1), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n254), .A2(G13), .A3(G20), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(new_n228), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n254), .A2(G20), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n257), .B1(new_n262), .B2(new_n253), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT3), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT72), .ZN(new_n265));
  INV_X1    g0065(.A(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(KEYINPUT72), .A2(G33), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n264), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n264), .A2(G33), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G1698), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n272), .B1(G226), .B2(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(G223), .A2(G1698), .ZN(new_n275));
  OAI22_X1  g0075(.A1(new_n274), .A2(new_n275), .B1(new_n266), .B2(new_n209), .ZN(new_n276));
  INV_X1    g0076(.A(G41), .ZN(new_n277));
  OAI211_X1 g0077(.A(G1), .B(G13), .C1(new_n266), .C2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT75), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n254), .B1(G41), .B2(G45), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n278), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n281), .B1(new_n283), .B2(new_n224), .ZN(new_n284));
  INV_X1    g0084(.A(G274), .ZN(new_n285));
  OR2_X1    g0085(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  NAND4_X1  g0086(.A1(new_n278), .A2(KEYINPUT75), .A3(G232), .A4(new_n282), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n284), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(KEYINPUT76), .ZN(new_n289));
  OR2_X1    g0089(.A1(new_n288), .A2(KEYINPUT76), .ZN(new_n290));
  AND4_X1   g0090(.A1(G190), .A2(new_n280), .A3(new_n289), .A4(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n232), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n223), .A2(new_n231), .ZN(new_n293));
  OR2_X1    g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(G20), .A2(G33), .ZN(new_n295));
  AOI22_X1  g0095(.A1(new_n294), .A2(G20), .B1(G159), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(KEYINPUT73), .B1(new_n269), .B2(new_n271), .ZN(new_n297));
  AND2_X1   g0097(.A1(KEYINPUT72), .A2(G33), .ZN(new_n298));
  NOR2_X1   g0098(.A1(KEYINPUT72), .A2(G33), .ZN(new_n299));
  OAI21_X1  g0099(.A(KEYINPUT3), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT73), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n300), .A2(new_n301), .A3(new_n270), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n297), .A2(new_n229), .A3(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT74), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT7), .ZN(new_n305));
  AND3_X1   g0105(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n304), .B1(new_n303), .B2(new_n305), .ZN(new_n307));
  NOR3_X1   g0107(.A1(new_n272), .A2(new_n305), .A3(G20), .ZN(new_n308));
  NOR3_X1   g0108(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  OAI211_X1 g0109(.A(KEYINPUT16), .B(new_n296), .C1(new_n309), .C2(new_n231), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n266), .A2(KEYINPUT3), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n267), .A2(new_n268), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n311), .B1(new_n312), .B2(KEYINPUT3), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n313), .A2(KEYINPUT7), .A3(new_n229), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n270), .A2(new_n311), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n305), .B1(new_n316), .B2(G20), .ZN(new_n317));
  AND2_X1   g0117(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n296), .B1(new_n318), .B2(new_n231), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT16), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n260), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  AOI211_X1 g0121(.A(new_n263), .B(new_n291), .C1(new_n310), .C2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT17), .ZN(new_n323));
  OR2_X1    g0123(.A1(new_n323), .A2(KEYINPUT78), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n280), .A2(new_n289), .A3(new_n290), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(G200), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n323), .A2(KEYINPUT78), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n322), .A2(new_n324), .A3(new_n326), .A4(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n310), .A2(new_n321), .ZN(new_n329));
  INV_X1    g0129(.A(new_n291), .ZN(new_n330));
  INV_X1    g0130(.A(new_n263), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n329), .A2(new_n326), .A3(new_n330), .A4(new_n331), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n332), .A2(KEYINPUT78), .A3(new_n323), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n328), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT77), .ZN(new_n335));
  INV_X1    g0135(.A(new_n296), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n303), .A2(new_n305), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(KEYINPUT74), .ZN(new_n338));
  INV_X1    g0138(.A(new_n308), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  AOI211_X1 g0141(.A(new_n320), .B(new_n336), .C1(new_n341), .C2(G68), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n319), .A2(new_n320), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(new_n259), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n331), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n325), .A2(G169), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n280), .A2(new_n290), .A3(G179), .A4(new_n289), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(KEYINPUT18), .B1(new_n345), .B2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n263), .B1(new_n310), .B2(new_n321), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT18), .ZN(new_n351));
  AND2_X1   g0151(.A1(new_n346), .A2(new_n347), .ZN(new_n352));
  NOR3_X1   g0152(.A1(new_n350), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n335), .B1(new_n349), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n351), .B1(new_n350), .B2(new_n352), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n336), .B1(new_n341), .B2(G68), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n344), .B1(new_n356), .B2(KEYINPUT16), .ZN(new_n357));
  OAI211_X1 g0157(.A(KEYINPUT18), .B(new_n348), .C1(new_n357), .C2(new_n263), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n355), .A2(new_n358), .A3(KEYINPUT77), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n334), .B1(new_n354), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n273), .A2(G222), .ZN(new_n361));
  NAND2_X1  g0161(.A1(G223), .A2(G1698), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n316), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n363), .B(new_n279), .C1(G77), .C2(new_n316), .ZN(new_n364));
  INV_X1    g0164(.A(G226), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n364), .B(new_n286), .C1(new_n365), .C2(new_n283), .ZN(new_n366));
  OR2_X1    g0166(.A1(new_n366), .A2(G179), .ZN(new_n367));
  OAI21_X1  g0167(.A(G20), .B1(new_n232), .B2(G50), .ZN(new_n368));
  INV_X1    g0168(.A(G150), .ZN(new_n369));
  INV_X1    g0169(.A(new_n295), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n229), .A2(G33), .ZN(new_n371));
  OAI221_X1 g0171(.A(new_n368), .B1(new_n369), .B2(new_n370), .C1(new_n371), .C2(new_n252), .ZN(new_n372));
  INV_X1    g0172(.A(G50), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n372), .A2(new_n259), .B1(new_n373), .B2(new_n256), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n374), .B1(new_n373), .B2(new_n262), .ZN(new_n375));
  INV_X1    g0175(.A(G169), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n366), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n367), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n253), .A2(new_n295), .B1(G20), .B2(G77), .ZN(new_n380));
  XNOR2_X1  g0180(.A(KEYINPUT15), .B(G87), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n380), .B1(new_n371), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n259), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n383), .B1(G77), .B2(new_n255), .ZN(new_n384));
  INV_X1    g0184(.A(new_n262), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n384), .B1(G77), .B2(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n279), .B1(new_n316), .B2(G107), .ZN(new_n387));
  NAND2_X1  g0187(.A1(G238), .A2(G1698), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(new_n224), .B2(G1698), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n315), .A2(new_n389), .ZN(new_n390));
  OAI221_X1 g0190(.A(new_n286), .B1(new_n283), .B2(new_n221), .C1(new_n387), .C2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(G190), .ZN(new_n392));
  OR2_X1    g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  XNOR2_X1  g0193(.A(KEYINPUT66), .B(G200), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n386), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n366), .A2(new_n394), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n366), .A2(new_n392), .ZN(new_n399));
  XNOR2_X1  g0199(.A(new_n375), .B(KEYINPUT68), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n399), .B1(new_n400), .B2(KEYINPUT9), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT69), .ZN(new_n402));
  NOR3_X1   g0202(.A1(new_n400), .A2(new_n402), .A3(KEYINPUT9), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT68), .ZN(new_n404));
  XNOR2_X1  g0204(.A(new_n375), .B(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT9), .ZN(new_n406));
  AOI21_X1  g0206(.A(KEYINPUT69), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n398), .B(new_n401), .C1(new_n403), .C2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(KEYINPUT10), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n402), .B1(new_n400), .B2(KEYINPUT9), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n405), .A2(KEYINPUT69), .A3(new_n406), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT10), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n412), .A2(new_n413), .A3(new_n398), .A4(new_n401), .ZN(new_n414));
  AOI211_X1 g0214(.A(new_n379), .B(new_n397), .C1(new_n409), .C2(new_n414), .ZN(new_n415));
  OAI22_X1  g0215(.A1(new_n370), .A2(new_n373), .B1(new_n229), .B2(G68), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n371), .A2(new_n220), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n259), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  XNOR2_X1  g0218(.A(new_n418), .B(KEYINPUT11), .ZN(new_n419));
  OAI21_X1  g0219(.A(KEYINPUT12), .B1(new_n255), .B2(G68), .ZN(new_n420));
  OR3_X1    g0220(.A1(new_n255), .A2(KEYINPUT12), .A3(G68), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n385), .A2(G68), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT14), .ZN(new_n425));
  INV_X1    g0225(.A(G238), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n286), .B1(new_n283), .B2(new_n426), .ZN(new_n427));
  XNOR2_X1  g0227(.A(new_n427), .B(KEYINPUT70), .ZN(new_n428));
  NAND2_X1  g0228(.A1(G33), .A2(G97), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n224), .A2(G1698), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n430), .B1(G226), .B2(G1698), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n429), .B1(new_n431), .B2(new_n315), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n279), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n428), .A2(new_n433), .ZN(new_n434));
  OR2_X1    g0234(.A1(new_n434), .A2(KEYINPUT13), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(KEYINPUT13), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n425), .B1(new_n437), .B2(G169), .ZN(new_n438));
  AOI211_X1 g0238(.A(KEYINPUT14), .B(new_n376), .C1(new_n435), .C2(new_n436), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n437), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(G179), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n424), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT71), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n437), .A2(G200), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n424), .B1(new_n437), .B2(new_n392), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n444), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n447), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n449), .A2(KEYINPUT71), .A3(new_n445), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n443), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  OR2_X1    g0251(.A1(new_n391), .A2(G179), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT67), .ZN(new_n453));
  OR2_X1    g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n452), .A2(new_n453), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n386), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n391), .A2(new_n376), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n360), .A2(new_n415), .A3(new_n451), .A4(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n215), .B1(new_n314), .B2(new_n317), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT6), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n211), .A2(new_n215), .ZN(new_n463));
  NOR2_X1   g0263(.A1(G97), .A2(G107), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n215), .A2(KEYINPUT6), .A3(G97), .ZN(new_n466));
  AND2_X1   g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI22_X1  g0267(.A1(new_n467), .A2(new_n229), .B1(new_n220), .B2(new_n370), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n259), .B1(new_n461), .B2(new_n468), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n260), .B(new_n255), .C1(G1), .C2(new_n266), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(G97), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n469), .B(new_n472), .C1(G97), .C2(new_n255), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT4), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n300), .A2(new_n270), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n221), .A2(G1698), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n474), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n316), .A2(G250), .A3(G1698), .ZN(new_n479));
  NAND2_X1  g0279(.A1(G33), .A2(G283), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n476), .A2(new_n270), .A3(new_n311), .A4(KEYINPUT4), .ZN(new_n482));
  XOR2_X1   g0282(.A(new_n482), .B(KEYINPUT79), .Z(new_n483));
  OAI21_X1  g0283(.A(new_n279), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(G45), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n485), .A2(G1), .ZN(new_n486));
  AND2_X1   g0286(.A1(KEYINPUT5), .A2(G41), .ZN(new_n487));
  NOR2_X1   g0287(.A1(KEYINPUT5), .A2(G41), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n489), .A2(G257), .A3(new_n278), .ZN(new_n490));
  OR2_X1    g0290(.A1(new_n489), .A2(new_n285), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n484), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n473), .B1(new_n493), .B2(G190), .ZN(new_n494));
  INV_X1    g0294(.A(G200), .ZN(new_n495));
  OAI21_X1  g0295(.A(KEYINPUT80), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT80), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n492), .A2(new_n497), .A3(G200), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n494), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n492), .A2(new_n376), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n500), .B(new_n473), .C1(G179), .C2(new_n492), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(KEYINPUT81), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT81), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n499), .A2(new_n504), .A3(new_n501), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(G116), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n312), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g0308(.A1(G238), .A2(G1698), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n509), .B1(new_n221), .B2(G1698), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n508), .B1(new_n272), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n278), .B1(G250), .B2(new_n486), .ZN(new_n512));
  NOR3_X1   g0312(.A1(new_n485), .A2(G1), .A3(G274), .ZN(new_n513));
  OAI22_X1  g0313(.A1(new_n511), .A2(new_n278), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n514), .A2(G179), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n514), .A2(new_n376), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT19), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n518), .A2(new_n229), .A3(G33), .A4(G97), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n464), .A2(new_n209), .B1(new_n429), .B2(new_n229), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n519), .B1(new_n520), .B2(new_n518), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n300), .A2(new_n229), .A3(G68), .A4(new_n270), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(KEYINPUT82), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT82), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n521), .A2(new_n522), .A3(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n524), .A2(new_n259), .A3(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n381), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n528), .A2(new_n255), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(KEYINPUT83), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT83), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n527), .A2(new_n533), .A3(new_n530), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n470), .A2(new_n381), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n516), .B(new_n517), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n514), .A2(new_n392), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT84), .ZN(new_n540));
  XNOR2_X1  g0340(.A(new_n539), .B(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n514), .A2(new_n394), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n470), .A2(new_n209), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n541), .A2(new_n535), .A3(new_n542), .A4(new_n544), .ZN(new_n545));
  NOR3_X1   g0345(.A1(new_n229), .A2(KEYINPUT23), .A3(G107), .ZN(new_n546));
  XNOR2_X1  g0346(.A(new_n546), .B(KEYINPUT87), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n270), .A2(new_n311), .A3(new_n229), .A4(G87), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT22), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT86), .ZN(new_n551));
  OR2_X1    g0351(.A1(new_n551), .A2(KEYINPUT23), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(KEYINPUT23), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n552), .B(new_n553), .C1(new_n229), .C2(G107), .ZN(new_n554));
  AND3_X1   g0354(.A1(new_n547), .A2(new_n550), .A3(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n272), .A2(KEYINPUT22), .A3(new_n229), .A4(G87), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n508), .A2(new_n229), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n555), .A2(KEYINPUT24), .A3(new_n556), .A4(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT24), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n557), .A2(new_n547), .A3(new_n550), .A4(new_n554), .ZN(new_n560));
  NOR4_X1   g0360(.A1(new_n475), .A2(new_n549), .A3(G20), .A4(new_n209), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n558), .A2(new_n562), .A3(new_n259), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n471), .A2(G107), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n255), .A2(G107), .ZN(new_n565));
  XNOR2_X1  g0365(.A(new_n565), .B(KEYINPUT25), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n563), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n210), .A2(new_n273), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n212), .A2(G1698), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n300), .A2(new_n270), .A3(new_n569), .A4(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n267), .A2(G294), .A3(new_n268), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n278), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n489), .A2(new_n278), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n574), .A2(new_n216), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n491), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n495), .ZN(new_n578));
  OR2_X1    g0378(.A1(new_n578), .A2(KEYINPUT88), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n578), .B(KEYINPUT88), .C1(G190), .C2(new_n577), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n568), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(G169), .B1(new_n576), .B2(new_n491), .ZN(new_n582));
  INV_X1    g0382(.A(new_n577), .ZN(new_n583));
  INV_X1    g0383(.A(G179), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n567), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n538), .A2(new_n545), .A3(new_n581), .A4(new_n586), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n574), .A2(new_n242), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n212), .A2(new_n273), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n216), .A2(G1698), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n300), .A2(new_n270), .A3(new_n589), .A4(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(G303), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n591), .B1(new_n592), .B2(new_n316), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n588), .B1(new_n593), .B2(new_n279), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n491), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n256), .A2(new_n507), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n480), .B(new_n229), .C1(G33), .C2(new_n211), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n597), .B(new_n259), .C1(new_n229), .C2(G116), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT20), .ZN(new_n599));
  AND2_X1   g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n598), .A2(new_n599), .ZN(new_n601));
  OAI221_X1 g0401(.A(new_n596), .B1(new_n507), .B2(new_n470), .C1(new_n600), .C2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n595), .A2(new_n602), .A3(G169), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT21), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n595), .A2(G200), .ZN(new_n606));
  INV_X1    g0406(.A(new_n602), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n606), .B(new_n607), .C1(new_n392), .C2(new_n595), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n595), .A2(KEYINPUT21), .A3(G169), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n594), .A2(G179), .A3(new_n491), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(KEYINPUT85), .B1(new_n611), .B2(new_n602), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT85), .ZN(new_n613));
  AOI211_X1 g0413(.A(new_n613), .B(new_n607), .C1(new_n609), .C2(new_n610), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n605), .B(new_n608), .C1(new_n612), .C2(new_n614), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n587), .A2(new_n615), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n460), .A2(new_n506), .A3(new_n616), .ZN(G372));
  INV_X1    g0417(.A(new_n438), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n437), .A2(new_n425), .A3(G169), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n618), .A2(new_n442), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n423), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT90), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n446), .A2(new_n447), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n621), .B(new_n622), .C1(new_n623), .C2(new_n458), .ZN(new_n624));
  INV_X1    g0424(.A(new_n334), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n623), .A2(new_n458), .ZN(new_n626));
  OAI21_X1  g0426(.A(KEYINPUT90), .B1(new_n443), .B2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n624), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n355), .A2(new_n358), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n409), .A2(new_n414), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n379), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n534), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n533), .B1(new_n527), .B2(new_n530), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n542), .B(new_n544), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n501), .B1(new_n636), .B2(new_n541), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT26), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n538), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  AOI211_X1 g0439(.A(new_n604), .B(new_n376), .C1(new_n594), .C2(new_n491), .ZN(new_n640));
  INV_X1    g0440(.A(new_n610), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n602), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n586), .A2(new_n605), .A3(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n499), .A2(new_n643), .A3(new_n581), .ZN(new_n644));
  AOI21_X1  g0444(.A(KEYINPUT26), .B1(new_n644), .B2(new_n501), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT89), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n539), .B1(new_n635), .B2(new_n646), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n535), .A2(KEYINPUT89), .A3(new_n542), .A4(new_n544), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n639), .B1(new_n645), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n632), .B1(new_n459), .B2(new_n650), .ZN(G369));
  NAND2_X1  g0451(.A1(new_n642), .A2(new_n605), .ZN(new_n652));
  INV_X1    g0452(.A(G13), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n653), .A2(G20), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  OR3_X1    g0455(.A1(new_n655), .A2(KEYINPUT27), .A3(G1), .ZN(new_n656));
  OAI21_X1  g0456(.A(KEYINPUT27), .B1(new_n655), .B2(G1), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n656), .A2(G213), .A3(new_n657), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n658), .A2(KEYINPUT91), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(KEYINPUT91), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(G343), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n663), .A2(new_n607), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n652), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n665), .B1(new_n615), .B2(new_n664), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n666), .A2(G330), .ZN(new_n667));
  INV_X1    g0467(.A(new_n663), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(new_n567), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n581), .A2(new_n586), .A3(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT92), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n581), .A2(KEYINPUT92), .A3(new_n586), .A4(new_n669), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n567), .A2(new_n585), .A3(new_n668), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n667), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n586), .A2(new_n668), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n672), .A2(new_n673), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n605), .B1(new_n612), .B2(new_n614), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(new_n663), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n677), .B1(new_n678), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n676), .A2(new_n682), .ZN(G399));
  NAND2_X1  g0483(.A1(new_n206), .A2(new_n277), .ZN(new_n684));
  XNOR2_X1  g0484(.A(new_n684), .B(KEYINPUT93), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n464), .A2(new_n209), .A3(new_n507), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AOI22_X1  g0487(.A1(new_n687), .A2(G1), .B1(new_n234), .B2(new_n685), .ZN(new_n688));
  XOR2_X1   g0488(.A(new_n688), .B(KEYINPUT28), .Z(new_n689));
  INV_X1    g0489(.A(KEYINPUT29), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n690), .B1(new_n650), .B2(new_n668), .ZN(new_n691));
  INV_X1    g0491(.A(new_n501), .ZN(new_n692));
  OAI211_X1 g0492(.A(new_n586), .B(new_n605), .C1(new_n612), .C2(new_n614), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n649), .A2(new_n693), .A3(new_n499), .A4(new_n581), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n692), .B1(new_n694), .B2(new_n638), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n637), .A2(new_n638), .ZN(new_n696));
  OAI211_X1 g0496(.A(new_n696), .B(new_n538), .C1(new_n638), .C2(new_n649), .ZN(new_n697));
  OAI211_X1 g0497(.A(KEYINPUT29), .B(new_n663), .C1(new_n695), .C2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n691), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(G330), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n506), .A2(new_n616), .A3(new_n663), .ZN(new_n701));
  NOR3_X1   g0501(.A1(new_n514), .A2(new_n575), .A3(new_n573), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n493), .A2(new_n641), .A3(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT30), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n493), .A2(new_n702), .A3(KEYINPUT30), .A4(new_n641), .ZN(new_n706));
  AOI21_X1  g0506(.A(G179), .B1(new_n594), .B2(new_n491), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n492), .A2(new_n514), .A3(new_n577), .A4(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n705), .A2(new_n706), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(new_n668), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n710), .B(KEYINPUT31), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n700), .B1(new_n701), .B2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n699), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n689), .B1(new_n715), .B2(G1), .ZN(G364));
  AOI21_X1  g0516(.A(new_n254), .B1(new_n654), .B2(G45), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n685), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n297), .A2(new_n302), .ZN(new_n721));
  INV_X1    g0521(.A(new_n206), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n234), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n723), .B1(G45), .B2(new_n724), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n725), .B(KEYINPUT95), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n726), .B1(new_n485), .B2(new_n247), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n722), .A2(new_n315), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(G355), .ZN(new_n729));
  OAI211_X1 g0529(.A(new_n727), .B(new_n729), .C1(G116), .C2(new_n206), .ZN(new_n730));
  NOR2_X1   g0530(.A1(G13), .A2(G33), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(G20), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n228), .B1(G20), .B2(new_n376), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XOR2_X1   g0535(.A(new_n735), .B(KEYINPUT96), .Z(new_n736));
  AOI21_X1  g0536(.A(new_n720), .B1(new_n730), .B2(new_n736), .ZN(new_n737));
  XOR2_X1   g0537(.A(new_n737), .B(KEYINPUT97), .Z(new_n738));
  NAND2_X1  g0538(.A1(new_n394), .A2(new_n584), .ZN(new_n739));
  NOR3_X1   g0539(.A1(new_n739), .A2(new_n229), .A3(new_n392), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(new_n209), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n584), .A2(new_n392), .A3(new_n495), .A4(G20), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT98), .ZN(new_n744));
  OR2_X1    g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n743), .A2(new_n744), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G159), .ZN(new_n749));
  OR2_X1    g0549(.A1(new_n749), .A2(KEYINPUT32), .ZN(new_n750));
  NOR3_X1   g0550(.A1(new_n392), .A2(G179), .A3(G200), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(new_n229), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  AOI22_X1  g0553(.A1(new_n749), .A2(KEYINPUT32), .B1(G97), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(G20), .A2(G179), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G190), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(G200), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n316), .B1(new_n759), .B2(new_n223), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n755), .A2(G190), .A3(G200), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n760), .B1(G77), .B2(new_n761), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n739), .A2(new_n229), .A3(G190), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n757), .A2(new_n495), .ZN(new_n764));
  AOI22_X1  g0564(.A1(new_n763), .A2(G107), .B1(G50), .B2(new_n764), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n750), .A2(new_n754), .A3(new_n762), .A4(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n756), .A2(new_n392), .A3(G200), .ZN(new_n767));
  OR2_X1    g0567(.A1(new_n767), .A2(KEYINPUT99), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(KEYINPUT99), .ZN(new_n769));
  AND2_X1   g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI211_X1 g0571(.A(new_n742), .B(new_n766), .C1(G68), .C2(new_n771), .ZN(new_n772));
  XNOR2_X1  g0572(.A(KEYINPUT33), .B(G317), .ZN(new_n773));
  AOI22_X1  g0573(.A1(new_n771), .A2(new_n773), .B1(G322), .B2(new_n758), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n774), .B1(new_n592), .B2(new_n741), .ZN(new_n775));
  AND2_X1   g0575(.A1(new_n764), .A2(G326), .ZN(new_n776));
  INV_X1    g0576(.A(G294), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n752), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n316), .B1(G311), .B2(new_n761), .ZN(new_n779));
  INV_X1    g0579(.A(G329), .ZN(new_n780));
  INV_X1    g0580(.A(new_n763), .ZN(new_n781));
  INV_X1    g0581(.A(G283), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n779), .B1(new_n780), .B2(new_n747), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  NOR4_X1   g0583(.A1(new_n775), .A2(new_n776), .A3(new_n778), .A4(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n734), .B1(new_n772), .B2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n733), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n738), .B(new_n785), .C1(new_n666), .C2(new_n786), .ZN(new_n787));
  AND3_X1   g0587(.A1(new_n666), .A2(KEYINPUT94), .A3(G330), .ZN(new_n788));
  AOI21_X1  g0588(.A(KEYINPUT94), .B1(new_n666), .B2(G330), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n720), .B1(G330), .B2(new_n666), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n787), .A2(new_n790), .ZN(G396));
  NOR2_X1   g0591(.A1(new_n650), .A2(new_n668), .ZN(new_n792));
  OR2_X1    g0592(.A1(new_n663), .A2(new_n386), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(new_n396), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(new_n458), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n456), .A2(new_n457), .A3(new_n663), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(KEYINPUT100), .ZN(new_n798));
  INV_X1    g0598(.A(KEYINPUT100), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n795), .A2(new_n799), .A3(new_n796), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n792), .B(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(new_n712), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(new_n720), .ZN(new_n804));
  INV_X1    g0604(.A(new_n734), .ZN(new_n805));
  AOI22_X1  g0605(.A1(G137), .A2(new_n764), .B1(new_n758), .B2(G143), .ZN(new_n806));
  INV_X1    g0606(.A(G159), .ZN(new_n807));
  INV_X1    g0607(.A(new_n761), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n806), .B1(new_n807), .B2(new_n808), .C1(new_n770), .C2(new_n369), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT34), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n763), .A2(G68), .B1(G58), .B2(new_n753), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n810), .A2(new_n721), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(G132), .B2(new_n748), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(new_n373), .B2(new_n741), .ZN(new_n814));
  INV_X1    g0614(.A(G311), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n315), .B1(new_n747), .B2(new_n815), .C1(new_n770), .C2(new_n782), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n816), .B1(G87), .B2(new_n763), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n761), .A2(G116), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n740), .A2(G107), .ZN(new_n819));
  INV_X1    g0619(.A(new_n764), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n759), .A2(new_n777), .B1(new_n820), .B2(new_n592), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n821), .B1(G97), .B2(new_n753), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n817), .A2(new_n818), .A3(new_n819), .A4(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n805), .B1(new_n814), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n734), .A2(new_n731), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n720), .B(new_n824), .C1(new_n220), .C2(new_n825), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(new_n732), .B2(new_n801), .ZN(new_n827));
  AND2_X1   g0627(.A1(new_n804), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(G384));
  NAND2_X1  g0629(.A1(new_n644), .A2(new_n501), .ZN(new_n830));
  AND3_X1   g0630(.A1(new_n830), .A2(new_n638), .A3(new_n649), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n801), .B(new_n663), .C1(new_n831), .C2(new_n639), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(new_n796), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT101), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n663), .A2(new_n424), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n623), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n621), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n835), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n837), .B1(new_n451), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n833), .A2(new_n834), .A3(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT38), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n342), .A2(new_n260), .ZN(new_n842));
  OR2_X1    g0642(.A1(new_n356), .A2(KEYINPUT16), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n263), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  OR2_X1    g0644(.A1(new_n844), .A2(new_n661), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n354), .A2(new_n359), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n845), .B1(new_n846), .B2(new_n625), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n348), .A2(new_n662), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n332), .B1(new_n844), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(KEYINPUT37), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n661), .B(KEYINPUT102), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n345), .B1(new_n348), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT37), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n853), .A2(new_n854), .A3(new_n332), .ZN(new_n855));
  AND2_X1   g0655(.A1(new_n850), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n841), .B1(new_n847), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n850), .A2(new_n855), .ZN(new_n858));
  OAI211_X1 g0658(.A(KEYINPUT38), .B(new_n858), .C1(new_n360), .C2(new_n845), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n796), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n861), .B1(new_n792), .B2(new_n801), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n450), .A2(new_n448), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n621), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n864), .A2(new_n835), .B1(new_n621), .B2(new_n836), .ZN(new_n865));
  OAI21_X1  g0665(.A(KEYINPUT101), .B1(new_n862), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n840), .A2(new_n860), .A3(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n629), .A2(new_n328), .A3(new_n333), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n350), .A2(new_n851), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n332), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n329), .A2(new_n331), .B1(new_n352), .B2(new_n851), .ZN(new_n872));
  OAI21_X1  g0672(.A(KEYINPUT37), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n873), .A2(KEYINPUT103), .A3(new_n855), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT103), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n875), .B(KEYINPUT37), .C1(new_n871), .C2(new_n872), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n870), .A2(new_n874), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n841), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n859), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT39), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n621), .A2(new_n668), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n857), .A2(KEYINPUT39), .A3(new_n859), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n867), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n355), .A2(new_n358), .A3(new_n851), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n630), .A2(new_n631), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n378), .ZN(new_n889));
  AND2_X1   g0689(.A1(new_n691), .A2(new_n698), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n890), .A2(KEYINPUT104), .A3(new_n460), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT104), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(new_n699), .B2(new_n459), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n889), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n887), .B(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT40), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n701), .A2(new_n711), .ZN(new_n897));
  AND3_X1   g0697(.A1(new_n839), .A2(new_n897), .A3(new_n801), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n896), .B1(new_n898), .B2(new_n879), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n839), .A2(new_n896), .A3(new_n897), .A4(new_n801), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n900), .B1(new_n859), .B2(new_n857), .ZN(new_n901));
  OAI21_X1  g0701(.A(G330), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n460), .A2(new_n712), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n897), .B1(new_n899), .B2(new_n901), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n904), .B1(new_n459), .B2(new_n905), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n895), .B(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n254), .B2(new_n654), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT35), .ZN(new_n909));
  AOI211_X1 g0709(.A(new_n229), .B(new_n228), .C1(new_n467), .C2(new_n909), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n910), .B(G116), .C1(new_n909), .C2(new_n467), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n911), .B(KEYINPUT36), .ZN(new_n912));
  NOR3_X1   g0712(.A1(new_n724), .A2(new_n220), .A3(new_n293), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n231), .A2(G50), .ZN(new_n914));
  OAI211_X1 g0714(.A(G1), .B(new_n653), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n908), .A2(new_n912), .A3(new_n915), .ZN(G367));
  AOI21_X1  g0716(.A(new_n680), .B1(new_n672), .B2(new_n673), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n917), .A2(new_n499), .A3(new_n501), .ZN(new_n918));
  OR2_X1    g0718(.A1(new_n918), .A2(KEYINPUT42), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(KEYINPUT42), .ZN(new_n920));
  AND2_X1   g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT43), .ZN(new_n922));
  INV_X1    g0722(.A(new_n538), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n668), .B1(new_n536), .B2(new_n543), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n649), .A2(new_n924), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n925), .B1(new_n926), .B2(new_n923), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(KEYINPUT105), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT105), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n929), .B(new_n925), .C1(new_n926), .C2(new_n923), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n668), .A2(new_n473), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n499), .A2(new_n501), .A3(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n501), .B1(new_n934), .B2(new_n586), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n663), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n921), .A2(new_n922), .A3(new_n932), .A4(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n692), .A2(new_n668), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n934), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n676), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n919), .A2(new_n936), .A3(new_n920), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n931), .A2(KEYINPUT43), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n928), .A2(new_n930), .A3(new_n922), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n937), .A2(new_n941), .A3(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT106), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n937), .A2(new_n945), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n676), .B2(new_n940), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n685), .B(KEYINPUT41), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT109), .ZN(new_n952));
  OAI21_X1  g0752(.A(KEYINPUT44), .B1(new_n682), .B2(new_n939), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT44), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n954), .B(new_n940), .C1(new_n917), .C2(new_n677), .ZN(new_n955));
  AOI21_X1  g0755(.A(KEYINPUT45), .B1(new_n682), .B2(new_n939), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT45), .ZN(new_n957));
  NOR4_X1   g0757(.A1(new_n917), .A2(new_n940), .A3(new_n957), .A4(new_n677), .ZN(new_n958));
  OAI211_X1 g0758(.A(new_n953), .B(new_n955), .C1(new_n956), .C2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n676), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n952), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  AND2_X1   g0761(.A1(new_n953), .A2(new_n955), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n682), .A2(new_n939), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n957), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n682), .A2(KEYINPUT45), .A3(new_n939), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n962), .A2(new_n966), .A3(KEYINPUT109), .A4(new_n676), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n961), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n678), .A2(new_n681), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n672), .A2(new_n680), .A3(new_n673), .A4(new_n674), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n788), .B2(new_n789), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(KEYINPUT108), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n667), .A2(new_n969), .A3(new_n970), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT108), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n971), .B(new_n975), .C1(new_n789), .C2(new_n788), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n973), .A2(new_n974), .A3(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n977), .A2(new_n714), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n959), .A2(new_n960), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(KEYINPUT107), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT107), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n959), .A2(new_n981), .A3(new_n960), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n968), .A2(new_n978), .A3(new_n980), .A4(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n951), .B1(new_n983), .B2(new_n715), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n947), .B(new_n949), .C1(new_n984), .C2(new_n718), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n932), .A2(new_n733), .ZN(new_n986));
  INV_X1    g0786(.A(G317), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n747), .A2(new_n987), .B1(new_n820), .B2(new_n815), .ZN(new_n988));
  AOI211_X1 g0788(.A(new_n721), .B(new_n988), .C1(G303), .C2(new_n758), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n771), .A2(G294), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n740), .A2(G116), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT46), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n752), .A2(new_n215), .B1(new_n808), .B2(new_n782), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(new_n763), .B2(G97), .ZN(new_n994));
  NAND4_X1  g0794(.A1(new_n989), .A2(new_n990), .A3(new_n992), .A4(new_n994), .ZN(new_n995));
  AOI22_X1  g0795(.A1(G143), .A2(new_n764), .B1(new_n758), .B2(G150), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n231), .B2(new_n752), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT110), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n763), .A2(G77), .ZN(new_n999));
  XNOR2_X1  g0799(.A(KEYINPUT111), .B(G137), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n748), .A2(new_n1000), .ZN(new_n1001));
  AND4_X1   g0801(.A1(new_n316), .A2(new_n998), .A3(new_n999), .A4(new_n1001), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n1002), .B1(new_n373), .B2(new_n808), .C1(new_n807), .C2(new_n770), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n741), .A2(new_n223), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n995), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT47), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(new_n734), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n723), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n735), .B1(new_n206), .B2(new_n381), .C1(new_n243), .C2(new_n1008), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n986), .A2(new_n719), .A3(new_n1007), .A4(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n985), .A2(new_n1010), .ZN(G387));
  INV_X1    g0811(.A(new_n978), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n977), .A2(new_n714), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n685), .B(KEYINPUT112), .Z(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1012), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n977), .A2(new_n717), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1008), .B1(new_n239), .B2(G45), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(new_n686), .B2(new_n728), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n253), .A2(new_n373), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT50), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n485), .B1(new_n231), .B2(new_n220), .ZN(new_n1022));
  NOR3_X1   g0822(.A1(new_n1021), .A2(new_n686), .A3(new_n1022), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n1019), .A2(new_n1023), .B1(G107), .B2(new_n206), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(new_n736), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n675), .A2(new_n786), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n741), .A2(new_n220), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n770), .A2(new_n252), .B1(new_n373), .B2(new_n759), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n1027), .B(new_n1028), .C1(G159), .C2(new_n764), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n748), .A2(G150), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n721), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n752), .A2(new_n381), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n763), .A2(G97), .B1(G68), .B2(new_n761), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1029), .A2(new_n1030), .A3(new_n1033), .A4(new_n1034), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n758), .A2(G317), .B1(G303), .B2(new_n761), .ZN(new_n1036));
  INV_X1    g0836(.A(G322), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1036), .B1(new_n1037), .B2(new_n820), .C1(new_n770), .C2(new_n815), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT48), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1039), .B1(new_n782), .B2(new_n752), .C1(new_n777), .C2(new_n741), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT49), .ZN(new_n1041));
  OR2_X1    g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n748), .A2(G326), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n763), .A2(G116), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1042), .A2(new_n1031), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1035), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n720), .B(new_n1026), .C1(new_n1047), .C2(new_n734), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1017), .B1(new_n1025), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1016), .A2(new_n1049), .ZN(G393));
  AOI22_X1  g0850(.A1(G311), .A2(new_n758), .B1(new_n764), .B2(G317), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT52), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(G107), .A2(new_n763), .B1(new_n740), .B2(G283), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1053), .B(new_n315), .C1(new_n1037), .C2(new_n747), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT114), .Z(new_n1055));
  AOI211_X1 g0855(.A(new_n1052), .B(new_n1055), .C1(G116), .C2(new_n753), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n1056), .B1(new_n777), .B2(new_n808), .C1(new_n592), .C2(new_n770), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(G150), .A2(new_n764), .B1(new_n758), .B2(G159), .ZN(new_n1058));
  XOR2_X1   g0858(.A(KEYINPUT113), .B(KEYINPUT51), .Z(new_n1059));
  XNOR2_X1  g0859(.A(new_n1058), .B(new_n1059), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n741), .A2(new_n231), .B1(new_n252), .B2(new_n808), .ZN(new_n1061));
  NOR3_X1   g0861(.A1(new_n1060), .A2(new_n1031), .A3(new_n1061), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n748), .A2(G143), .B1(new_n763), .B2(G87), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n753), .A2(G77), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n771), .A2(G50), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n805), .B1(new_n1057), .B2(new_n1066), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n735), .B1(new_n211), .B2(new_n206), .C1(new_n1008), .C2(new_n250), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(new_n1069));
  NOR3_X1   g0869(.A1(new_n1067), .A2(new_n720), .A3(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n786), .B2(new_n939), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n968), .A2(new_n979), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1071), .B1(new_n1072), .B2(new_n717), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1014), .B1(new_n1072), .B2(new_n1012), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1073), .B1(new_n983), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(G390));
  NAND3_X1  g0876(.A1(new_n712), .A2(new_n839), .A3(new_n801), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n882), .B1(new_n833), .B2(new_n839), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(new_n881), .B2(new_n883), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n801), .B(new_n663), .C1(new_n695), .C2(new_n697), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(new_n796), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n839), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n882), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1083), .A2(new_n879), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1078), .B1(new_n1080), .B2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1084), .B1(new_n862), .B2(new_n865), .ZN(new_n1088));
  AND3_X1   g0888(.A1(new_n857), .A2(KEYINPUT39), .A3(new_n859), .ZN(new_n1089));
  AOI21_X1  g0889(.A(KEYINPUT39), .B1(new_n878), .B2(new_n859), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1088), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1091), .A2(new_n1085), .A3(new_n1077), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1087), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(KEYINPUT104), .B1(new_n890), .B2(new_n460), .ZN(new_n1094));
  NOR3_X1   g0894(.A1(new_n699), .A2(new_n459), .A3(new_n892), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n632), .B(new_n903), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n897), .A2(G330), .A3(new_n801), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n865), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT115), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1099), .A2(new_n1100), .A3(new_n1077), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1098), .A2(KEYINPUT115), .A3(new_n865), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1101), .A2(new_n833), .A3(new_n1102), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1099), .A2(new_n796), .A3(new_n1077), .A4(new_n1081), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1097), .A2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g0906(.A(KEYINPUT116), .B1(new_n1093), .B2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1096), .B1(new_n1104), .B2(new_n1103), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT116), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1108), .A2(new_n1109), .A3(new_n1087), .A4(new_n1092), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1107), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1014), .B1(new_n1093), .B2(new_n1106), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1087), .A2(new_n1092), .A3(new_n718), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n731), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1115));
  XOR2_X1   g0915(.A(KEYINPUT54), .B(G143), .Z(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n781), .A2(new_n373), .B1(new_n808), .B2(new_n1117), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n315), .B(new_n1118), .C1(G132), .C2(new_n758), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n753), .A2(G159), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n771), .A2(new_n1000), .B1(new_n748), .B2(G125), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n740), .A2(G150), .ZN(new_n1122));
  XOR2_X1   g0922(.A(new_n1122), .B(KEYINPUT53), .Z(new_n1123));
  NAND4_X1  g0923(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .A4(new_n1123), .ZN(new_n1124));
  AND2_X1   g0924(.A1(new_n764), .A2(G128), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n808), .A2(new_n211), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n771), .A2(G107), .B1(G68), .B2(new_n763), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n742), .A2(new_n316), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1064), .B1(new_n747), .B2(new_n777), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(G283), .B2(new_n764), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n758), .A2(G116), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n1127), .A2(new_n1128), .A3(new_n1130), .A4(new_n1131), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n1124), .A2(new_n1125), .B1(new_n1126), .B2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n720), .B1(new_n1133), .B2(new_n734), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n825), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1115), .B(new_n1134), .C1(new_n253), .C2(new_n1135), .ZN(new_n1136));
  AND2_X1   g0936(.A1(new_n1114), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1113), .A2(new_n1137), .ZN(G378));
  NAND2_X1  g0938(.A1(new_n1111), .A2(new_n1097), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n631), .A2(new_n378), .ZN(new_n1140));
  XOR2_X1   g0940(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1141));
  XNOR2_X1  g0941(.A(new_n1140), .B(new_n1141), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n400), .A2(new_n661), .ZN(new_n1143));
  XOR2_X1   g0943(.A(new_n1142), .B(new_n1143), .Z(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n902), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1144), .B(G330), .C1(new_n899), .C2(new_n901), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n887), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1146), .A2(new_n1147), .A3(new_n885), .A4(new_n886), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1139), .A2(KEYINPUT57), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT57), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1096), .B1(new_n1107), .B2(new_n1110), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1154), .B1(new_n1155), .B2(new_n1151), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1153), .A2(new_n1015), .A3(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1144), .A2(new_n731), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1135), .A2(G50), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n1031), .B1(new_n215), .B2(new_n759), .C1(new_n782), .C2(new_n747), .ZN(new_n1160));
  OAI221_X1 g0960(.A(new_n277), .B1(new_n808), .B2(new_n381), .C1(new_n781), .C2(new_n223), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n752), .A2(new_n231), .ZN(new_n1162));
  NOR4_X1   g0962(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .A4(new_n1027), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n1163), .B1(new_n211), .B2(new_n770), .C1(new_n507), .C2(new_n820), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1164), .B(KEYINPUT58), .ZN(new_n1165));
  AOI21_X1  g0965(.A(G41), .B1(new_n721), .B2(G33), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n741), .A2(new_n1117), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n1168), .A2(KEYINPUT117), .B1(G137), .B2(new_n761), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n753), .A2(G150), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n758), .A2(G128), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT117), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n1167), .A2(new_n1172), .B1(new_n771), .B2(G132), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .A4(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(G125), .B2(new_n764), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT59), .ZN(new_n1176));
  AOI21_X1  g0976(.A(G33), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(G41), .B1(new_n748), .B2(G124), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1177), .B(new_n1178), .C1(new_n807), .C2(new_n781), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n1165), .B1(G50), .B2(new_n1166), .C1(new_n1179), .C2(new_n1180), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1181), .B(KEYINPUT118), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n720), .B(new_n1159), .C1(new_n1182), .C2(new_n734), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1158), .A2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(new_n1151), .B2(new_n717), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1157), .A2(new_n1186), .ZN(G375));
  AOI21_X1  g0987(.A(KEYINPUT119), .B1(new_n1105), .B2(new_n718), .ZN(new_n1188));
  AND3_X1   g0988(.A1(new_n1105), .A2(KEYINPUT119), .A3(new_n718), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n865), .A2(new_n731), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1032), .B1(G283), .B2(new_n758), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(new_n777), .B2(new_n820), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n748), .A2(G303), .B1(new_n740), .B2(G97), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n1193), .B(KEYINPUT120), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n1192), .B(new_n1194), .C1(G107), .C2(new_n761), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n771), .A2(G116), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1195), .A2(new_n315), .A3(new_n999), .A4(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n758), .A2(new_n1000), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1198), .B1(new_n781), .B2(new_n223), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n752), .A2(new_n373), .B1(new_n808), .B2(new_n369), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n1200), .B(KEYINPUT121), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n1199), .B(new_n1201), .C1(new_n771), .C2(new_n1116), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n764), .A2(G132), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n748), .A2(G128), .B1(new_n740), .B2(G159), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1202), .A2(new_n721), .A3(new_n1203), .A4(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n805), .B1(new_n1197), .B2(new_n1205), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n720), .B(new_n1206), .C1(new_n231), .C2(new_n825), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n1188), .B(new_n1189), .C1(new_n1190), .C2(new_n1207), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n950), .B1(new_n1097), .B2(new_n1105), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1208), .B1(new_n1108), .B2(new_n1209), .ZN(G381));
  AOI21_X1  g1010(.A(new_n1151), .B1(new_n1111), .B2(new_n1097), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1014), .B1(new_n1211), .B2(KEYINPUT57), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1185), .B1(new_n1212), .B2(new_n1156), .ZN(new_n1213));
  INV_X1    g1013(.A(G378), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  NOR3_X1   g1015(.A1(new_n1215), .A2(G384), .A3(G381), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n985), .A2(new_n1010), .A3(new_n1075), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1016), .A2(new_n1049), .A3(new_n787), .A4(new_n790), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1216), .A2(new_n1217), .A3(new_n1219), .ZN(G407));
  OAI211_X1 g1020(.A(G407), .B(G213), .C1(G343), .C2(new_n1215), .ZN(G409));
  AOI21_X1  g1021(.A(new_n1075), .B1(new_n985), .B2(new_n1010), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT122), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(G393), .A2(G396), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1223), .B1(new_n1224), .B2(new_n1218), .ZN(new_n1225));
  AND3_X1   g1025(.A1(new_n1224), .A2(new_n1223), .A3(new_n1218), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n1217), .A2(new_n1222), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(G387), .A2(G390), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n985), .A2(new_n1010), .A3(new_n1075), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1226), .A2(new_n1225), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1228), .A2(new_n1229), .A3(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1227), .A2(new_n1231), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(new_n1232), .B(KEYINPUT125), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT61), .ZN(new_n1234));
  NOR3_X1   g1034(.A1(new_n1155), .A2(new_n951), .A3(new_n1151), .ZN(new_n1235));
  OR3_X1    g1035(.A1(new_n1235), .A2(G378), .A3(new_n1185), .ZN(new_n1236));
  INV_X1    g1036(.A(G213), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1237), .A2(G343), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1236), .B(new_n1239), .C1(new_n1213), .C2(new_n1214), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1097), .A2(new_n1105), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1014), .B1(new_n1241), .B2(KEYINPUT60), .ZN(new_n1242));
  AND2_X1   g1042(.A1(new_n1106), .A2(KEYINPUT60), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1242), .B1(new_n1243), .B2(new_n1241), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1208), .A2(G384), .A3(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(G384), .B1(new_n1208), .B2(new_n1244), .ZN(new_n1247));
  OAI211_X1 g1047(.A(G2897), .B(new_n1238), .C1(new_n1246), .C2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1247), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1238), .A2(G2897), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1249), .A2(new_n1245), .A3(new_n1250), .ZN(new_n1251));
  AND2_X1   g1051(.A1(new_n1248), .A2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(KEYINPUT62), .B1(new_n1240), .B2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1214), .B1(new_n1157), .B2(new_n1186), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1249), .A2(new_n1245), .ZN(new_n1255));
  NOR3_X1   g1055(.A1(new_n1235), .A2(G378), .A3(new_n1185), .ZN(new_n1256));
  NOR4_X1   g1056(.A1(new_n1254), .A2(new_n1255), .A3(new_n1238), .A4(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1234), .B1(new_n1253), .B2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(G375), .A2(G378), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1259), .A2(new_n1260), .A3(new_n1239), .A4(new_n1236), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1261), .A2(KEYINPUT62), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1233), .B1(new_n1258), .B2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1240), .A2(new_n1252), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1257), .B1(new_n1264), .B2(KEYINPUT63), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT63), .ZN(new_n1266));
  AOI21_X1  g1066(.A(KEYINPUT123), .B1(new_n1232), .B2(new_n1234), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT123), .ZN(new_n1268));
  AOI211_X1 g1068(.A(new_n1268), .B(KEYINPUT61), .C1(new_n1227), .C2(new_n1231), .ZN(new_n1269));
  OAI22_X1  g1069(.A1(new_n1261), .A2(new_n1266), .B1(new_n1267), .B2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT124), .ZN(new_n1271));
  NOR3_X1   g1071(.A1(new_n1265), .A2(new_n1270), .A3(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1248), .A2(new_n1251), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1238), .B1(G375), .B2(G378), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1273), .B1(new_n1274), .B2(new_n1236), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1261), .B1(new_n1275), .B2(new_n1266), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1267), .A2(new_n1269), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1277), .B1(new_n1257), .B2(KEYINPUT63), .ZN(new_n1278));
  AOI21_X1  g1078(.A(KEYINPUT124), .B1(new_n1276), .B2(new_n1278), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1263), .B1(new_n1272), .B2(new_n1279), .ZN(G405));
  INV_X1    g1080(.A(KEYINPUT127), .ZN(new_n1281));
  AND3_X1   g1081(.A1(new_n1260), .A2(KEYINPUT126), .A3(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1281), .B1(new_n1260), .B2(KEYINPUT126), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1259), .A2(new_n1215), .ZN(new_n1285));
  OR2_X1    g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1232), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1288));
  AND3_X1   g1088(.A1(new_n1286), .A2(new_n1287), .A3(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1287), .B1(new_n1286), .B2(new_n1288), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1289), .A2(new_n1290), .ZN(G402));
endmodule


