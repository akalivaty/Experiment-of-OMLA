//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 1 1 0 0 0 0 1 1 1 0 0 0 1 0 0 1 0 1 1 0 1 1 1 1 0 1 0 0 1 1 1 0 1 1 1 0 1 0 0 1 1 0 1 1 1 0 0 0 0 0 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:34 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n542, new_n543, new_n544, new_n545, new_n546, new_n548,
    new_n549, new_n550, new_n551, new_n554, new_n555, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n577, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n613, new_n616, new_n618, new_n619,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1201, new_n1202,
    new_n1203;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT64), .Z(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n455), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n453), .A2(G2106), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n458), .B1(new_n459), .B2(KEYINPUT65), .ZN(new_n460));
  AOI21_X1  g035(.A(new_n460), .B1(KEYINPUT65), .B2(new_n459), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT66), .Z(G319));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT67), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT67), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n464), .A2(new_n466), .A3(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  OAI21_X1  g043(.A(KEYINPUT68), .B1(new_n463), .B2(KEYINPUT3), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT68), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n470), .A2(new_n471), .A3(G2104), .ZN(new_n472));
  NAND4_X1  g047(.A1(new_n467), .A2(new_n468), .A3(new_n469), .A4(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G137), .ZN(new_n474));
  XNOR2_X1  g049(.A(KEYINPUT3), .B(G2104), .ZN(new_n475));
  AOI22_X1  g050(.A1(new_n475), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n476));
  OAI22_X1  g051(.A1(new_n473), .A2(new_n474), .B1(new_n476), .B2(new_n468), .ZN(new_n477));
  INV_X1    g052(.A(G101), .ZN(new_n478));
  XNOR2_X1  g053(.A(KEYINPUT67), .B(G2104), .ZN(new_n479));
  OAI21_X1  g054(.A(KEYINPUT69), .B1(new_n479), .B2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n464), .A2(new_n466), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT69), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n481), .A2(new_n482), .A3(new_n468), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n478), .B1(new_n480), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n477), .A2(new_n484), .ZN(G160));
  NAND4_X1  g060(.A1(new_n467), .A2(G2105), .A3(new_n469), .A4(new_n472), .ZN(new_n486));
  INV_X1    g061(.A(G124), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n468), .A2(G112), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n489));
  OAI22_X1  g064(.A1(new_n486), .A2(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(G136), .ZN(new_n491));
  OR3_X1    g066(.A1(new_n473), .A2(KEYINPUT70), .A3(new_n491), .ZN(new_n492));
  OAI21_X1  g067(.A(KEYINPUT70), .B1(new_n473), .B2(new_n491), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n490), .B1(new_n492), .B2(new_n493), .ZN(G162));
  INV_X1    g069(.A(G126), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n468), .A2(G114), .ZN(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n497));
  OAI22_X1  g072(.A1(new_n486), .A2(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n471), .A2(G2104), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n502), .A2(new_n468), .A3(G138), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  AND2_X1   g079(.A1(new_n468), .A2(G138), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n467), .A2(new_n469), .A3(new_n472), .A4(new_n505), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n504), .B1(new_n506), .B2(KEYINPUT4), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n498), .A2(new_n507), .ZN(G164));
  INV_X1    g083(.A(KEYINPUT71), .ZN(new_n509));
  OR2_X1    g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  AND2_X1   g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  AND2_X1   g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  OAI22_X1  g094(.A1(new_n516), .A2(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G88), .ZN(new_n521));
  OAI21_X1  g096(.A(G543), .B1(new_n518), .B2(new_n519), .ZN(new_n522));
  INV_X1    g097(.A(G50), .ZN(new_n523));
  OAI22_X1  g098(.A1(new_n520), .A2(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n509), .B1(new_n515), .B2(new_n524), .ZN(new_n525));
  OR2_X1    g100(.A1(KEYINPUT6), .A2(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(KEYINPUT6), .A2(G651), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n510), .A2(new_n511), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(G543), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n529), .B1(new_n526), .B2(new_n527), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n528), .A2(G88), .B1(new_n530), .B2(G50), .ZN(new_n531));
  OAI211_X1 g106(.A(new_n531), .B(KEYINPUT71), .C1(new_n514), .C2(new_n513), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n525), .A2(new_n532), .ZN(G166));
  XNOR2_X1  g108(.A(KEYINPUT72), .B(KEYINPUT7), .ZN(new_n534));
  AND3_X1   g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n534), .B(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n512), .A2(G63), .A3(G651), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n530), .A2(G51), .ZN(new_n538));
  XOR2_X1   g113(.A(KEYINPUT73), .B(G89), .Z(new_n539));
  NAND2_X1  g114(.A1(new_n528), .A2(new_n539), .ZN(new_n540));
  AND4_X1   g115(.A1(new_n536), .A2(new_n537), .A3(new_n538), .A4(new_n540), .ZN(G168));
  AOI22_X1  g116(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(new_n514), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n530), .A2(G52), .ZN(new_n544));
  INV_X1    g119(.A(G90), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n545), .B2(new_n520), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n543), .A2(new_n546), .ZN(G171));
  AOI22_X1  g122(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n548));
  OR2_X1    g123(.A1(new_n548), .A2(new_n514), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n528), .A2(G81), .B1(new_n530), .B2(G43), .ZN(new_n550));
  AND2_X1   g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  INV_X1    g131(.A(G53), .ZN(new_n557));
  OAI21_X1  g132(.A(KEYINPUT9), .B1(new_n522), .B2(new_n557), .ZN(new_n558));
  OR3_X1    g133(.A1(new_n522), .A2(KEYINPUT9), .A3(new_n557), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n528), .A2(KEYINPUT74), .A3(G91), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT74), .ZN(new_n561));
  INV_X1    g136(.A(G91), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n520), .B2(new_n562), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n558), .A2(new_n559), .B1(new_n560), .B2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(G65), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT75), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n512), .A2(new_n566), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n517), .A2(new_n516), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(KEYINPUT75), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n565), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  AND2_X1   g145(.A1(G78), .A2(G543), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n564), .A2(new_n572), .ZN(G299));
  OAI221_X1 g148(.A(new_n544), .B1(new_n545), .B2(new_n520), .C1(new_n542), .C2(new_n514), .ZN(G301));
  NAND4_X1  g149(.A1(new_n536), .A2(new_n537), .A3(new_n538), .A4(new_n540), .ZN(G286));
  INV_X1    g150(.A(G166), .ZN(G303));
  INV_X1    g151(.A(G74), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n510), .A2(new_n577), .A3(new_n511), .ZN(new_n578));
  AOI22_X1  g153(.A1(G49), .A2(new_n530), .B1(new_n578), .B2(G651), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n528), .A2(G87), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(G288));
  INV_X1    g156(.A(G86), .ZN(new_n582));
  INV_X1    g157(.A(G48), .ZN(new_n583));
  OAI22_X1  g158(.A1(new_n520), .A2(new_n582), .B1(new_n522), .B2(new_n583), .ZN(new_n584));
  OAI21_X1  g159(.A(G61), .B1(new_n517), .B2(new_n516), .ZN(new_n585));
  NAND2_X1  g160(.A1(G73), .A2(G543), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n514), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G305));
  AND2_X1   g164(.A1(G72), .A2(G543), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n590), .B1(new_n512), .B2(G60), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n591), .A2(new_n514), .ZN(new_n592));
  INV_X1    g167(.A(G85), .ZN(new_n593));
  INV_X1    g168(.A(G47), .ZN(new_n594));
  OAI22_X1  g169(.A1(new_n520), .A2(new_n593), .B1(new_n522), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n530), .A2(G54), .ZN(new_n599));
  INV_X1    g174(.A(G92), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n520), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n601), .A2(KEYINPUT10), .ZN(new_n602));
  AND3_X1   g177(.A1(new_n528), .A2(KEYINPUT10), .A3(G92), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n599), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n567), .A2(new_n569), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(G66), .ZN(new_n606));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n514), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n598), .B1(new_n609), .B2(G868), .ZN(G284));
  OAI21_X1  g185(.A(new_n598), .B1(new_n609), .B2(G868), .ZN(G321));
  NAND2_X1  g186(.A1(G286), .A2(G868), .ZN(new_n612));
  INV_X1    g187(.A(G299), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(G868), .ZN(G297));
  XNOR2_X1  g189(.A(G297), .B(KEYINPUT76), .ZN(G280));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n609), .B1(new_n616), .B2(G860), .ZN(G148));
  NAND2_X1  g192(.A1(new_n609), .A2(new_n616), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(G868), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(G868), .B2(new_n551), .ZN(G323));
  XNOR2_X1  g195(.A(KEYINPUT77), .B(KEYINPUT11), .ZN(new_n621));
  XNOR2_X1  g196(.A(G323), .B(new_n621), .ZN(G282));
  INV_X1    g197(.A(new_n473), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(G135), .ZN(new_n624));
  AND4_X1   g199(.A1(G2105), .A2(new_n467), .A3(new_n469), .A4(new_n472), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G123), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n468), .A2(G111), .ZN(new_n627));
  OAI21_X1  g202(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n628));
  OAI211_X1 g203(.A(new_n624), .B(new_n626), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(KEYINPUT79), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n631), .A2(G2096), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n631), .A2(G2096), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n480), .A2(new_n483), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(new_n475), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT12), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT78), .B(G2100), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT13), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n636), .B(new_n638), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n632), .A2(new_n633), .A3(new_n639), .ZN(G156));
  INV_X1    g215(.A(KEYINPUT14), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2427), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2430), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT15), .B(G2435), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n641), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n645), .B1(new_n644), .B2(new_n643), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2451), .B(G2454), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT16), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n646), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(G14), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n651), .A2(new_n652), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(G401));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT80), .ZN(new_n658));
  NOR2_X1   g233(.A1(G2072), .A2(G2078), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n442), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2084), .B(G2090), .ZN(new_n661));
  NOR3_X1   g236(.A1(new_n658), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT18), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n658), .A2(new_n660), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n660), .B(KEYINPUT17), .ZN(new_n665));
  OAI211_X1 g240(.A(new_n664), .B(new_n661), .C1(new_n658), .C2(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n661), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n665), .A2(new_n658), .A3(new_n667), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n663), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(G2096), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT81), .B(G2100), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(G227));
  XOR2_X1   g247(.A(G1991), .B(G1996), .Z(new_n673));
  XNOR2_X1  g248(.A(G1971), .B(G1976), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G1956), .B(G2474), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT82), .ZN(new_n678));
  XOR2_X1   g253(.A(G1961), .B(G1966), .Z(new_n679));
  NAND3_X1  g254(.A1(new_n676), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT20), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n676), .B1(new_n678), .B2(new_n679), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n678), .A2(new_n679), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OAI211_X1 g259(.A(new_n681), .B(new_n684), .C1(new_n675), .C2(new_n683), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT83), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n685), .A2(new_n686), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n687), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n689), .B1(new_n687), .B2(new_n688), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n673), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n692), .ZN(new_n694));
  INV_X1    g269(.A(new_n673), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n694), .A2(new_n695), .A3(new_n690), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1981), .B(G1986), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n693), .A2(new_n696), .A3(new_n698), .ZN(new_n701));
  AND2_X1   g276(.A1(new_n700), .A2(new_n701), .ZN(G229));
  XOR2_X1   g277(.A(KEYINPUT92), .B(KEYINPUT24), .Z(new_n703));
  AOI21_X1  g278(.A(G29), .B1(new_n703), .B2(G34), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G34), .B2(new_n703), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT93), .ZN(new_n706));
  INV_X1    g281(.A(G160), .ZN(new_n707));
  INV_X1    g282(.A(G29), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n706), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(G2084), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  MUX2_X1   g286(.A(G5), .B(G301), .S(G16), .Z(new_n712));
  OAI21_X1  g287(.A(new_n711), .B1(G1961), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n708), .A2(G32), .ZN(new_n714));
  NAND3_X1  g289(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT26), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n634), .A2(G105), .ZN(new_n717));
  AOI211_X1 g292(.A(new_n716), .B(new_n717), .C1(G129), .C2(new_n625), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n623), .A2(G141), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT94), .Z(new_n720));
  NAND2_X1  g295(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n714), .B1(new_n722), .B2(new_n708), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT27), .B(G1996), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n713), .B1(new_n723), .B2(new_n725), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT97), .Z(new_n727));
  NOR2_X1   g302(.A1(new_n631), .A2(new_n708), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT96), .Z(new_n729));
  NOR2_X1   g304(.A1(G29), .A2(G33), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT90), .Z(new_n731));
  NAND2_X1  g306(.A1(new_n623), .A2(G139), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n475), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n733), .A2(new_n468), .ZN(new_n734));
  XOR2_X1   g309(.A(KEYINPUT91), .B(KEYINPUT25), .Z(new_n735));
  NAND3_X1  g310(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n732), .A2(new_n734), .A3(new_n737), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n731), .B1(new_n738), .B2(new_n708), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(G2072), .Z(new_n740));
  NOR2_X1   g315(.A1(new_n709), .A2(new_n710), .ZN(new_n741));
  INV_X1    g316(.A(G1966), .ZN(new_n742));
  INV_X1    g317(.A(G21), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n743), .A2(G16), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G286), .B2(G16), .ZN(new_n745));
  AOI22_X1  g320(.A1(new_n712), .A2(G1961), .B1(new_n742), .B2(new_n745), .ZN(new_n746));
  XOR2_X1   g321(.A(KEYINPUT31), .B(G11), .Z(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT95), .ZN(new_n748));
  INV_X1    g323(.A(G28), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n749), .A2(KEYINPUT30), .ZN(new_n750));
  AOI21_X1  g325(.A(G29), .B1(new_n749), .B2(KEYINPUT30), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n748), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n746), .B(new_n752), .C1(new_n742), .C2(new_n745), .ZN(new_n753));
  NOR4_X1   g328(.A1(new_n729), .A2(new_n740), .A3(new_n741), .A4(new_n753), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT85), .B(G16), .Z(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n756), .A2(G19), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(new_n551), .B2(new_n756), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT89), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(G1341), .Z(new_n760));
  NAND2_X1  g335(.A1(new_n708), .A2(G26), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT28), .ZN(new_n762));
  INV_X1    g337(.A(G128), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n468), .A2(G116), .ZN(new_n764));
  OAI21_X1  g339(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n765));
  OAI22_X1  g340(.A1(new_n486), .A2(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(G140), .B2(new_n623), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n762), .B1(new_n767), .B2(new_n708), .ZN(new_n768));
  INV_X1    g343(.A(G2067), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(new_n723), .B2(new_n725), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n708), .A2(G27), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G164), .B2(new_n708), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT98), .B(G2078), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NOR3_X1   g350(.A1(new_n760), .A2(new_n771), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n755), .A2(G20), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT99), .Z(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT23), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G16), .B2(G299), .ZN(new_n780));
  INV_X1    g355(.A(G1956), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(G4), .A2(G16), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n609), .B2(G16), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT88), .B(G1348), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(G29), .A2(G35), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G162), .B2(G29), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT29), .B(G2090), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NOR3_X1   g365(.A1(new_n782), .A2(new_n786), .A3(new_n790), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n727), .A2(new_n754), .A3(new_n776), .A4(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(G6), .A2(G16), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(new_n588), .B2(G16), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT32), .ZN(new_n795));
  INV_X1    g370(.A(G1981), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  MUX2_X1   g372(.A(G23), .B(G288), .S(G16), .Z(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT33), .B(G1976), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT86), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n798), .B(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n755), .A2(G22), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G166), .B2(new_n755), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n801), .B1(new_n803), .B2(G1971), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n803), .A2(G1971), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n797), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT87), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g383(.A1(new_n797), .A2(new_n804), .A3(KEYINPUT87), .A4(new_n805), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT34), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n808), .A2(KEYINPUT34), .A3(new_n809), .ZN(new_n813));
  NOR2_X1   g388(.A1(G25), .A2(G29), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n623), .A2(G131), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n625), .A2(G119), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n468), .A2(G107), .ZN(new_n817));
  OAI21_X1  g392(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n818));
  OAI211_X1 g393(.A(new_n815), .B(new_n816), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT84), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n819), .A2(new_n820), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n814), .B1(new_n824), .B2(G29), .ZN(new_n825));
  XOR2_X1   g400(.A(KEYINPUT35), .B(G1991), .Z(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n756), .A2(G24), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n828), .B1(new_n596), .B2(new_n756), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(G1986), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n812), .A2(new_n813), .A3(new_n827), .A4(new_n831), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n832), .A2(KEYINPUT36), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(KEYINPUT36), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n792), .B1(new_n833), .B2(new_n834), .ZN(G311));
  INV_X1    g410(.A(G311), .ZN(G150));
  NAND2_X1  g411(.A1(new_n609), .A2(G559), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT38), .ZN(new_n838));
  AOI22_X1  g413(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n839), .A2(new_n514), .ZN(new_n840));
  INV_X1    g415(.A(G93), .ZN(new_n841));
  INV_X1    g416(.A(G55), .ZN(new_n842));
  OAI22_X1  g417(.A1(new_n520), .A2(new_n841), .B1(new_n522), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n551), .B(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n838), .B(new_n846), .ZN(new_n847));
  OR2_X1    g422(.A1(new_n847), .A2(KEYINPUT39), .ZN(new_n848));
  INV_X1    g423(.A(G860), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(KEYINPUT39), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n844), .A2(new_n849), .ZN(new_n852));
  XNOR2_X1  g427(.A(KEYINPUT100), .B(KEYINPUT37), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n851), .A2(new_n854), .ZN(G145));
  XNOR2_X1  g430(.A(new_n631), .B(G160), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(G162), .ZN(new_n857));
  XNOR2_X1  g432(.A(KEYINPUT102), .B(KEYINPUT103), .ZN(new_n858));
  INV_X1    g433(.A(new_n738), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n718), .A2(new_n720), .A3(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n859), .B1(new_n718), .B2(new_n720), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n858), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n862), .ZN(new_n864));
  INV_X1    g439(.A(new_n858), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n864), .A2(new_n860), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n496), .A2(new_n497), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n868), .B1(new_n625), .B2(G126), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n506), .A2(KEYINPUT4), .ZN(new_n870));
  INV_X1    g445(.A(new_n504), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n767), .B(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n867), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n623), .A2(G142), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n625), .A2(G130), .ZN(new_n877));
  NOR3_X1   g452(.A1(new_n468), .A2(KEYINPUT101), .A3(G118), .ZN(new_n878));
  OAI21_X1  g453(.A(KEYINPUT101), .B1(new_n468), .B2(G118), .ZN(new_n879));
  OR2_X1    g454(.A1(G106), .A2(G2105), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n879), .A2(G2104), .A3(new_n880), .ZN(new_n881));
  OAI211_X1 g456(.A(new_n876), .B(new_n877), .C1(new_n878), .C2(new_n881), .ZN(new_n882));
  OR2_X1    g457(.A1(new_n636), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n636), .A2(new_n882), .ZN(new_n884));
  AND3_X1   g459(.A1(new_n823), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n823), .B1(new_n883), .B2(new_n884), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n874), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n863), .A2(new_n866), .A3(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n875), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(KEYINPUT104), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n887), .B1(new_n875), .B2(new_n889), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n857), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n875), .A2(new_n889), .ZN(new_n894));
  INV_X1    g469(.A(new_n887), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n857), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n896), .A2(KEYINPUT104), .A3(new_n897), .A4(new_n890), .ZN(new_n898));
  INV_X1    g473(.A(G37), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n893), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(KEYINPUT40), .ZN(G395));
  AOI21_X1  g476(.A(G305), .B1(new_n525), .B2(new_n532), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  AND2_X1   g478(.A1(new_n512), .A2(G60), .ZN(new_n904));
  OAI21_X1  g479(.A(G651), .B1(new_n904), .B2(new_n590), .ZN(new_n905));
  AOI22_X1  g480(.A1(new_n528), .A2(G85), .B1(new_n530), .B2(G47), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT106), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(KEYINPUT106), .B1(new_n592), .B2(new_n595), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(G288), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n525), .A2(new_n532), .A3(G305), .ZN(new_n912));
  INV_X1    g487(.A(G288), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n908), .A2(new_n909), .A3(new_n913), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n903), .A2(new_n911), .A3(new_n912), .A4(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT108), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n914), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n913), .B1(new_n908), .B2(new_n909), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n525), .A2(new_n532), .A3(G305), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n921), .A2(new_n902), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n920), .A2(new_n922), .A3(KEYINPUT108), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n917), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT107), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n925), .B1(new_n920), .B2(new_n922), .ZN(new_n926));
  OAI221_X1 g501(.A(KEYINPUT107), .B1(new_n921), .B2(new_n902), .C1(new_n918), .C2(new_n919), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n924), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT109), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n924), .A2(new_n928), .A3(KEYINPUT109), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(KEYINPUT42), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n609), .A2(G299), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT105), .ZN(new_n936));
  OAI211_X1 g511(.A(new_n572), .B(new_n564), .C1(new_n604), .C2(new_n608), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n609), .A2(KEYINPUT105), .A3(G299), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n938), .A2(KEYINPUT41), .A3(new_n939), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT41), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n935), .A2(new_n942), .A3(new_n937), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n846), .B(new_n618), .ZN(new_n945));
  MUX2_X1   g520(.A(new_n940), .B(new_n944), .S(new_n945), .Z(new_n946));
  INV_X1    g521(.A(KEYINPUT42), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n929), .A2(new_n947), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n934), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n946), .B1(new_n934), .B2(new_n948), .ZN(new_n950));
  OAI21_X1  g525(.A(G868), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n951), .B1(G868), .B2(new_n844), .ZN(G295));
  OAI21_X1  g527(.A(new_n951), .B1(G868), .B2(new_n844), .ZN(G331));
  INV_X1    g528(.A(KEYINPUT43), .ZN(new_n954));
  AND3_X1   g529(.A1(G171), .A2(KEYINPUT111), .A3(G286), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT111), .B1(G171), .B2(G286), .ZN(new_n956));
  OR2_X1    g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NOR3_X1   g532(.A1(G171), .A2(G286), .A3(KEYINPUT110), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(KEYINPUT110), .B1(G171), .B2(G286), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n551), .B(new_n844), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n957), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(new_n960), .ZN(new_n964));
  OAI22_X1  g539(.A1(new_n964), .A2(new_n958), .B1(new_n955), .B2(new_n956), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(new_n846), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n963), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT41), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(new_n940), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n935), .A2(new_n937), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n967), .A2(KEYINPUT41), .A3(new_n970), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n924), .A2(new_n928), .A3(KEYINPUT109), .ZN(new_n972));
  AOI21_X1  g547(.A(KEYINPUT109), .B1(new_n924), .B2(new_n928), .ZN(new_n973));
  OAI211_X1 g548(.A(new_n969), .B(new_n971), .C1(new_n972), .C2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n944), .A2(new_n967), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n940), .A2(new_n963), .A3(new_n966), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n977), .A2(new_n931), .A3(new_n932), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n974), .A2(new_n978), .A3(new_n899), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT112), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n974), .A2(new_n978), .A3(KEYINPUT112), .A4(new_n899), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n954), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  AND2_X1   g558(.A1(new_n978), .A2(new_n899), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n933), .A2(new_n976), .A3(new_n975), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT43), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(KEYINPUT44), .B1(new_n983), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT44), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n954), .B1(new_n984), .B2(new_n985), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n979), .A2(KEYINPUT43), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n988), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n987), .A2(new_n991), .ZN(G397));
  INV_X1    g567(.A(G1384), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n993), .B1(new_n498), .B2(new_n507), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT45), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n482), .B1(new_n481), .B2(new_n468), .ZN(new_n997));
  AOI211_X1 g572(.A(KEYINPUT69), .B(G2105), .C1(new_n464), .C2(new_n466), .ZN(new_n998));
  OAI21_X1  g573(.A(G101), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(G113), .A2(G2104), .ZN(new_n1000));
  INV_X1    g575(.A(G125), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n1000), .B1(new_n501), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(G2105), .ZN(new_n1003));
  AND2_X1   g578(.A1(new_n469), .A2(new_n472), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n1004), .A2(G137), .A3(new_n468), .A4(new_n467), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n999), .A2(G40), .A3(new_n1003), .A4(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n996), .A2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n767), .B(G2067), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n722), .A2(G1996), .ZN(new_n1009));
  INV_X1    g584(.A(G1996), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n721), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1008), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  XOR2_X1   g587(.A(new_n823), .B(new_n826), .Z(new_n1013));
  OR2_X1    g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G1986), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n596), .B(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1007), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT50), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1018), .B1(new_n873), .B2(new_n993), .ZN(new_n1019));
  INV_X1    g594(.A(G40), .ZN(new_n1020));
  NOR3_X1   g595(.A1(new_n477), .A2(new_n1020), .A3(new_n484), .ZN(new_n1021));
  NOR2_X1   g596(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1022), .B1(new_n498), .B2(new_n507), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n781), .B1(new_n1019), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT57), .ZN(new_n1026));
  AND3_X1   g601(.A1(new_n564), .A2(new_n1026), .A3(new_n572), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1026), .B1(new_n564), .B2(new_n572), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1006), .B1(new_n994), .B2(new_n995), .ZN(new_n1030));
  OAI211_X1 g605(.A(KEYINPUT45), .B(new_n993), .C1(new_n498), .C2(new_n507), .ZN(new_n1031));
  XNOR2_X1  g606(.A(KEYINPUT56), .B(G2072), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1025), .A2(new_n1029), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(new_n609), .ZN(new_n1035));
  OAI21_X1  g610(.A(KEYINPUT119), .B1(new_n1019), .B2(new_n1024), .ZN(new_n1036));
  INV_X1    g611(.A(G1348), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n994), .A2(KEYINPUT50), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT119), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1038), .A2(new_n1039), .A3(new_n1021), .A4(new_n1023), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1036), .A2(new_n1037), .A3(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n994), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1042), .A2(new_n769), .A3(new_n1021), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1035), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1029), .B1(new_n1025), .B2(new_n1033), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1034), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT120), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT120), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1048), .B(new_n1034), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT121), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1034), .B1(new_n1045), .B2(new_n1050), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1025), .A2(new_n1033), .A3(KEYINPUT121), .A4(new_n1029), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1051), .A2(KEYINPUT61), .A3(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT61), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1034), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1054), .B1(new_n1055), .B2(new_n1045), .ZN(new_n1056));
  XOR2_X1   g631(.A(KEYINPUT58), .B(G1341), .Z(new_n1057));
  OAI21_X1  g632(.A(new_n1057), .B1(new_n994), .B2(new_n1006), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n996), .A2(new_n1021), .A3(new_n1031), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1058), .B1(new_n1059), .B2(G1996), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(new_n551), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(KEYINPUT59), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT59), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1060), .A2(new_n1063), .A3(new_n551), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1053), .A2(new_n1056), .A3(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(KEYINPUT60), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1041), .A2(KEYINPUT60), .A3(new_n1043), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(new_n609), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1041), .A2(KEYINPUT60), .A3(new_n1035), .A4(new_n1043), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1067), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1047), .B(new_n1049), .C1(new_n1066), .C2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT54), .ZN(new_n1073));
  INV_X1    g648(.A(G1961), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1036), .A2(new_n1074), .A3(new_n1040), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(KEYINPUT123), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT123), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1036), .A2(new_n1077), .A3(new_n1074), .A4(new_n1040), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT53), .ZN(new_n1080));
  OR3_X1    g655(.A1(new_n1059), .A2(new_n1080), .A3(G2078), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1080), .B1(new_n1059), .B2(G2078), .ZN(new_n1082));
  AND2_X1   g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1079), .A2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1084), .A2(G171), .ZN(new_n1085));
  AOI21_X1  g660(.A(G301), .B1(new_n1083), .B2(new_n1075), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1073), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(G1976), .B1(new_n579), .B2(new_n580), .ZN(new_n1088));
  OR3_X1    g663(.A1(new_n1088), .A2(KEYINPUT114), .A3(KEYINPUT52), .ZN(new_n1089));
  OAI21_X1  g664(.A(KEYINPUT114), .B1(new_n1088), .B2(KEYINPUT52), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n913), .A2(G1976), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1092), .B(G8), .C1(new_n994), .C2(new_n1006), .ZN(new_n1093));
  OR2_X1    g668(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(KEYINPUT115), .A2(KEYINPUT49), .ZN(new_n1095));
  AOI22_X1  g670(.A1(new_n528), .A2(G86), .B1(new_n530), .B2(G48), .ZN(new_n1096));
  INV_X1    g671(.A(new_n587), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n796), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NOR3_X1   g673(.A1(new_n584), .A2(new_n587), .A3(G1981), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1095), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1096), .A2(new_n1097), .A3(new_n796), .ZN(new_n1101));
  OAI21_X1  g676(.A(G1981), .B1(new_n584), .B2(new_n587), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n1101), .B(new_n1102), .C1(KEYINPUT115), .C2(KEYINPUT49), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1100), .A2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(G8), .B1(new_n994), .B2(new_n1006), .ZN(new_n1105));
  OR2_X1    g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1093), .A2(KEYINPUT52), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1094), .A2(new_n1106), .A3(KEYINPUT117), .A4(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT117), .ZN(new_n1109));
  OAI22_X1  g684(.A1(new_n1091), .A2(new_n1093), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1110));
  AND2_X1   g685(.A1(new_n1093), .A2(KEYINPUT52), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1109), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1108), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT124), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n525), .A2(new_n532), .A3(G8), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT55), .ZN(new_n1116));
  XNOR2_X1  g691(.A(new_n1115), .B(new_n1116), .ZN(new_n1117));
  NOR3_X1   g692(.A1(new_n1019), .A2(new_n1024), .A3(G2090), .ZN(new_n1118));
  XOR2_X1   g693(.A(KEYINPUT113), .B(G1971), .Z(new_n1119));
  INV_X1    g694(.A(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1120), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1117), .B(G8), .C1(new_n1118), .C2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(G8), .B1(new_n1118), .B2(new_n1121), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1117), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1113), .A2(new_n1114), .A3(new_n1122), .A4(new_n1125), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1125), .A2(new_n1122), .A3(new_n1112), .A4(new_n1108), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(KEYINPUT124), .ZN(new_n1128));
  AND2_X1   g703(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1084), .A2(G171), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1081), .A2(new_n1075), .A3(G301), .A4(new_n1082), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1131), .A2(KEYINPUT54), .ZN(new_n1132));
  NOR2_X1   g707(.A1(KEYINPUT122), .A2(KEYINPUT51), .ZN(new_n1133));
  INV_X1    g708(.A(G8), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1059), .A2(new_n742), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1038), .A2(new_n710), .A3(new_n1021), .A4(new_n1023), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1134), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(G286), .A2(G8), .ZN(new_n1138));
  NAND2_X1  g713(.A1(KEYINPUT122), .A2(KEYINPUT51), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1133), .B1(new_n1137), .B2(new_n1140), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1019), .A2(new_n1024), .ZN(new_n1142));
  AOI22_X1  g717(.A1(new_n1142), .A2(new_n710), .B1(new_n1059), .B2(new_n742), .ZN(new_n1143));
  OR2_X1    g718(.A1(new_n1143), .A2(new_n1138), .ZN(new_n1144));
  AND2_X1   g719(.A1(new_n1141), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1140), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1133), .ZN(new_n1147));
  OAI211_X1 g722(.A(new_n1146), .B(new_n1147), .C1(new_n1143), .C2(new_n1134), .ZN(new_n1148));
  AOI22_X1  g723(.A1(new_n1130), .A2(new_n1132), .B1(new_n1145), .B2(new_n1148), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1072), .A2(new_n1087), .A3(new_n1129), .A4(new_n1149), .ZN(new_n1150));
  AND3_X1   g725(.A1(new_n1126), .A2(new_n1128), .A3(new_n1086), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1141), .A2(new_n1148), .A3(new_n1144), .ZN(new_n1152));
  OR2_X1    g727(.A1(new_n1152), .A2(KEYINPUT62), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT125), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1152), .A2(new_n1154), .A3(KEYINPUT62), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1152), .A2(KEYINPUT62), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(KEYINPUT125), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1151), .A2(new_n1153), .A3(new_n1155), .A4(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1150), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT118), .ZN(new_n1160));
  AOI211_X1 g735(.A(new_n1134), .B(G286), .C1(new_n1135), .C2(new_n1136), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT63), .ZN(new_n1162));
  NOR3_X1   g737(.A1(new_n1110), .A2(new_n1111), .A3(new_n1162), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1125), .A2(new_n1161), .A3(new_n1122), .A4(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1164), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1113), .A2(new_n1122), .A3(new_n1125), .A4(new_n1161), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1165), .B1(new_n1166), .B2(new_n1162), .ZN(new_n1167));
  NOR3_X1   g742(.A1(new_n1122), .A2(new_n1111), .A3(new_n1110), .ZN(new_n1168));
  INV_X1    g743(.A(G1976), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1106), .A2(new_n1169), .A3(new_n913), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n1099), .B(KEYINPUT116), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1105), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1168), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1160), .B1(new_n1167), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1161), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1162), .B1(new_n1127), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1177), .A2(new_n1164), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1178), .A2(KEYINPUT118), .A3(new_n1173), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1175), .A2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1017), .B1(new_n1159), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1182));
  OR2_X1    g757(.A1(new_n1182), .A2(KEYINPUT46), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1182), .A2(KEYINPUT46), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n722), .A2(new_n1008), .ZN(new_n1185));
  AOI22_X1  g760(.A1(new_n1183), .A2(new_n1184), .B1(new_n1185), .B2(new_n1007), .ZN(new_n1186));
  XNOR2_X1  g761(.A(new_n1186), .B(KEYINPUT47), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1014), .A2(new_n1007), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1007), .A2(new_n1015), .A3(new_n596), .ZN(new_n1189));
  XOR2_X1   g764(.A(new_n1189), .B(KEYINPUT127), .Z(new_n1190));
  XOR2_X1   g765(.A(KEYINPUT126), .B(KEYINPUT48), .Z(new_n1191));
  OR2_X1    g766(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1193));
  AND3_X1   g768(.A1(new_n1188), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n767), .A2(new_n769), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n824), .A2(new_n826), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1195), .B1(new_n1012), .B2(new_n1196), .ZN(new_n1197));
  AOI211_X1 g772(.A(new_n1187), .B(new_n1194), .C1(new_n1007), .C2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1181), .A2(new_n1198), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g774(.A(new_n461), .B1(new_n654), .B2(new_n655), .ZN(new_n1201));
  OR2_X1    g775(.A1(G227), .A2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g776(.A(new_n1202), .B1(new_n700), .B2(new_n701), .ZN(new_n1203));
  OAI211_X1 g777(.A(new_n1203), .B(new_n900), .C1(new_n989), .C2(new_n990), .ZN(G225));
  INV_X1    g778(.A(G225), .ZN(G308));
endmodule


