//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 1 0 1 0 1 0 1 0 1 0 1 0 0 1 1 0 0 1 1 0 0 0 1 1 1 0 0 1 1 0 0 1 1 1 1 1 0 1 1 1 1 0 1 1 0 0 0 0 1 0 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n748, new_n749, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n816, new_n817, new_n818, new_n820, new_n821,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n918, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n991, new_n992, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1033, new_n1034, new_n1035;
  INV_X1    g000(.A(KEYINPUT91), .ZN(new_n202));
  XNOR2_X1  g001(.A(G127gat), .B(G134gat), .ZN(new_n203));
  INV_X1    g002(.A(G113gat), .ZN(new_n204));
  INV_X1    g003(.A(G120gat), .ZN(new_n205));
  AOI21_X1  g004(.A(KEYINPUT1), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  AND2_X1   g005(.A1(new_n203), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(KEYINPUT69), .B(G120gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G113gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n206), .B1(new_n204), .B2(new_n205), .ZN(new_n210));
  INV_X1    g009(.A(new_n203), .ZN(new_n211));
  AOI22_X1  g010(.A1(new_n207), .A2(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G183gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT27), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT27), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G183gat), .ZN(new_n216));
  INV_X1    g015(.A(G190gat), .ZN(new_n217));
  NAND4_X1  g016(.A1(new_n214), .A2(new_n216), .A3(KEYINPUT28), .A4(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT67), .ZN(new_n219));
  XNOR2_X1  g018(.A(KEYINPUT27), .B(G183gat), .ZN(new_n220));
  AOI21_X1  g019(.A(KEYINPUT28), .B1(new_n220), .B2(new_n217), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n214), .A2(new_n216), .A3(new_n217), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT67), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT28), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(G183gat), .A2(G190gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(G169gat), .A2(G176gat), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT26), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(G169gat), .ZN(new_n232));
  INV_X1    g031(.A(G176gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n231), .A2(KEYINPUT68), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT68), .ZN(new_n236));
  AOI21_X1  g035(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n237));
  NOR2_X1   g036(.A1(G169gat), .A2(G176gat), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n236), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n230), .ZN(new_n240));
  AND3_X1   g039(.A1(new_n235), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  NOR3_X1   g040(.A1(new_n222), .A2(new_n228), .A3(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT23), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n243), .B1(G169gat), .B2(G176gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(new_n229), .ZN(new_n245));
  NOR3_X1   g044(.A1(new_n243), .A2(G169gat), .A3(G176gat), .ZN(new_n246));
  OAI21_X1  g045(.A(KEYINPUT64), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n238), .A2(KEYINPUT23), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT25), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(KEYINPUT64), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n248), .A2(new_n229), .A3(new_n244), .A4(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n252));
  NOR2_X1   g051(.A1(G183gat), .A2(G190gat), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n247), .A2(new_n251), .A3(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n248), .A2(new_n229), .A3(new_n244), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT65), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT24), .ZN(new_n260));
  AND3_X1   g059(.A1(new_n227), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n259), .B1(new_n227), .B2(new_n260), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT66), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n264), .A2(new_n213), .A3(new_n217), .ZN(new_n265));
  OAI21_X1  g064(.A(KEYINPUT66), .B1(G183gat), .B2(G190gat), .ZN(new_n266));
  AND3_X1   g065(.A1(new_n265), .A2(new_n255), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n258), .B1(new_n263), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n257), .B1(new_n268), .B2(new_n249), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n212), .B1(new_n242), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(G227gat), .ZN(new_n271));
  INV_X1    g070(.A(G233gat), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n245), .A2(new_n246), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n227), .A2(new_n260), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(KEYINPUT65), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n252), .A2(new_n259), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n265), .A2(new_n255), .A3(new_n266), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n274), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  AOI22_X1  g079(.A1(new_n258), .A2(KEYINPUT64), .B1(new_n255), .B2(new_n254), .ZN(new_n281));
  AOI22_X1  g080(.A1(new_n280), .A2(KEYINPUT25), .B1(new_n281), .B2(new_n251), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n209), .A2(new_n206), .A3(new_n203), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n210), .A2(new_n211), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n223), .A2(new_n225), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n286), .A2(KEYINPUT67), .A3(new_n218), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n235), .A2(new_n239), .A3(new_n240), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n287), .A2(new_n288), .A3(new_n227), .A4(new_n226), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n282), .A2(new_n285), .A3(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n270), .A2(new_n273), .A3(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT33), .ZN(new_n292));
  XNOR2_X1  g091(.A(G15gat), .B(G43gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(G71gat), .B(G99gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n293), .B(new_n294), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n291), .B(KEYINPUT32), .C1(new_n292), .C2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n295), .B1(new_n291), .B2(new_n292), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT70), .ZN(new_n299));
  AND3_X1   g098(.A1(new_n291), .A2(new_n299), .A3(KEYINPUT32), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n299), .B1(new_n291), .B2(KEYINPUT32), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n298), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT71), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OAI211_X1 g103(.A(KEYINPUT71), .B(new_n298), .C1(new_n300), .C2(new_n301), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n297), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n270), .A2(new_n290), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n307), .B1(new_n271), .B2(new_n272), .ZN(new_n308));
  AND3_X1   g107(.A1(new_n308), .A2(KEYINPUT72), .A3(KEYINPUT34), .ZN(new_n309));
  AOI21_X1  g108(.A(KEYINPUT34), .B1(new_n308), .B2(KEYINPUT72), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(KEYINPUT36), .B1(new_n306), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n291), .A2(KEYINPUT32), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT70), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n291), .A2(new_n299), .A3(KEYINPUT32), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(KEYINPUT71), .B1(new_n316), .B2(new_n298), .ZN(new_n317));
  INV_X1    g116(.A(new_n305), .ZN(new_n318));
  OAI211_X1 g117(.A(new_n296), .B(new_n311), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT73), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n306), .A2(KEYINPUT73), .A3(new_n311), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n312), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT74), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n324), .B1(new_n306), .B2(new_n311), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n296), .B1(new_n317), .B2(new_n318), .ZN(new_n326));
  INV_X1    g125(.A(new_n311), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n326), .A2(new_n327), .A3(KEYINPUT74), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n319), .A2(new_n320), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT73), .B1(new_n306), .B2(new_n311), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n325), .B(new_n328), .C1(new_n329), .C2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT36), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n323), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(G225gat), .A2(G233gat), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(G155gat), .A2(G162gat), .ZN(new_n336));
  INV_X1    g135(.A(G155gat), .ZN(new_n337));
  INV_X1    g136(.A(G162gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  OR2_X1    g138(.A1(G141gat), .A2(G148gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(G141gat), .A2(G148gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n336), .B(new_n339), .C1(new_n342), .C2(KEYINPUT2), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT80), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n340), .A2(new_n344), .A3(new_n341), .ZN(new_n345));
  AND2_X1   g144(.A1(G141gat), .A2(G148gat), .ZN(new_n346));
  NOR2_X1   g145(.A1(G141gat), .A2(G148gat), .ZN(new_n347));
  OAI21_X1  g146(.A(KEYINPUT80), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n339), .A2(new_n336), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n345), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n336), .A2(KEYINPUT81), .A3(KEYINPUT2), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT81), .B1(new_n336), .B2(KEYINPUT2), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n343), .B1(new_n350), .B2(new_n354), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n355), .A2(new_n285), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n336), .A2(KEYINPUT2), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT81), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(new_n351), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n360), .A2(new_n349), .A3(new_n345), .A4(new_n348), .ZN(new_n361));
  AOI22_X1  g160(.A1(new_n361), .A2(new_n343), .B1(new_n283), .B2(new_n284), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n335), .B1(new_n356), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT5), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n355), .A2(KEYINPUT3), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT3), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n361), .A2(new_n366), .A3(new_n343), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n365), .A2(new_n367), .A3(new_n285), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT4), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n369), .B1(new_n355), .B2(new_n285), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n212), .A2(KEYINPUT4), .A3(new_n343), .A4(new_n361), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n368), .A2(new_n334), .A3(new_n370), .A4(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n364), .A2(new_n372), .ZN(new_n373));
  AND2_X1   g172(.A1(new_n370), .A2(new_n371), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n374), .A2(KEYINPUT5), .A3(new_n334), .A4(new_n368), .ZN(new_n375));
  XNOR2_X1  g174(.A(G1gat), .B(G29gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n376), .B(KEYINPUT0), .ZN(new_n377));
  XNOR2_X1  g176(.A(G57gat), .B(G85gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n377), .B(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n379), .B(KEYINPUT84), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n373), .A2(new_n375), .A3(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT39), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n368), .A2(new_n370), .A3(new_n371), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT85), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n384), .A2(new_n385), .A3(new_n335), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n385), .B1(new_n384), .B2(new_n335), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n383), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n384), .A2(new_n335), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(KEYINPUT85), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n356), .A2(new_n362), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n383), .B1(new_n392), .B2(new_n334), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n391), .A2(new_n386), .A3(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n380), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n389), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT86), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n382), .B1(new_n398), .B2(KEYINPUT40), .ZN(new_n399));
  XNOR2_X1  g198(.A(G8gat), .B(G36gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(G64gat), .B(G92gat), .ZN(new_n401));
  XOR2_X1   g200(.A(new_n400), .B(new_n401), .Z(new_n402));
  NAND2_X1  g201(.A1(G211gat), .A2(G218gat), .ZN(new_n403));
  INV_X1    g202(.A(G211gat), .ZN(new_n404));
  INV_X1    g203(.A(G218gat), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AND2_X1   g205(.A1(G197gat), .A2(G204gat), .ZN(new_n407));
  NOR2_X1   g206(.A1(G197gat), .A2(G204gat), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT22), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n403), .B(new_n406), .C1(new_n409), .C2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n406), .A2(new_n403), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n403), .A2(new_n410), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n412), .B(new_n413), .C1(new_n408), .C2(new_n407), .ZN(new_n414));
  AND3_X1   g213(.A1(new_n411), .A2(new_n414), .A3(KEYINPUT75), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT75), .B1(new_n411), .B2(new_n414), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n280), .A2(KEYINPUT25), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n289), .A2(new_n419), .A3(new_n257), .ZN(new_n420));
  NAND2_X1  g219(.A1(G226gat), .A2(G233gat), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(KEYINPUT76), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n422), .B1(new_n242), .B2(new_n269), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT29), .B1(new_n282), .B2(new_n289), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n424), .B1(new_n425), .B2(new_n422), .ZN(new_n426));
  AOI211_X1 g225(.A(new_n418), .B(new_n423), .C1(new_n426), .C2(KEYINPUT76), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n421), .B1(new_n282), .B2(new_n289), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT29), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n429), .B1(new_n242), .B2(new_n269), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n428), .B1(new_n430), .B2(new_n421), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n431), .A2(new_n417), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n402), .B1(new_n427), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT30), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n423), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT76), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n417), .B(new_n436), .C1(new_n431), .C2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n426), .A2(new_n418), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n402), .B(KEYINPUT77), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT78), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  OAI211_X1 g242(.A(KEYINPUT30), .B(new_n402), .C1(new_n427), .C2(new_n432), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n438), .A2(KEYINPUT78), .A3(new_n439), .A4(new_n440), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n435), .A2(new_n443), .A3(new_n444), .A4(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT40), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n396), .A2(new_n397), .A3(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n399), .A2(new_n446), .A3(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(G78gat), .ZN(new_n450));
  INV_X1    g249(.A(G22gat), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n367), .A2(new_n429), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(new_n417), .ZN(new_n453));
  AND2_X1   g252(.A1(G228gat), .A2(G233gat), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT29), .B1(new_n411), .B2(new_n414), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(new_n355), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n453), .A2(new_n365), .A3(new_n454), .A4(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT83), .ZN(new_n458));
  AND2_X1   g257(.A1(new_n411), .A2(new_n414), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n458), .B1(new_n459), .B2(KEYINPUT29), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n455), .A2(KEYINPUT83), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(new_n366), .A3(new_n461), .ZN(new_n462));
  AOI22_X1  g261(.A1(new_n462), .A2(new_n355), .B1(new_n417), .B2(new_n452), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n451), .B(new_n457), .C1(new_n463), .C2(new_n454), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n366), .B1(new_n455), .B2(KEYINPUT83), .ZN(new_n465));
  AOI211_X1 g264(.A(new_n458), .B(KEYINPUT29), .C1(new_n411), .C2(new_n414), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n355), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n454), .B1(new_n467), .B2(new_n453), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n456), .A2(new_n365), .A3(new_n454), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n469), .B1(new_n417), .B2(new_n452), .ZN(new_n470));
  OAI21_X1  g269(.A(G22gat), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n450), .B1(new_n464), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n464), .A2(new_n471), .A3(new_n450), .ZN(new_n474));
  XNOR2_X1  g273(.A(KEYINPUT31), .B(G50gat), .ZN(new_n475));
  INV_X1    g274(.A(G106gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n475), .B(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n473), .A2(new_n474), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n477), .ZN(new_n479));
  AND3_X1   g278(.A1(new_n464), .A2(new_n471), .A3(new_n450), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n479), .B1(new_n480), .B2(new_n472), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT89), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n423), .B1(new_n426), .B2(KEYINPUT76), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n432), .B1(new_n417), .B2(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(KEYINPUT88), .B(KEYINPUT37), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n484), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n438), .A2(new_n439), .ZN(new_n489));
  INV_X1    g288(.A(new_n487), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n489), .A2(KEYINPUT89), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT38), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n440), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT37), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n495), .B1(new_n431), .B2(new_n417), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n496), .B1(new_n485), .B2(new_n417), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT87), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT87), .ZN(new_n499));
  OAI211_X1 g298(.A(new_n496), .B(new_n499), .C1(new_n485), .C2(new_n417), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n494), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n492), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n373), .A2(new_n375), .ZN(new_n503));
  INV_X1    g302(.A(new_n379), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT6), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n505), .A2(new_n506), .A3(new_n381), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n373), .A2(new_n375), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT90), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n508), .A2(new_n509), .A3(KEYINPUT6), .A4(new_n379), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n373), .A2(new_n375), .A3(KEYINPUT6), .A4(new_n379), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT90), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n507), .A2(new_n433), .A3(new_n510), .A4(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n502), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n402), .B1(new_n486), .B2(KEYINPUT37), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n493), .B1(new_n492), .B2(new_n516), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n449), .B(new_n483), .C1(new_n515), .C2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT79), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n443), .A2(new_n444), .A3(KEYINPUT79), .A4(new_n445), .ZN(new_n522));
  OAI21_X1  g321(.A(KEYINPUT82), .B1(new_n503), .B2(new_n504), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT82), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n373), .A2(new_n375), .A3(new_n524), .A4(new_n379), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n523), .A2(new_n506), .A3(new_n525), .A4(new_n505), .ZN(new_n526));
  AOI22_X1  g325(.A1(new_n526), .A2(new_n511), .B1(new_n434), .B2(new_n433), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n521), .A2(new_n522), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(new_n482), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n518), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n333), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n331), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n507), .A2(new_n510), .A3(new_n512), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT35), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n478), .A2(new_n481), .A3(new_n533), .A4(new_n534), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n535), .A2(new_n446), .ZN(new_n536));
  AND3_X1   g335(.A1(new_n521), .A2(new_n522), .A3(new_n527), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n321), .A2(new_n322), .ZN(new_n538));
  OAI211_X1 g337(.A(new_n478), .B(new_n481), .C1(new_n306), .C2(new_n311), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n537), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  AOI22_X1  g340(.A1(new_n532), .A2(new_n536), .B1(new_n541), .B2(KEYINPUT35), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n202), .B1(new_n531), .B2(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n513), .B1(new_n492), .B2(new_n501), .ZN(new_n544));
  AOI21_X1  g343(.A(KEYINPUT89), .B1(new_n489), .B2(new_n490), .ZN(new_n545));
  AOI211_X1 g344(.A(new_n484), .B(new_n487), .C1(new_n438), .C2(new_n439), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n516), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT38), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n482), .B1(new_n544), .B2(new_n548), .ZN(new_n549));
  AOI22_X1  g348(.A1(new_n549), .A2(new_n449), .B1(new_n528), .B2(new_n482), .ZN(new_n550));
  AOI21_X1  g349(.A(KEYINPUT74), .B1(new_n326), .B2(new_n327), .ZN(new_n551));
  NOR3_X1   g350(.A1(new_n306), .A2(new_n324), .A3(new_n311), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(KEYINPUT36), .B1(new_n553), .B2(new_n538), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n550), .B1(new_n554), .B2(new_n323), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n541), .A2(KEYINPUT35), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n553), .A2(new_n538), .A3(new_n536), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n555), .A2(new_n558), .A3(KEYINPUT91), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(G8gat), .ZN(new_n561));
  XOR2_X1   g360(.A(G15gat), .B(G22gat), .Z(new_n562));
  INV_X1    g361(.A(G1gat), .ZN(new_n563));
  AOI21_X1  g362(.A(KEYINPUT95), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G15gat), .B(G22gat), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT16), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n565), .B1(new_n566), .B2(G1gat), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n561), .B1(new_n564), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n564), .A2(new_n561), .A3(new_n567), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(G29gat), .A2(G36gat), .ZN(new_n572));
  OAI21_X1  g371(.A(KEYINPUT93), .B1(G29gat), .B2(G36gat), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n572), .B1(new_n573), .B2(KEYINPUT14), .ZN(new_n574));
  INV_X1    g373(.A(new_n573), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT14), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT93), .ZN(new_n578));
  INV_X1    g377(.A(G29gat), .ZN(new_n579));
  INV_X1    g378(.A(G36gat), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n574), .B1(new_n577), .B2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(G43gat), .ZN(new_n583));
  INV_X1    g382(.A(G50gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT15), .ZN(new_n586));
  NAND2_X1  g385(.A1(G43gat), .A2(G50gat), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT94), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n585), .A2(new_n587), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n590), .A2(new_n586), .ZN(new_n591));
  OAI211_X1 g390(.A(new_n582), .B(new_n588), .C1(new_n589), .C2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n591), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n581), .A2(KEYINPUT14), .A3(new_n573), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n575), .A2(new_n576), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n594), .A2(new_n595), .A3(new_n589), .A4(new_n572), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n594), .A2(new_n595), .A3(new_n572), .A4(new_n588), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n593), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n571), .A2(new_n592), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(G229gat), .A2(G233gat), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT17), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n592), .A2(new_n598), .A3(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n570), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n603), .A2(new_n568), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n601), .B1(new_n592), .B2(new_n598), .ZN(new_n606));
  OAI211_X1 g405(.A(new_n599), .B(new_n600), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT18), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n606), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n610), .A2(new_n604), .A3(new_n602), .ZN(new_n611));
  NAND4_X1  g410(.A1(new_n611), .A2(KEYINPUT18), .A3(new_n600), .A4(new_n599), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n592), .A2(new_n598), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n604), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT96), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n599), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  XOR2_X1   g415(.A(new_n600), .B(KEYINPUT13), .Z(new_n617));
  NAND3_X1  g416(.A1(new_n604), .A2(new_n613), .A3(KEYINPUT96), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n609), .A2(new_n612), .A3(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G113gat), .B(G141gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(G197gat), .ZN(new_n622));
  XOR2_X1   g421(.A(KEYINPUT11), .B(G169gat), .Z(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT92), .B(KEYINPUT12), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n624), .B(new_n625), .Z(new_n626));
  NAND2_X1  g425(.A1(new_n620), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n626), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n628), .A2(new_n609), .A3(new_n612), .A4(new_n619), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(G232gat), .A2(G233gat), .ZN(new_n631));
  XOR2_X1   g430(.A(new_n631), .B(KEYINPUT100), .Z(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n633), .A2(KEYINPUT41), .ZN(new_n634));
  XNOR2_X1  g433(.A(G134gat), .B(G162gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT102), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(G92gat), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n639), .A2(KEYINPUT7), .A3(G85gat), .ZN(new_n640));
  NAND2_X1  g439(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(G92gat), .ZN(new_n642));
  NOR2_X1   g441(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n640), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(G99gat), .B(G106gat), .ZN(new_n645));
  NAND2_X1  g444(.A1(G99gat), .A2(G106gat), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT101), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(KEYINPUT101), .A2(G99gat), .A3(G106gat), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n648), .A2(KEYINPUT8), .A3(new_n649), .ZN(new_n650));
  AND3_X1   g449(.A1(new_n644), .A2(new_n645), .A3(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n645), .B1(new_n644), .B2(new_n650), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n613), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n653), .B1(KEYINPUT41), .B2(new_n633), .ZN(new_n654));
  OAI211_X1 g453(.A(new_n610), .B(new_n602), .C1(new_n651), .C2(new_n652), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g455(.A(G190gat), .B(G218gat), .Z(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n657), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n654), .A2(new_n659), .A3(new_n655), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n638), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  AND2_X1   g460(.A1(new_n658), .A2(new_n660), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n636), .B(new_n637), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(G120gat), .B(G148gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(G176gat), .B(G204gat), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n666), .B(new_n667), .Z(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n644), .A2(new_n650), .ZN(new_n670));
  INV_X1    g469(.A(new_n645), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n644), .A2(new_n645), .A3(new_n650), .ZN(new_n673));
  XNOR2_X1  g472(.A(G71gat), .B(G78gat), .ZN(new_n674));
  NAND2_X1  g473(.A1(G71gat), .A2(G78gat), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT9), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  OR2_X1    g476(.A1(G57gat), .A2(G64gat), .ZN(new_n678));
  NAND2_X1  g477(.A1(G57gat), .A2(G64gat), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n674), .B1(new_n680), .B2(KEYINPUT97), .ZN(new_n681));
  AND3_X1   g480(.A1(new_n680), .A2(KEYINPUT97), .A3(new_n674), .ZN(new_n682));
  OAI211_X1 g481(.A(new_n672), .B(new_n673), .C1(new_n681), .C2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n680), .A2(KEYINPUT97), .ZN(new_n684));
  INV_X1    g483(.A(new_n674), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n680), .A2(KEYINPUT97), .A3(new_n674), .ZN(new_n687));
  OAI211_X1 g486(.A(new_n686), .B(new_n687), .C1(new_n651), .C2(new_n652), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT10), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n683), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(KEYINPUT103), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT103), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n683), .A2(new_n688), .A3(new_n692), .A4(new_n689), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(KEYINPUT104), .B1(new_n683), .B2(new_n689), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n651), .A2(new_n652), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n686), .A2(new_n687), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT104), .ZN(new_n698));
  NAND4_X1  g497(.A1(new_n696), .A2(new_n697), .A3(new_n698), .A4(KEYINPUT10), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n694), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT105), .ZN(new_n702));
  NAND2_X1  g501(.A1(G230gat), .A2(G233gat), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  AOI22_X1  g503(.A1(new_n691), .A2(new_n693), .B1(new_n695), .B2(new_n699), .ZN(new_n705));
  INV_X1    g504(.A(new_n703), .ZN(new_n706));
  OAI21_X1  g505(.A(KEYINPUT105), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n683), .A2(new_n688), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(new_n706), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n669), .B1(new_n708), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n701), .A2(new_n703), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n711), .A2(new_n669), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n697), .A2(KEYINPUT21), .ZN(new_n717));
  XNOR2_X1  g516(.A(KEYINPUT99), .B(KEYINPUT19), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n571), .B1(KEYINPUT21), .B2(new_n697), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n719), .B(new_n720), .ZN(new_n721));
  XNOR2_X1  g520(.A(G127gat), .B(G155gat), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(KEYINPUT20), .ZN(new_n723));
  NAND2_X1  g522(.A1(G231gat), .A2(G233gat), .ZN(new_n724));
  XOR2_X1   g523(.A(new_n724), .B(KEYINPUT98), .Z(new_n725));
  XNOR2_X1  g524(.A(new_n723), .B(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(G183gat), .B(G211gat), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n721), .B(new_n728), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n665), .A2(new_n716), .A3(new_n729), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n560), .A2(new_n630), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n526), .A2(new_n511), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(new_n563), .ZN(G1324gat));
  INV_X1    g533(.A(new_n446), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n731), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n736), .A2(new_n561), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n566), .A2(new_n561), .ZN(new_n738));
  NOR2_X1   g537(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n739));
  NOR4_X1   g538(.A1(new_n731), .A2(new_n735), .A3(new_n738), .A4(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(KEYINPUT42), .B1(new_n737), .B2(new_n740), .ZN(new_n741));
  OR2_X1    g540(.A1(new_n740), .A2(KEYINPUT42), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(G1325gat));
  INV_X1    g542(.A(new_n333), .ZN(new_n744));
  OAI21_X1  g543(.A(G15gat), .B1(new_n731), .B2(new_n744), .ZN(new_n745));
  OR2_X1    g544(.A1(new_n331), .A2(G15gat), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n745), .B1(new_n731), .B2(new_n746), .ZN(G1326gat));
  NOR2_X1   g546(.A1(new_n731), .A2(new_n483), .ZN(new_n748));
  XOR2_X1   g547(.A(KEYINPUT43), .B(G22gat), .Z(new_n749));
  XNOR2_X1  g548(.A(new_n748), .B(new_n749), .ZN(G1327gat));
  INV_X1    g549(.A(new_n716), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(new_n729), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n752), .A2(new_n664), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n560), .A2(new_n630), .A3(new_n753), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n754), .A2(G29gat), .A3(new_n732), .ZN(new_n755));
  OR2_X1    g554(.A1(new_n755), .A2(KEYINPUT45), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(KEYINPUT45), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n539), .B1(new_n321), .B2(new_n322), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n534), .B1(new_n758), .B2(new_n537), .ZN(new_n759));
  AND4_X1   g558(.A1(new_n538), .A2(new_n536), .A3(new_n325), .A4(new_n328), .ZN(new_n760));
  OAI22_X1  g559(.A1(new_n333), .A2(new_n530), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  AOI21_X1  g560(.A(KEYINPUT44), .B1(new_n761), .B2(new_n665), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT44), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n664), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n762), .B1(new_n560), .B2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(new_n732), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT106), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n630), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n627), .A2(KEYINPUT106), .A3(new_n629), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n752), .A2(new_n771), .ZN(new_n772));
  AND3_X1   g571(.A1(new_n765), .A2(new_n766), .A3(new_n772), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n756), .B(new_n757), .C1(new_n773), .C2(new_n579), .ZN(G1328gat));
  NAND3_X1  g573(.A1(new_n765), .A2(new_n446), .A3(new_n772), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT107), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n765), .A2(KEYINPUT107), .A3(new_n446), .A4(new_n772), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n777), .A2(G36gat), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n446), .A2(new_n580), .ZN(new_n780));
  OAI21_X1  g579(.A(KEYINPUT46), .B1(new_n754), .B2(new_n780), .ZN(new_n781));
  OR3_X1    g580(.A1(new_n754), .A2(KEYINPUT46), .A3(new_n780), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n779), .A2(new_n781), .A3(new_n782), .ZN(G1329gat));
  NAND4_X1  g582(.A1(new_n765), .A2(G43gat), .A3(new_n333), .A4(new_n772), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n754), .A2(new_n331), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n784), .B1(new_n785), .B2(G43gat), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(KEYINPUT47), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT47), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n784), .B(new_n788), .C1(new_n785), .C2(G43gat), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n787), .A2(new_n789), .ZN(G1330gat));
  AND3_X1   g589(.A1(new_n555), .A2(new_n558), .A3(KEYINPUT91), .ZN(new_n791));
  AOI21_X1  g590(.A(KEYINPUT91), .B1(new_n555), .B2(new_n558), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n764), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n531), .A2(new_n542), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n763), .B1(new_n794), .B2(new_n664), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n793), .A2(new_n482), .A3(new_n795), .A4(new_n772), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(G50gat), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n482), .A2(new_n584), .ZN(new_n798));
  OR2_X1    g597(.A1(new_n754), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT48), .ZN(new_n800));
  AND3_X1   g599(.A1(new_n797), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n800), .B1(new_n797), .B2(new_n799), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n801), .A2(new_n802), .ZN(G1331gat));
  INV_X1    g602(.A(new_n729), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n771), .A2(new_n804), .A3(new_n664), .A4(new_n716), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n794), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n766), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(G57gat), .ZN(G1332gat));
  OR3_X1    g607(.A1(new_n794), .A2(KEYINPUT108), .A3(new_n805), .ZN(new_n809));
  OAI21_X1  g608(.A(KEYINPUT108), .B1(new_n794), .B2(new_n805), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n446), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n812), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n813));
  XOR2_X1   g612(.A(KEYINPUT49), .B(G64gat), .Z(new_n814));
  OAI21_X1  g613(.A(new_n813), .B1(new_n812), .B2(new_n814), .ZN(G1333gat));
  NAND4_X1  g614(.A1(new_n809), .A2(G71gat), .A3(new_n333), .A4(new_n810), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n794), .A2(new_n331), .A3(new_n805), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n816), .B1(G71gat), .B2(new_n817), .ZN(new_n818));
  XNOR2_X1  g617(.A(new_n818), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g618(.A1(new_n811), .A2(new_n482), .ZN(new_n820));
  XNOR2_X1  g619(.A(KEYINPUT109), .B(G78gat), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n820), .B(new_n821), .ZN(G1335gat));
  INV_X1    g621(.A(new_n765), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n770), .A2(new_n804), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n825), .A2(new_n751), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n823), .A2(new_n732), .A3(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(G85gat), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n761), .A2(new_n665), .A3(new_n824), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT51), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n830), .B(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n716), .A2(new_n766), .A3(new_n829), .ZN(new_n834));
  OAI22_X1  g633(.A1(new_n828), .A2(new_n829), .B1(new_n833), .B2(new_n834), .ZN(G1336gat));
  NAND3_X1  g634(.A1(new_n716), .A2(new_n639), .A3(new_n446), .ZN(new_n836));
  XOR2_X1   g635(.A(new_n836), .B(KEYINPUT110), .Z(new_n837));
  NAND2_X1  g636(.A1(new_n832), .A2(new_n837), .ZN(new_n838));
  AND4_X1   g637(.A1(new_n446), .A2(new_n793), .A3(new_n795), .A4(new_n826), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n838), .B1(new_n839), .B2(new_n639), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(KEYINPUT52), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT52), .ZN(new_n842));
  OAI211_X1 g641(.A(new_n838), .B(new_n842), .C1(new_n839), .C2(new_n639), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n841), .A2(new_n843), .ZN(G1337gat));
  NOR3_X1   g643(.A1(new_n823), .A2(new_n744), .A3(new_n827), .ZN(new_n845));
  INV_X1    g644(.A(G99gat), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n532), .A2(new_n846), .A3(new_n716), .ZN(new_n847));
  OAI22_X1  g646(.A1(new_n845), .A2(new_n846), .B1(new_n833), .B2(new_n847), .ZN(G1338gat));
  NAND4_X1  g647(.A1(new_n793), .A2(new_n482), .A3(new_n795), .A4(new_n826), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT112), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n765), .A2(KEYINPUT112), .A3(new_n482), .A4(new_n826), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n851), .A2(new_n852), .A3(G106gat), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n716), .A2(new_n482), .A3(new_n476), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n854), .B(KEYINPUT111), .ZN(new_n855));
  AOI21_X1  g654(.A(KEYINPUT53), .B1(new_n832), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n849), .A2(G106gat), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n832), .A2(new_n855), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(KEYINPUT53), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n857), .A2(new_n861), .ZN(G1339gat));
  INV_X1    g661(.A(KEYINPUT54), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n704), .A2(new_n707), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n705), .A2(new_n706), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n713), .A2(KEYINPUT54), .A3(new_n865), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n864), .A2(new_n866), .A3(KEYINPUT55), .A4(new_n669), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT114), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT55), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n863), .B1(new_n701), .B2(new_n703), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n870), .B1(new_n871), .B2(new_n865), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n872), .A2(KEYINPUT114), .A3(new_n669), .A4(new_n864), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n864), .A2(new_n669), .A3(new_n866), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n870), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n874), .A2(new_n715), .A3(new_n770), .A4(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT115), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n617), .B1(new_n616), .B2(new_n618), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n600), .B1(new_n611), .B2(new_n599), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n624), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n629), .A2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n716), .A2(new_n883), .ZN(new_n884));
  AND3_X1   g683(.A1(new_n877), .A2(new_n878), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n878), .B1(new_n877), .B2(new_n884), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n885), .A2(new_n886), .A3(new_n665), .ZN(new_n887));
  AOI22_X1  g686(.A1(new_n869), .A2(new_n873), .B1(new_n713), .B2(new_n714), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n664), .A2(new_n882), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n888), .A2(new_n876), .A3(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n729), .B1(new_n887), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n730), .A2(new_n771), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n893), .B(KEYINPUT113), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n482), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n446), .A2(new_n732), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n895), .A2(new_n532), .A3(new_n896), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n627), .A2(new_n629), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n897), .A2(new_n204), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n877), .A2(new_n884), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n665), .B1(new_n900), .B2(KEYINPUT115), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n877), .A2(new_n878), .A3(new_n884), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n891), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n894), .B1(new_n903), .B2(new_n804), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n904), .A2(new_n896), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n905), .A2(new_n758), .A3(new_n770), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n899), .B1(new_n906), .B2(new_n204), .ZN(G1340gat));
  OAI21_X1  g706(.A(G120gat), .B1(new_n897), .B2(new_n751), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n905), .A2(new_n758), .ZN(new_n909));
  OR2_X1    g708(.A1(new_n751), .A2(new_n208), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(G1341gat));
  OAI21_X1  g710(.A(G127gat), .B1(new_n897), .B2(new_n729), .ZN(new_n912));
  OR2_X1    g711(.A1(new_n729), .A2(G127gat), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n912), .B1(new_n909), .B2(new_n913), .ZN(G1342gat));
  OR2_X1    g713(.A1(new_n664), .A2(G134gat), .ZN(new_n915));
  OR3_X1    g714(.A1(new_n909), .A2(KEYINPUT56), .A3(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(G134gat), .B1(new_n897), .B2(new_n664), .ZN(new_n917));
  OAI21_X1  g716(.A(KEYINPUT56), .B1(new_n909), .B2(new_n915), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(G1343gat));
  NAND2_X1  g718(.A1(new_n744), .A2(new_n896), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g720(.A(KEYINPUT57), .B1(new_n904), .B2(new_n482), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT57), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n483), .A2(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  XNOR2_X1  g724(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n898), .B1(new_n875), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n874), .A2(new_n927), .A3(new_n715), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n665), .B1(new_n928), .B2(new_n884), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n729), .B1(new_n929), .B2(new_n891), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n925), .B1(new_n894), .B2(new_n930), .ZN(new_n931));
  OAI211_X1 g730(.A(new_n630), .B(new_n921), .C1(new_n922), .C2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(G141gat), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n333), .A2(new_n483), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n898), .A2(G141gat), .ZN(new_n935));
  AND4_X1   g734(.A1(new_n904), .A2(new_n896), .A3(new_n934), .A4(new_n935), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n936), .A2(KEYINPUT58), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n933), .A2(new_n937), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT58), .ZN(new_n939));
  OAI211_X1 g738(.A(new_n770), .B(new_n921), .C1(new_n922), .C2(new_n931), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n936), .B1(new_n940), .B2(G141gat), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n938), .B1(new_n939), .B2(new_n941), .ZN(G1344gat));
  INV_X1    g741(.A(KEYINPUT117), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n905), .A2(new_n934), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n751), .A2(G148gat), .ZN(new_n945));
  INV_X1    g744(.A(new_n945), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n943), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  NAND4_X1  g746(.A1(new_n905), .A2(KEYINPUT117), .A3(new_n934), .A4(new_n945), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT59), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(G148gat), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n904), .A2(new_n482), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(new_n923), .ZN(new_n953));
  INV_X1    g752(.A(new_n931), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n920), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n951), .B1(new_n955), .B2(new_n716), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT118), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n730), .A2(new_n898), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n483), .B1(new_n930), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n957), .B1(new_n959), .B2(KEYINPUT57), .ZN(new_n960));
  AOI22_X1  g759(.A1(new_n888), .A2(new_n927), .B1(new_n716), .B2(new_n883), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n890), .B1(new_n961), .B2(new_n665), .ZN(new_n962));
  AOI22_X1  g761(.A1(new_n962), .A2(new_n729), .B1(new_n898), .B2(new_n730), .ZN(new_n963));
  OAI211_X1 g762(.A(KEYINPUT118), .B(new_n923), .C1(new_n963), .C2(new_n483), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n960), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n925), .B1(new_n892), .B2(new_n894), .ZN(new_n966));
  OAI211_X1 g765(.A(new_n716), .B(new_n921), .C1(new_n965), .C2(new_n966), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n950), .B1(new_n967), .B2(G148gat), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n949), .B1(new_n956), .B2(new_n968), .ZN(G1345gat));
  NAND4_X1  g768(.A1(new_n904), .A2(new_n804), .A3(new_n896), .A4(new_n934), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n970), .A2(new_n337), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n921), .B1(new_n922), .B2(new_n931), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n729), .A2(new_n337), .ZN(new_n973));
  XNOR2_X1  g772(.A(new_n973), .B(KEYINPUT119), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n971), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT120), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OAI211_X1 g776(.A(KEYINPUT120), .B(new_n971), .C1(new_n972), .C2(new_n974), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n977), .A2(new_n978), .ZN(G1346gat));
  NAND3_X1  g778(.A1(new_n955), .A2(G162gat), .A3(new_n665), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n338), .B1(new_n944), .B2(new_n664), .ZN(new_n981));
  AND2_X1   g780(.A1(new_n980), .A2(new_n981), .ZN(G1347gat));
  NOR2_X1   g781(.A1(new_n735), .A2(new_n766), .ZN(new_n983));
  XNOR2_X1  g782(.A(new_n983), .B(KEYINPUT121), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n984), .A2(new_n331), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n895), .A2(new_n985), .ZN(new_n986));
  NOR3_X1   g785(.A1(new_n986), .A2(new_n232), .A3(new_n898), .ZN(new_n987));
  AND3_X1   g786(.A1(new_n904), .A2(new_n758), .A3(new_n983), .ZN(new_n988));
  AOI21_X1  g787(.A(G169gat), .B1(new_n988), .B2(new_n770), .ZN(new_n989));
  NOR2_X1   g788(.A1(new_n987), .A2(new_n989), .ZN(G1348gat));
  OAI21_X1  g789(.A(G176gat), .B1(new_n986), .B2(new_n751), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n988), .A2(new_n233), .A3(new_n716), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n991), .A2(new_n992), .ZN(G1349gat));
  INV_X1    g792(.A(KEYINPUT60), .ZN(new_n994));
  NOR2_X1   g793(.A1(new_n994), .A2(KEYINPUT123), .ZN(new_n995));
  AND2_X1   g794(.A1(new_n804), .A2(new_n220), .ZN(new_n996));
  AOI21_X1  g795(.A(new_n995), .B1(new_n988), .B2(new_n996), .ZN(new_n997));
  NAND3_X1  g796(.A1(new_n895), .A2(new_n804), .A3(new_n985), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n998), .A2(G183gat), .ZN(new_n999));
  OAI21_X1  g798(.A(KEYINPUT123), .B1(new_n994), .B2(KEYINPUT122), .ZN(new_n1000));
  XOR2_X1   g799(.A(new_n1000), .B(KEYINPUT124), .Z(new_n1001));
  AND3_X1   g800(.A1(new_n997), .A2(new_n999), .A3(new_n1001), .ZN(new_n1002));
  AOI21_X1  g801(.A(new_n1001), .B1(new_n997), .B2(new_n999), .ZN(new_n1003));
  NOR2_X1   g802(.A1(new_n1002), .A2(new_n1003), .ZN(G1350gat));
  NAND4_X1  g803(.A1(new_n904), .A2(new_n483), .A3(new_n665), .A4(new_n985), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1005), .A2(G190gat), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1006), .A2(KEYINPUT125), .ZN(new_n1007));
  INV_X1    g806(.A(KEYINPUT125), .ZN(new_n1008));
  NAND3_X1  g807(.A1(new_n1005), .A2(new_n1008), .A3(G190gat), .ZN(new_n1009));
  NAND3_X1  g808(.A1(new_n1007), .A2(KEYINPUT61), .A3(new_n1009), .ZN(new_n1010));
  NAND3_X1  g809(.A1(new_n988), .A2(new_n217), .A3(new_n665), .ZN(new_n1011));
  OAI211_X1 g810(.A(new_n1010), .B(new_n1011), .C1(KEYINPUT61), .C2(new_n1007), .ZN(G1351gat));
  NOR3_X1   g811(.A1(new_n333), .A2(new_n483), .A3(new_n735), .ZN(new_n1013));
  XNOR2_X1  g812(.A(new_n1013), .B(KEYINPUT126), .ZN(new_n1014));
  AND3_X1   g813(.A1(new_n1014), .A2(new_n732), .A3(new_n904), .ZN(new_n1015));
  AOI21_X1  g814(.A(G197gat), .B1(new_n1015), .B2(new_n770), .ZN(new_n1016));
  NOR2_X1   g815(.A1(new_n984), .A2(new_n333), .ZN(new_n1017));
  AND2_X1   g816(.A1(new_n630), .A2(G197gat), .ZN(new_n1018));
  OAI211_X1 g817(.A(new_n1017), .B(new_n1018), .C1(new_n965), .C2(new_n966), .ZN(new_n1019));
  INV_X1    g818(.A(new_n1019), .ZN(new_n1020));
  NOR2_X1   g819(.A1(new_n1016), .A2(new_n1020), .ZN(G1352gat));
  NOR2_X1   g820(.A1(new_n751), .A2(G204gat), .ZN(new_n1022));
  NAND4_X1  g821(.A1(new_n1014), .A2(new_n732), .A3(new_n904), .A4(new_n1022), .ZN(new_n1023));
  XOR2_X1   g822(.A(new_n1023), .B(KEYINPUT62), .Z(new_n1024));
  OAI21_X1  g823(.A(new_n1017), .B1(new_n965), .B2(new_n966), .ZN(new_n1025));
  OAI21_X1  g824(.A(G204gat), .B1(new_n1025), .B2(new_n751), .ZN(new_n1026));
  NAND2_X1  g825(.A1(new_n1024), .A2(new_n1026), .ZN(G1353gat));
  NAND3_X1  g826(.A1(new_n1015), .A2(new_n404), .A3(new_n804), .ZN(new_n1028));
  OAI211_X1 g827(.A(new_n804), .B(new_n1017), .C1(new_n965), .C2(new_n966), .ZN(new_n1029));
  AND3_X1   g828(.A1(new_n1029), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1030));
  AOI21_X1  g829(.A(KEYINPUT63), .B1(new_n1029), .B2(G211gat), .ZN(new_n1031));
  OAI21_X1  g830(.A(new_n1028), .B1(new_n1030), .B2(new_n1031), .ZN(G1354gat));
  NAND3_X1  g831(.A1(new_n1015), .A2(new_n405), .A3(new_n665), .ZN(new_n1033));
  OAI211_X1 g832(.A(new_n665), .B(new_n1017), .C1(new_n965), .C2(new_n966), .ZN(new_n1034));
  INV_X1    g833(.A(new_n1034), .ZN(new_n1035));
  OAI21_X1  g834(.A(new_n1033), .B1(new_n1035), .B2(new_n405), .ZN(G1355gat));
endmodule


