//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 0 1 0 1 1 0 1 1 1 0 1 1 0 1 0 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 0 1 1 0 1 0 0 0 1 0 1 1 0 0 0 1 0 1 1 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:32 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n554, new_n556, new_n557,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n584, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n626, new_n627, new_n629, new_n630, new_n632, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n868, new_n869, new_n870, new_n871,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT66), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT67), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(KEYINPUT68), .B(KEYINPUT2), .Z(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  OR4_X1    g028(.A1(G235), .A2(G238), .A3(G236), .A4(G237), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n454), .A2(G567), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT69), .Z(new_n458));
  NAND2_X1  g033(.A1(new_n453), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n462), .A2(G101), .A3(G2104), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT70), .ZN(new_n464));
  OR2_X1    g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n464), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G137), .ZN(new_n468));
  XNOR2_X1  g043(.A(KEYINPUT3), .B(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(new_n462), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n467), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  AOI22_X1  g046(.A1(new_n469), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(new_n462), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n471), .A2(new_n473), .ZN(G160));
  INV_X1    g049(.A(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(KEYINPUT3), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT3), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n479), .A2(new_n462), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n481), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  NAND4_X1  g062(.A1(new_n476), .A2(new_n478), .A3(G138), .A4(new_n462), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n469), .A2(KEYINPUT4), .A3(G138), .A4(new_n462), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n476), .A2(new_n478), .A3(G126), .A4(G2105), .ZN(new_n493));
  OR2_X1    g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n494), .A2(new_n496), .A3(G2104), .ZN(new_n497));
  AND3_X1   g072(.A1(new_n493), .A2(KEYINPUT71), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g073(.A(KEYINPUT71), .B1(new_n493), .B2(new_n497), .ZN(new_n499));
  NOR3_X1   g074(.A1(new_n492), .A2(new_n498), .A3(new_n499), .ZN(G164));
  XNOR2_X1  g075(.A(KEYINPUT5), .B(G543), .ZN(new_n501));
  AND2_X1   g076(.A1(new_n501), .A2(G62), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT73), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(G75), .A2(G543), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n506), .B1(new_n502), .B2(new_n503), .ZN(new_n507));
  OAI21_X1  g082(.A(G651), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n501), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT72), .A2(G651), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT6), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g087(.A1(KEYINPUT72), .A2(KEYINPUT6), .A3(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  OR2_X1    g090(.A1(new_n509), .A2(new_n515), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n508), .A2(new_n516), .ZN(G166));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  XNOR2_X1  g093(.A(new_n501), .B(KEYINPUT74), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G63), .ZN(new_n520));
  NAND3_X1  g095(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n518), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT75), .ZN(new_n523));
  INV_X1    g098(.A(new_n513), .ZN(new_n524));
  AOI21_X1  g099(.A(KEYINPUT6), .B1(KEYINPUT72), .B2(G651), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n512), .A2(KEYINPUT75), .A3(new_n513), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n526), .A2(G543), .A3(new_n527), .ZN(new_n528));
  XNOR2_X1  g103(.A(KEYINPUT76), .B(G51), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n514), .A2(new_n501), .ZN(new_n531));
  INV_X1    g106(.A(G89), .ZN(new_n532));
  AND3_X1   g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  OAI22_X1  g108(.A1(new_n531), .A2(new_n532), .B1(KEYINPUT7), .B2(new_n533), .ZN(new_n534));
  NOR3_X1   g109(.A1(new_n522), .A2(new_n530), .A3(new_n534), .ZN(G168));
  INV_X1    g110(.A(G52), .ZN(new_n536));
  INV_X1    g111(.A(G90), .ZN(new_n537));
  OAI22_X1  g112(.A1(new_n528), .A2(new_n536), .B1(new_n537), .B2(new_n531), .ZN(new_n538));
  NAND2_X1  g113(.A1(G77), .A2(G543), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT74), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n501), .B(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(G64), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n539), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n538), .B1(new_n543), .B2(G651), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT77), .ZN(G171));
  NAND2_X1  g120(.A1(new_n519), .A2(G56), .ZN(new_n546));
  NAND2_X1  g121(.A1(G68), .A2(G543), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n518), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(G43), .ZN(new_n549));
  INV_X1    g124(.A(G81), .ZN(new_n550));
  OAI22_X1  g125(.A1(new_n528), .A2(new_n549), .B1(new_n550), .B2(new_n531), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  AND3_X1   g128(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G36), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n554), .A2(new_n557), .ZN(G188));
  NAND4_X1  g133(.A1(new_n526), .A2(G53), .A3(new_n527), .A4(G543), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(KEYINPUT9), .ZN(new_n560));
  INV_X1    g135(.A(G543), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n561), .B1(new_n514), .B2(new_n523), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n562), .A2(new_n563), .A3(G53), .A4(new_n527), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT78), .ZN(new_n565));
  AND3_X1   g140(.A1(new_n560), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n565), .B1(new_n560), .B2(new_n564), .ZN(new_n567));
  OR2_X1    g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(G78), .ZN(new_n569));
  OAI21_X1  g144(.A(KEYINPUT79), .B1(new_n569), .B2(new_n561), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT79), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n571), .A2(G78), .A3(G543), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n501), .A2(G65), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT80), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n518), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n570), .A2(new_n572), .ZN(new_n576));
  XOR2_X1   g151(.A(KEYINPUT5), .B(G543), .Z(new_n577));
  INV_X1    g152(.A(G65), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(KEYINPUT80), .ZN(new_n580));
  AND2_X1   g155(.A1(new_n514), .A2(new_n501), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n575), .A2(new_n580), .B1(G91), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n568), .A2(new_n582), .ZN(G299));
  INV_X1    g158(.A(KEYINPUT77), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n544), .B(new_n584), .ZN(G301));
  INV_X1    g160(.A(G168), .ZN(G286));
  NAND2_X1  g161(.A1(new_n508), .A2(new_n516), .ZN(G303));
  NAND2_X1  g162(.A1(new_n581), .A2(G87), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n588), .B(KEYINPUT81), .ZN(new_n589));
  INV_X1    g164(.A(G74), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n541), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n528), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n591), .A2(G651), .B1(G49), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n589), .A2(new_n593), .ZN(G288));
  NAND2_X1  g169(.A1(new_n501), .A2(G61), .ZN(new_n595));
  NAND2_X1  g170(.A1(G73), .A2(G543), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n518), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT82), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n597), .B(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n501), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n600), .A2(new_n515), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n599), .A2(new_n602), .ZN(G305));
  AOI22_X1  g178(.A1(new_n592), .A2(G47), .B1(G85), .B2(new_n581), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n519), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(new_n518), .ZN(G290));
  INV_X1    g181(.A(KEYINPUT10), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT83), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n608), .B1(new_n581), .B2(G92), .ZN(new_n609));
  INV_X1    g184(.A(G92), .ZN(new_n610));
  NOR3_X1   g185(.A1(new_n531), .A2(KEYINPUT83), .A3(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n607), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n581), .A2(new_n608), .A3(G92), .ZN(new_n613));
  OAI21_X1  g188(.A(KEYINPUT83), .B1(new_n531), .B2(new_n610), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n613), .A2(KEYINPUT10), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(G79), .A2(G543), .ZN(new_n616));
  INV_X1    g191(.A(G66), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n577), .B2(new_n617), .ZN(new_n618));
  AOI22_X1  g193(.A1(new_n592), .A2(G54), .B1(G651), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n612), .A2(new_n615), .A3(new_n619), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n620), .A2(G868), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n621), .B1(G171), .B2(G868), .ZN(G284));
  AOI21_X1  g197(.A(new_n621), .B1(G171), .B2(G868), .ZN(G321));
  MUX2_X1   g198(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g199(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g200(.A(new_n620), .ZN(new_n626));
  INV_X1    g201(.A(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(G860), .ZN(G148));
  NAND2_X1  g203(.A1(new_n626), .A2(new_n627), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(G868), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(G868), .B2(new_n552), .ZN(G323));
  XNOR2_X1  g206(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n632));
  XNOR2_X1  g207(.A(G323), .B(new_n632), .ZN(G282));
  NAND2_X1  g208(.A1(new_n480), .A2(G2104), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT12), .ZN(new_n635));
  XOR2_X1   g210(.A(KEYINPUT85), .B(KEYINPUT13), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2100), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n635), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n480), .A2(G135), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n482), .A2(G123), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n462), .A2(G111), .ZN(new_n641));
  OAI21_X1  g216(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n642));
  OAI211_X1 g217(.A(new_n639), .B(new_n640), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(G2096), .Z(new_n644));
  NAND2_X1  g219(.A1(new_n638), .A2(new_n644), .ZN(G156));
  XNOR2_X1  g220(.A(G2451), .B(G2454), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n646), .B(new_n647), .Z(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2435), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2438), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2427), .B(G2430), .ZN(new_n651));
  INV_X1    g226(.A(KEYINPUT87), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n654), .A2(KEYINPUT14), .ZN(new_n655));
  AND2_X1   g230(.A1(new_n655), .A2(KEYINPUT88), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n655), .A2(KEYINPUT88), .ZN(new_n657));
  OAI22_X1  g232(.A1(new_n656), .A2(new_n657), .B1(new_n650), .B2(new_n653), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1341), .B(G1348), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n658), .A2(new_n659), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n648), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n662), .ZN(new_n664));
  INV_X1    g239(.A(new_n648), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n664), .A2(new_n665), .A3(new_n660), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n663), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n668), .A2(G14), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n667), .B1(new_n663), .B2(new_n666), .ZN(new_n670));
  OAI21_X1  g245(.A(KEYINPUT89), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(new_n670), .ZN(new_n672));
  INV_X1    g247(.A(KEYINPUT89), .ZN(new_n673));
  NAND4_X1  g248(.A1(new_n672), .A2(new_n673), .A3(G14), .A4(new_n668), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(G401));
  XOR2_X1   g251(.A(G2084), .B(G2090), .Z(new_n677));
  XNOR2_X1  g252(.A(G2072), .B(G2078), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT90), .ZN(new_n679));
  XNOR2_X1  g254(.A(G2067), .B(G2678), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n677), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n679), .B(KEYINPUT17), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n682), .B1(new_n683), .B2(new_n681), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT91), .Z(new_n685));
  INV_X1    g260(.A(new_n677), .ZN(new_n686));
  NOR3_X1   g261(.A1(new_n679), .A2(new_n681), .A3(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n687), .B(KEYINPUT18), .Z(new_n688));
  NOR2_X1   g263(.A1(new_n686), .A2(new_n680), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n688), .B1(new_n683), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n685), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(G2096), .B(G2100), .Z(new_n692));
  OR2_X1    g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n691), .A2(new_n692), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(G227));
  XNOR2_X1  g270(.A(G1971), .B(G1976), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT19), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(G1956), .B(G2474), .Z(new_n699));
  XOR2_X1   g274(.A(G1961), .B(G1966), .Z(new_n700));
  AND2_X1   g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(KEYINPUT20), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n699), .A2(new_n700), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n701), .A2(new_n705), .ZN(new_n706));
  MUX2_X1   g281(.A(new_n706), .B(new_n705), .S(new_n698), .Z(new_n707));
  NOR2_X1   g282(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(G1991), .B(G1996), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(G1981), .B(G1986), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(G229));
  INV_X1    g289(.A(G16), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G21), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G168), .B2(new_n715), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G1966), .ZN(new_n718));
  INV_X1    g293(.A(G29), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G27), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G164), .B2(new_n719), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT99), .B(G2078), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n721), .B(new_n722), .Z(new_n723));
  NAND2_X1  g298(.A1(new_n718), .A2(new_n723), .ZN(new_n724));
  AND2_X1   g299(.A1(KEYINPUT24), .A2(G34), .ZN(new_n725));
  NOR2_X1   g300(.A1(KEYINPUT24), .A2(G34), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n719), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT96), .Z(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(G160), .B2(G29), .ZN(new_n729));
  INV_X1    g304(.A(G2084), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT30), .B(G28), .ZN(new_n732));
  OR2_X1    g307(.A1(KEYINPUT31), .A2(G11), .ZN(new_n733));
  NAND2_X1  g308(.A1(KEYINPUT31), .A2(G11), .ZN(new_n734));
  AOI22_X1  g309(.A1(new_n732), .A2(new_n719), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(new_n643), .B2(new_n719), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n719), .A2(G33), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT25), .Z(new_n739));
  INV_X1    g314(.A(G139), .ZN(new_n740));
  AOI22_X1  g315(.A1(new_n469), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n741));
  OAI221_X1 g316(.A(new_n739), .B1(new_n470), .B2(new_n740), .C1(new_n741), .C2(new_n462), .ZN(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n737), .B1(new_n743), .B2(new_n719), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n736), .B1(new_n744), .B2(G2072), .ZN(new_n745));
  OAI211_X1 g320(.A(new_n731), .B(new_n745), .C1(G2072), .C2(new_n744), .ZN(new_n746));
  INV_X1    g321(.A(G1966), .ZN(new_n747));
  INV_X1    g322(.A(new_n717), .ZN(new_n748));
  AOI211_X1 g323(.A(new_n724), .B(new_n746), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(G171), .A2(G16), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G5), .B2(G16), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(G1961), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT100), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n480), .A2(G141), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT97), .ZN(new_n755));
  AND3_X1   g330(.A1(new_n462), .A2(G105), .A3(G2104), .ZN(new_n756));
  NAND3_X1  g331(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT26), .ZN(new_n758));
  AOI211_X1 g333(.A(new_n756), .B(new_n758), .C1(G129), .C2(new_n482), .ZN(new_n759));
  AOI21_X1  g334(.A(KEYINPUT98), .B1(new_n755), .B2(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(new_n760), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n755), .A2(KEYINPUT98), .A3(new_n759), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n719), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  AND2_X1   g338(.A1(new_n719), .A2(G32), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT27), .B(G1996), .ZN(new_n765));
  OR3_X1    g340(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n765), .B1(new_n763), .B2(new_n764), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND4_X1  g343(.A1(new_n749), .A2(new_n752), .A3(new_n753), .A4(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n770));
  INV_X1    g345(.A(new_n724), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n770), .A2(new_n768), .A3(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(G1961), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n751), .B(new_n773), .ZN(new_n774));
  OAI21_X1  g349(.A(KEYINPUT100), .B1(new_n772), .B2(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(G2067), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n480), .A2(G140), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n482), .A2(G128), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n462), .A2(G116), .ZN(new_n779));
  OAI21_X1  g354(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n780));
  OAI211_X1 g355(.A(new_n777), .B(new_n778), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n781), .A2(KEYINPUT95), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n781), .A2(KEYINPUT95), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n719), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n719), .A2(G26), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT28), .Z(new_n786));
  OAI21_X1  g361(.A(new_n776), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  OR3_X1    g362(.A1(new_n784), .A2(new_n776), .A3(new_n786), .ZN(new_n788));
  INV_X1    g363(.A(G2090), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n719), .A2(G35), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G162), .B2(new_n719), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n791), .A2(KEYINPUT29), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(KEYINPUT29), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n789), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT101), .ZN(new_n795));
  AOI22_X1  g370(.A1(new_n787), .A2(new_n788), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  OR2_X1    g371(.A1(new_n794), .A2(new_n795), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n792), .A2(new_n789), .A3(new_n793), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n715), .A2(G19), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(new_n552), .B2(new_n715), .ZN(new_n800));
  INV_X1    g375(.A(G1341), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NAND4_X1  g377(.A1(new_n796), .A2(new_n797), .A3(new_n798), .A4(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n715), .A2(G20), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT23), .Z(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(G299), .B2(G16), .ZN(new_n806));
  INV_X1    g381(.A(G1956), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(G4), .A2(G16), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT94), .Z(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(new_n620), .B2(new_n715), .ZN(new_n811));
  INV_X1    g386(.A(G1348), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NOR3_X1   g388(.A1(new_n803), .A2(new_n808), .A3(new_n813), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n769), .A2(new_n775), .A3(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT34), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n715), .A2(G22), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(G166), .B2(new_n715), .ZN(new_n818));
  INV_X1    g393(.A(G1971), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n818), .A2(new_n819), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(G288), .A2(G16), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n715), .A2(G23), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT33), .B(G1976), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n822), .A2(new_n828), .ZN(new_n829));
  MUX2_X1   g404(.A(G6), .B(G305), .S(G16), .Z(new_n830));
  XOR2_X1   g405(.A(KEYINPUT32), .B(G1981), .Z(new_n831));
  AND2_X1   g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n830), .A2(new_n831), .ZN(new_n833));
  OAI22_X1  g408(.A1(new_n832), .A2(new_n833), .B1(new_n826), .B2(new_n827), .ZN(new_n834));
  NOR3_X1   g409(.A1(new_n829), .A2(new_n834), .A3(KEYINPUT92), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT92), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n830), .A2(new_n831), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n830), .A2(new_n831), .ZN(new_n838));
  INV_X1    g413(.A(new_n827), .ZN(new_n839));
  AOI22_X1  g414(.A1(new_n837), .A2(new_n838), .B1(new_n825), .B2(new_n839), .ZN(new_n840));
  AOI22_X1  g415(.A1(new_n820), .A2(new_n821), .B1(new_n826), .B2(new_n827), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n836), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n816), .B1(new_n835), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(KEYINPUT92), .B1(new_n829), .B2(new_n834), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n840), .A2(new_n836), .A3(new_n841), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n844), .A2(KEYINPUT34), .A3(new_n845), .ZN(new_n846));
  MUX2_X1   g421(.A(G24), .B(G290), .S(G16), .Z(new_n847));
  AND2_X1   g422(.A1(new_n847), .A2(G1986), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n847), .A2(G1986), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n719), .A2(G25), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n480), .A2(G131), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n482), .A2(G119), .ZN(new_n852));
  OR2_X1    g427(.A1(G95), .A2(G2105), .ZN(new_n853));
  OAI211_X1 g428(.A(new_n853), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n851), .A2(new_n852), .A3(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n850), .B1(new_n856), .B2(new_n719), .ZN(new_n857));
  XOR2_X1   g432(.A(KEYINPUT35), .B(G1991), .Z(new_n858));
  XOR2_X1   g433(.A(new_n857), .B(new_n858), .Z(new_n859));
  NOR3_X1   g434(.A1(new_n848), .A2(new_n849), .A3(new_n859), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n843), .A2(new_n846), .A3(new_n860), .ZN(new_n861));
  AND2_X1   g436(.A1(KEYINPUT93), .A2(KEYINPUT36), .ZN(new_n862));
  NOR2_X1   g437(.A1(KEYINPUT93), .A2(KEYINPUT36), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n815), .B1(new_n861), .B2(new_n864), .ZN(new_n865));
  NAND4_X1  g440(.A1(new_n843), .A2(new_n846), .A3(new_n860), .A4(new_n862), .ZN(new_n866));
  AND2_X1   g441(.A1(new_n865), .A2(new_n866), .ZN(G311));
  NAND2_X1  g442(.A1(new_n861), .A2(new_n864), .ZN(new_n868));
  INV_X1    g443(.A(new_n815), .ZN(new_n869));
  AND4_X1   g444(.A1(KEYINPUT102), .A2(new_n868), .A3(new_n866), .A4(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(KEYINPUT102), .B1(new_n865), .B2(new_n866), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n870), .A2(new_n871), .ZN(G150));
  NAND2_X1  g447(.A1(new_n519), .A2(G67), .ZN(new_n873));
  NAND2_X1  g448(.A1(G80), .A2(G543), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n518), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(G55), .ZN(new_n876));
  INV_X1    g451(.A(G93), .ZN(new_n877));
  OAI22_X1  g452(.A1(new_n528), .A2(new_n876), .B1(new_n877), .B2(new_n531), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(G860), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT37), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n626), .A2(G559), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT38), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n552), .A2(new_n879), .ZN(new_n885));
  OAI22_X1  g460(.A1(new_n548), .A2(new_n551), .B1(new_n875), .B2(new_n878), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n884), .B(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(KEYINPUT39), .ZN(new_n890));
  XOR2_X1   g465(.A(new_n890), .B(KEYINPUT103), .Z(new_n891));
  OAI21_X1  g466(.A(new_n880), .B1(new_n889), .B2(KEYINPUT39), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n882), .B1(new_n891), .B2(new_n892), .ZN(G145));
  XNOR2_X1  g468(.A(G162), .B(new_n643), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(G160), .ZN(new_n895));
  AND2_X1   g470(.A1(new_n782), .A2(new_n783), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n896), .A2(new_n761), .A3(new_n762), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n782), .A2(new_n783), .ZN(new_n898));
  INV_X1    g473(.A(new_n762), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n898), .B1(new_n899), .B2(new_n760), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n742), .B1(new_n897), .B2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n490), .A2(new_n491), .A3(KEYINPUT104), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n493), .A2(new_n497), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT104), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n904), .B1(new_n492), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n897), .A2(new_n900), .A3(new_n742), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n902), .A2(new_n903), .A3(new_n906), .A4(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n480), .A2(G142), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n482), .A2(G130), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n462), .A2(G118), .ZN(new_n911));
  OAI21_X1  g486(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n912));
  OAI211_X1 g487(.A(new_n909), .B(new_n910), .C1(new_n911), .C2(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n635), .B(new_n913), .ZN(new_n914));
  OR2_X1    g489(.A1(new_n914), .A2(new_n856), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n856), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT105), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n915), .A2(KEYINPUT105), .A3(new_n916), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n492), .A2(new_n905), .ZN(new_n922));
  INV_X1    g497(.A(new_n904), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n922), .A2(new_n923), .A3(new_n903), .ZN(new_n924));
  INV_X1    g499(.A(new_n907), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n924), .B1(new_n925), .B2(new_n901), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n908), .A2(new_n921), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n921), .B1(new_n908), .B2(new_n926), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n895), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT106), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI211_X1 g506(.A(KEYINPUT106), .B(new_n895), .C1(new_n927), .C2(new_n928), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n928), .A2(new_n895), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n908), .A2(new_n926), .A3(new_n916), .A4(new_n915), .ZN(new_n935));
  AOI21_X1  g510(.A(G37), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n933), .A2(KEYINPUT40), .A3(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(KEYINPUT40), .B1(new_n933), .B2(new_n936), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n938), .A2(new_n939), .ZN(G395));
  XNOR2_X1  g515(.A(new_n887), .B(new_n629), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n626), .B1(new_n568), .B2(new_n582), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n568), .A2(new_n626), .A3(new_n582), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n941), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT41), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n944), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n949), .A2(new_n942), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(KEYINPUT41), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n948), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n946), .B1(new_n952), .B2(new_n941), .ZN(new_n953));
  OR2_X1    g528(.A1(new_n953), .A2(KEYINPUT42), .ZN(new_n954));
  XOR2_X1   g529(.A(G288), .B(G305), .Z(new_n955));
  XNOR2_X1  g530(.A(G166), .B(G290), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n955), .B(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n953), .A2(KEYINPUT42), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n954), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n958), .B1(new_n954), .B2(new_n959), .ZN(new_n961));
  OAI21_X1  g536(.A(G868), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n962), .B1(G868), .B2(new_n879), .ZN(G295));
  OAI21_X1  g538(.A(new_n962), .B1(G868), .B2(new_n879), .ZN(G331));
  XNOR2_X1  g539(.A(KEYINPUT107), .B(KEYINPUT44), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n887), .A2(G301), .ZN(new_n966));
  NAND3_X1  g541(.A1(G171), .A2(new_n886), .A3(new_n885), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(G286), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n966), .A2(new_n967), .A3(G168), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n952), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n969), .A2(new_n950), .A3(new_n970), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n972), .A2(new_n973), .A3(new_n957), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n957), .B1(new_n972), .B2(new_n973), .ZN(new_n976));
  NOR4_X1   g551(.A1(new_n975), .A2(new_n976), .A3(KEYINPUT43), .A4(G37), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT43), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n972), .A2(new_n973), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n957), .A2(KEYINPUT108), .ZN(new_n980));
  AOI21_X1  g555(.A(G37), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n972), .B(new_n973), .C1(KEYINPUT108), .C2(new_n957), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n978), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n965), .B1(new_n977), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n981), .A2(new_n978), .A3(new_n982), .ZN(new_n985));
  NOR3_X1   g560(.A1(new_n975), .A2(G37), .A3(new_n976), .ZN(new_n986));
  OAI211_X1 g561(.A(new_n985), .B(KEYINPUT44), .C1(new_n986), .C2(new_n978), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n984), .A2(new_n987), .ZN(G397));
  INV_X1    g563(.A(G1384), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n924), .A2(new_n989), .ZN(new_n990));
  XOR2_X1   g565(.A(KEYINPUT109), .B(KEYINPUT45), .Z(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  AOI22_X1  g567(.A1(new_n480), .A2(G137), .B1(new_n465), .B2(new_n466), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n993), .B(G40), .C1(new_n462), .C2(new_n472), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n761), .A2(new_n762), .ZN(new_n996));
  INV_X1    g571(.A(G1996), .ZN(new_n997));
  XNOR2_X1  g572(.A(new_n996), .B(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n896), .A2(new_n776), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n898), .A2(G2067), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n998), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n856), .A2(new_n858), .ZN(new_n1004));
  OR2_X1    g579(.A1(new_n856), .A2(new_n858), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g581(.A(G290), .B(G1986), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n995), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT63), .ZN(new_n1009));
  NOR2_X1   g584(.A1(KEYINPUT112), .A2(KEYINPUT55), .ZN(new_n1010));
  AND2_X1   g585(.A1(KEYINPUT112), .A2(KEYINPUT55), .ZN(new_n1011));
  OAI211_X1 g586(.A(G303), .B(G8), .C1(new_n1010), .C2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(G8), .ZN(new_n1013));
  NOR2_X1   g588(.A1(G166), .A2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1012), .B1(new_n1014), .B2(new_n1011), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT71), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n904), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n493), .A2(KEYINPUT71), .A3(new_n497), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n989), .B1(new_n1020), .B2(new_n492), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n994), .B1(new_n1021), .B2(new_n991), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n924), .A2(KEYINPUT45), .A3(new_n989), .ZN(new_n1023));
  AOI21_X1  g598(.A(G1971), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G40), .ZN(new_n1025));
  NOR3_X1   g600(.A1(new_n471), .A2(new_n473), .A3(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(G1384), .B1(new_n906), .B2(new_n903), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT50), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1026), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n498), .A2(new_n499), .ZN(new_n1030));
  INV_X1    g605(.A(new_n492), .ZN(new_n1031));
  AOI21_X1  g606(.A(G1384), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1032), .A2(KEYINPUT117), .A3(new_n1028), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT117), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1034), .B1(new_n1021), .B2(KEYINPUT50), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1029), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g611(.A(KEYINPUT110), .B(G2090), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1024), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1016), .B1(new_n1038), .B2(new_n1013), .ZN(new_n1039));
  INV_X1    g614(.A(G1976), .ZN(new_n1040));
  OR3_X1    g615(.A1(G288), .A2(KEYINPUT114), .A3(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1013), .B1(new_n1027), .B2(new_n1026), .ZN(new_n1042));
  OAI21_X1  g617(.A(KEYINPUT114), .B1(G288), .B2(new_n1040), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT52), .ZN(new_n1045));
  INV_X1    g620(.A(G1981), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n599), .A2(new_n1046), .A3(new_n602), .ZN(new_n1047));
  OAI21_X1  g622(.A(G1981), .B1(new_n601), .B2(new_n597), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  OR2_X1    g624(.A1(KEYINPUT115), .A2(KEYINPUT49), .ZN(new_n1050));
  XNOR2_X1  g625(.A(new_n1049), .B(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(new_n1042), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT52), .B1(G288), .B2(new_n1040), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .A4(new_n1053), .ZN(new_n1054));
  AND3_X1   g629(.A1(new_n1045), .A2(new_n1052), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT111), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n994), .B1(new_n1021), .B2(KEYINPUT50), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n924), .A2(new_n1028), .A3(new_n989), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n1057), .A2(new_n1037), .A3(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1056), .B1(new_n1059), .B2(new_n1024), .ZN(new_n1060));
  INV_X1    g635(.A(new_n991), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1026), .B1(new_n1032), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT45), .ZN(new_n1063));
  AOI211_X1 g638(.A(new_n1063), .B(G1384), .C1(new_n906), .C2(new_n903), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n819), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1057), .A2(new_n1037), .A3(new_n1058), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1065), .A2(KEYINPUT111), .A3(new_n1066), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1060), .A2(G8), .A3(new_n1015), .A4(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT113), .ZN(new_n1069));
  AND2_X1   g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1039), .B(new_n1055), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1027), .A2(KEYINPUT45), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1026), .B1(new_n1021), .B2(new_n991), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n747), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1057), .A2(new_n730), .A3(new_n1058), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1077), .A2(G8), .A3(G168), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1009), .B1(new_n1072), .B2(new_n1078), .ZN(new_n1079));
  AND2_X1   g654(.A1(new_n1067), .A2(G8), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1015), .B1(new_n1080), .B2(new_n1060), .ZN(new_n1081));
  NOR3_X1   g656(.A1(new_n1081), .A2(new_n1009), .A3(new_n1078), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1080), .A2(KEYINPUT113), .A3(new_n1015), .A4(new_n1060), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1082), .A2(new_n1085), .A3(new_n1055), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1079), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1072), .A2(KEYINPUT126), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1075), .A2(G168), .A3(new_n1076), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(G8), .ZN(new_n1090));
  AOI21_X1  g665(.A(G168), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1091));
  OAI21_X1  g666(.A(KEYINPUT51), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT62), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT51), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1089), .A2(new_n1094), .A3(G8), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n1092), .A2(new_n1093), .A3(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1093), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1097));
  AOI21_X1  g672(.A(G1961), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT53), .ZN(new_n1099));
  INV_X1    g674(.A(G2078), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1022), .A2(new_n1100), .A3(new_n1023), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1098), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1099), .A2(G2078), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(G301), .B1(new_n1102), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  NOR3_X1   g682(.A1(new_n1096), .A2(new_n1097), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT126), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1085), .A2(new_n1109), .A3(new_n1039), .A4(new_n1055), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1088), .A2(new_n1108), .A3(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1055), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1112));
  AOI211_X1 g687(.A(G1976), .B(G288), .C1(new_n1051), .C2(new_n1042), .ZN(new_n1113));
  XOR2_X1   g688(.A(new_n1047), .B(KEYINPUT116), .Z(new_n1114));
  OAI21_X1  g689(.A(new_n1042), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  AND2_X1   g690(.A1(new_n1112), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1087), .A2(new_n1111), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1029), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1035), .A2(new_n1033), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1121));
  XOR2_X1   g696(.A(KEYINPUT120), .B(KEYINPUT56), .Z(new_n1122));
  XNOR2_X1  g697(.A(new_n1122), .B(G2072), .ZN(new_n1123));
  AOI22_X1  g698(.A1(new_n1120), .A2(new_n807), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT119), .ZN(new_n1125));
  XOR2_X1   g700(.A(KEYINPUT118), .B(KEYINPUT57), .Z(new_n1126));
  INV_X1    g701(.A(new_n582), .ZN(new_n1127));
  AND2_X1   g702(.A1(new_n560), .A2(new_n564), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1126), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  OAI211_X1 g704(.A(KEYINPUT57), .B(new_n582), .C1(new_n566), .C2(new_n567), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1125), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1129), .A2(new_n1130), .A3(new_n1125), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1124), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1124), .A2(new_n1134), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1026), .B1(new_n1032), .B2(new_n1028), .ZN(new_n1138));
  AOI211_X1 g713(.A(KEYINPUT50), .B(G1384), .C1(new_n906), .C2(new_n903), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n812), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1027), .A2(new_n776), .A3(new_n1026), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n620), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1137), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT61), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1144), .A2(KEYINPUT123), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1146), .B1(new_n1036), .B2(G1956), .ZN(new_n1147));
  AND3_X1   g722(.A1(new_n1129), .A2(new_n1130), .A3(new_n1125), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1148), .A2(new_n1131), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1145), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1145), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1124), .A2(new_n1134), .A3(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT124), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n612), .A2(new_n1154), .A3(new_n619), .A4(new_n615), .ZN(new_n1155));
  AND2_X1   g730(.A1(new_n1155), .A2(KEYINPUT60), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1140), .A2(new_n1141), .A3(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n620), .A2(KEYINPUT124), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1140), .A2(new_n1156), .A3(new_n1141), .A4(new_n1158), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT60), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1160), .A2(new_n1161), .A3(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n991), .B1(G164), .B2(G1384), .ZN(new_n1166));
  XNOR2_X1  g741(.A(KEYINPUT121), .B(G1996), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1023), .A2(new_n1166), .A3(new_n1026), .A4(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g743(.A(KEYINPUT122), .B(KEYINPUT58), .ZN(new_n1169));
  XNOR2_X1  g744(.A(new_n1169), .B(new_n801), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1170), .B1(new_n990), .B2(new_n994), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1168), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(new_n552), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1173), .A2(KEYINPUT59), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT59), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1172), .A2(new_n1175), .A3(new_n552), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1165), .A2(new_n1177), .ZN(new_n1178));
  OAI211_X1 g753(.A(new_n1136), .B(new_n1143), .C1(new_n1153), .C2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1179), .A2(KEYINPUT125), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT125), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1135), .B1(new_n1137), .B2(new_n1142), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1135), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1183));
  OAI211_X1 g758(.A(new_n1181), .B(new_n1182), .C1(new_n1183), .C2(new_n1178), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT54), .ZN(new_n1185));
  NAND4_X1  g760(.A1(new_n992), .A2(new_n1023), .A3(new_n1026), .A4(new_n1104), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1102), .A2(new_n1186), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n1187), .A2(G171), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1185), .B1(new_n1188), .B2(new_n1106), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1187), .A2(G171), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1102), .A2(G301), .A3(new_n1105), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1191), .A2(KEYINPUT54), .A3(new_n1192), .ZN(new_n1193));
  AND3_X1   g768(.A1(new_n1189), .A2(new_n1190), .A3(new_n1193), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1180), .A2(new_n1184), .A3(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1088), .A2(new_n1110), .ZN(new_n1196));
  NOR2_X1   g771(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1008), .B1(new_n1117), .B2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1006), .A2(new_n995), .ZN(new_n1199));
  OR2_X1    g774(.A1(new_n1199), .A2(KEYINPUT127), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1199), .A2(KEYINPUT127), .ZN(new_n1201));
  NOR2_X1   g776(.A1(G290), .A2(G1986), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n995), .A2(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g778(.A(new_n1203), .B(KEYINPUT48), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1200), .A2(new_n1201), .A3(new_n1204), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n995), .B1(new_n1001), .B2(new_n996), .ZN(new_n1206));
  NOR3_X1   g781(.A1(new_n992), .A2(G1996), .A3(new_n994), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1207), .A2(KEYINPUT46), .ZN(new_n1208));
  OR2_X1    g783(.A1(new_n1207), .A2(KEYINPUT46), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1206), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  XNOR2_X1  g785(.A(new_n1210), .B(KEYINPUT47), .ZN(new_n1211));
  INV_X1    g786(.A(new_n1003), .ZN(new_n1212));
  OAI21_X1  g787(.A(new_n999), .B1(new_n1212), .B2(new_n1004), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1213), .A2(new_n995), .ZN(new_n1214));
  AND3_X1   g789(.A1(new_n1205), .A2(new_n1211), .A3(new_n1214), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1198), .A2(new_n1215), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g791(.A1(new_n976), .A2(G37), .ZN(new_n1218));
  NAND3_X1  g792(.A1(new_n1218), .A2(new_n978), .A3(new_n974), .ZN(new_n1219));
  NAND2_X1  g793(.A1(new_n979), .A2(new_n980), .ZN(new_n1220));
  INV_X1    g794(.A(G37), .ZN(new_n1221));
  AND3_X1   g795(.A1(new_n1220), .A2(new_n1221), .A3(new_n982), .ZN(new_n1222));
  OAI21_X1  g796(.A(new_n1219), .B1(new_n1222), .B2(new_n978), .ZN(new_n1223));
  NAND3_X1  g797(.A1(new_n693), .A2(G319), .A3(new_n694), .ZN(new_n1224));
  NOR2_X1   g798(.A1(G229), .A2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g799(.A1(new_n1225), .A2(new_n675), .ZN(new_n1226));
  AOI21_X1  g800(.A(new_n1226), .B1(new_n933), .B2(new_n936), .ZN(new_n1227));
  AND2_X1   g801(.A1(new_n1223), .A2(new_n1227), .ZN(G308));
  NAND2_X1  g802(.A1(new_n1223), .A2(new_n1227), .ZN(G225));
endmodule


