//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 1 1 0 1 1 1 0 1 1 1 1 1 0 1 0 0 1 0 0 1 1 0 1 0 0 0 0 1 1 1 0 1 0 1 0 0 0 1 0 0 0 1 1 1 0 0 1 0 1 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:23 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n701, new_n702, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G107), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G104), .ZN(new_n191));
  AND2_X1   g005(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n192));
  NOR2_X1   g006(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n191), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G101), .ZN(new_n195));
  XNOR2_X1  g009(.A(G104), .B(G107), .ZN(new_n196));
  OAI211_X1 g010(.A(new_n194), .B(new_n195), .C1(new_n196), .C2(new_n192), .ZN(new_n197));
  OR2_X1    g011(.A1(new_n196), .A2(new_n195), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT78), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT78), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n197), .A2(new_n201), .A3(new_n198), .ZN(new_n202));
  INV_X1    g016(.A(G146), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G143), .ZN(new_n204));
  INV_X1    g018(.A(G143), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G146), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT1), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n204), .A2(new_n206), .A3(new_n207), .A4(G128), .ZN(new_n208));
  INV_X1    g022(.A(G128), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n209), .B1(new_n204), .B2(KEYINPUT1), .ZN(new_n210));
  XNOR2_X1  g024(.A(G143), .B(G146), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n208), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AND2_X1   g026(.A1(new_n212), .A2(KEYINPUT10), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n200), .A2(new_n202), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT79), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT79), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n200), .A2(new_n216), .A3(new_n202), .A4(new_n213), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G134), .ZN(new_n219));
  OAI21_X1  g033(.A(KEYINPUT11), .B1(new_n219), .B2(G137), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT11), .ZN(new_n221));
  INV_X1    g035(.A(G137), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n221), .A2(new_n222), .A3(G134), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT65), .B1(new_n222), .B2(G134), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT65), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n226), .A2(new_n219), .A3(G137), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n224), .A2(new_n225), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G131), .ZN(new_n229));
  INV_X1    g043(.A(G131), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n224), .A2(new_n230), .A3(new_n225), .A4(new_n227), .ZN(new_n231));
  AND2_X1   g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  NOR3_X1   g046(.A1(new_n211), .A2(KEYINPUT0), .A3(new_n209), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n204), .A2(new_n206), .A3(G128), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT0), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n235), .A2(new_n209), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n234), .B1(new_n211), .B2(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n233), .B1(KEYINPUT0), .B2(new_n237), .ZN(new_n238));
  OR2_X1    g052(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n239));
  NAND2_X1  g053(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n240));
  AOI22_X1  g054(.A1(new_n239), .A2(new_n240), .B1(G104), .B2(new_n190), .ZN(new_n241));
  INV_X1    g055(.A(G104), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G107), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n192), .B1(new_n243), .B2(new_n191), .ZN(new_n244));
  OAI21_X1  g058(.A(G101), .B1(new_n241), .B2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n245), .A2(KEYINPUT4), .A3(new_n197), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n247), .B(G101), .C1(new_n241), .C2(new_n244), .ZN(new_n248));
  AND2_X1   g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  AND2_X1   g063(.A1(new_n197), .A2(new_n198), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT77), .ZN(new_n251));
  INV_X1    g065(.A(new_n211), .ZN(new_n252));
  OAI211_X1 g066(.A(KEYINPUT76), .B(KEYINPUT1), .C1(new_n205), .C2(G146), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G128), .ZN(new_n254));
  AOI21_X1  g068(.A(KEYINPUT76), .B1(new_n204), .B2(KEYINPUT1), .ZN(new_n255));
  OAI211_X1 g069(.A(new_n251), .B(new_n252), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(new_n208), .ZN(new_n257));
  OAI21_X1  g071(.A(KEYINPUT1), .B1(new_n205), .B2(G146), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT76), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n260), .A2(G128), .A3(new_n253), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n251), .B1(new_n261), .B2(new_n252), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n250), .B1(new_n257), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT10), .ZN(new_n264));
  AOI22_X1  g078(.A1(new_n238), .A2(new_n249), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n218), .A2(new_n232), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(KEYINPUT80), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT80), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n218), .A2(new_n268), .A3(new_n265), .A4(new_n232), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n218), .A2(new_n265), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n229), .A2(new_n231), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g088(.A(G110), .B(G140), .ZN(new_n275));
  INV_X1    g089(.A(G953), .ZN(new_n276));
  AND2_X1   g090(.A1(new_n276), .A2(G227), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n275), .B(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n274), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n212), .ZN(new_n280));
  INV_X1    g094(.A(new_n202), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n201), .B1(new_n197), .B2(new_n198), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(new_n263), .ZN(new_n284));
  AOI21_X1  g098(.A(KEYINPUT12), .B1(new_n284), .B2(new_n272), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT12), .ZN(new_n286));
  AOI211_X1 g100(.A(new_n286), .B(new_n232), .C1(new_n283), .C2(new_n263), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n278), .B1(new_n267), .B2(new_n269), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT81), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n289), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  AOI211_X1 g106(.A(KEYINPUT81), .B(new_n278), .C1(new_n267), .C2(new_n269), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n279), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G469), .ZN(new_n295));
  INV_X1    g109(.A(G902), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n288), .B1(new_n267), .B2(new_n269), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  AOI22_X1  g113(.A1(new_n299), .A2(new_n278), .B1(new_n290), .B2(new_n273), .ZN(new_n300));
  OAI21_X1  g114(.A(G469), .B1(new_n300), .B2(G902), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n189), .B1(new_n297), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT67), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n219), .A2(G137), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n222), .A2(G134), .ZN(new_n305));
  OAI21_X1  g119(.A(G131), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AND3_X1   g120(.A1(new_n231), .A2(new_n212), .A3(new_n306), .ZN(new_n307));
  AOI22_X1  g121(.A1(new_n303), .A2(new_n307), .B1(new_n272), .B2(new_n238), .ZN(new_n308));
  NOR2_X1   g122(.A1(KEYINPUT2), .A2(G113), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(KEYINPUT66), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT66), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n311), .B1(KEYINPUT2), .B2(G113), .ZN(new_n312));
  AOI22_X1  g126(.A1(new_n310), .A2(new_n312), .B1(KEYINPUT2), .B2(G113), .ZN(new_n313));
  XNOR2_X1  g127(.A(G116), .B(G119), .ZN(new_n314));
  XOR2_X1   g128(.A(new_n313), .B(new_n314), .Z(new_n315));
  NAND3_X1  g129(.A1(new_n231), .A2(new_n212), .A3(new_n306), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(KEYINPUT67), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n308), .A2(KEYINPUT68), .A3(new_n315), .A4(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n272), .A2(new_n238), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n231), .A2(new_n212), .A3(new_n303), .A4(new_n306), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n319), .A2(new_n315), .A3(new_n317), .A4(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT68), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n318), .A2(new_n323), .A3(KEYINPUT28), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n307), .B1(new_n272), .B2(new_n238), .ZN(new_n325));
  AOI21_X1  g139(.A(KEYINPUT28), .B1(new_n325), .B2(new_n315), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n325), .A2(new_n315), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n324), .A2(new_n328), .ZN(new_n329));
  NOR2_X1   g143(.A1(G237), .A2(G953), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G210), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n331), .B(KEYINPUT27), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT26), .B(G101), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n332), .B(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n329), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n318), .A2(new_n323), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n319), .A2(new_n316), .ZN(new_n338));
  XNOR2_X1  g152(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n319), .A2(KEYINPUT30), .A3(new_n317), .A4(new_n320), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n313), .B(new_n314), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n337), .A2(new_n334), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(KEYINPUT31), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT31), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n337), .A2(new_n346), .A3(new_n343), .A4(new_n334), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n336), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(G472), .A2(G902), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(KEYINPUT69), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT32), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT69), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n348), .A2(new_n353), .A3(new_n349), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n351), .A2(new_n352), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n337), .A2(new_n343), .ZN(new_n356));
  AOI21_X1  g170(.A(KEYINPUT29), .B1(new_n356), .B2(new_n335), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n357), .B1(new_n335), .B2(new_n329), .ZN(new_n358));
  INV_X1    g172(.A(new_n326), .ZN(new_n359));
  AND2_X1   g173(.A1(new_n334), .A2(KEYINPUT29), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n308), .A2(new_n317), .ZN(new_n361));
  AOI22_X1  g175(.A1(new_n318), .A2(new_n323), .B1(new_n342), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT28), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n359), .B(new_n360), .C1(new_n362), .C2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(KEYINPUT70), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n358), .A2(new_n296), .A3(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n364), .A2(KEYINPUT70), .ZN(new_n367));
  OAI21_X1  g181(.A(G472), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n348), .A2(KEYINPUT32), .A3(new_n349), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n355), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT72), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT23), .ZN(new_n372));
  AOI22_X1  g186(.A1(new_n371), .A2(new_n372), .B1(new_n209), .B2(G119), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n373), .B1(new_n371), .B2(new_n372), .ZN(new_n374));
  OAI21_X1  g188(.A(KEYINPUT71), .B1(new_n209), .B2(G119), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n209), .A2(KEYINPUT23), .A3(G119), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT71), .ZN(new_n378));
  OAI211_X1 g192(.A(new_n374), .B(new_n377), .C1(new_n378), .C2(new_n376), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G110), .ZN(new_n380));
  XNOR2_X1  g194(.A(G125), .B(G140), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(KEYINPUT16), .ZN(new_n382));
  INV_X1    g196(.A(G125), .ZN(new_n383));
  OR3_X1    g197(.A1(new_n383), .A2(KEYINPUT16), .A3(G140), .ZN(new_n384));
  AOI21_X1  g198(.A(G146), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n382), .A2(G146), .A3(new_n384), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  XOR2_X1   g201(.A(G119), .B(G128), .Z(new_n388));
  XNOR2_X1  g202(.A(KEYINPUT24), .B(G110), .ZN(new_n389));
  OAI221_X1 g203(.A(new_n380), .B1(new_n385), .B2(new_n387), .C1(new_n388), .C2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n388), .A2(new_n389), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n391), .B1(new_n379), .B2(G110), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n381), .A2(new_n203), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n392), .A2(new_n386), .A3(new_n393), .ZN(new_n394));
  AND2_X1   g208(.A1(new_n390), .A2(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(KEYINPUT22), .B(G137), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n276), .A2(G221), .A3(G234), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n396), .B(new_n397), .ZN(new_n398));
  XOR2_X1   g212(.A(new_n398), .B(KEYINPUT73), .Z(new_n399));
  OR2_X1    g213(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n395), .A2(new_n398), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n400), .A2(new_n296), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT25), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n400), .A2(KEYINPUT25), .A3(new_n296), .A4(new_n401), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(G217), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n407), .B1(G234), .B2(new_n296), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  AND2_X1   g223(.A1(new_n400), .A2(new_n401), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n408), .A2(G902), .ZN(new_n411));
  XOR2_X1   g225(.A(new_n411), .B(KEYINPUT74), .Z(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n409), .A2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(G214), .B1(G237), .B2(G902), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  AND3_X1   g232(.A1(new_n342), .A2(new_n246), .A3(new_n248), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(G110), .B(G122), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n313), .A2(new_n314), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n314), .A2(KEYINPUT5), .ZN(new_n423));
  INV_X1    g237(.A(G116), .ZN(new_n424));
  OR2_X1    g238(.A1(new_n424), .A2(G119), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n423), .B(G113), .C1(KEYINPUT5), .C2(new_n425), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n200), .A2(new_n422), .A3(new_n202), .A4(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n420), .A2(new_n421), .A3(new_n427), .ZN(new_n428));
  AND2_X1   g242(.A1(new_n237), .A2(KEYINPUT0), .ZN(new_n429));
  OAI21_X1  g243(.A(G125), .B1(new_n429), .B2(new_n233), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n280), .A2(new_n383), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT84), .ZN(new_n432));
  INV_X1    g246(.A(G224), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n433), .A2(G953), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT7), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n430), .B(new_n431), .C1(new_n432), .C2(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n436), .B1(new_n430), .B2(new_n432), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n430), .A2(new_n431), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  AND3_X1   g254(.A1(new_n428), .A2(new_n437), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n426), .A2(new_n422), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(new_n199), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n427), .A2(new_n443), .ZN(new_n444));
  XOR2_X1   g258(.A(new_n421), .B(KEYINPUT8), .Z(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(KEYINPUT83), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n444), .A2(new_n446), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT83), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n441), .B1(new_n447), .B2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n421), .ZN(new_n452));
  INV_X1    g266(.A(new_n427), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n452), .B1(new_n453), .B2(new_n419), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n454), .A2(new_n428), .A3(KEYINPUT6), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n434), .B(KEYINPUT82), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n439), .B(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT6), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n458), .B(new_n452), .C1(new_n453), .C2(new_n419), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n455), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n451), .A2(new_n296), .A3(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(G210), .B1(G237), .B2(G902), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n448), .B(new_n449), .ZN(new_n465));
  AOI21_X1  g279(.A(G902), .B1(new_n465), .B2(new_n441), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n466), .A2(new_n462), .A3(new_n460), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n418), .B1(new_n464), .B2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(G952), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n469), .A2(G953), .ZN(new_n470));
  INV_X1    g284(.A(G234), .ZN(new_n471));
  INV_X1    g285(.A(G237), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  AOI211_X1 g288(.A(new_n296), .B(new_n276), .C1(G234), .C2(G237), .ZN(new_n475));
  XNOR2_X1  g289(.A(KEYINPUT21), .B(G898), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT85), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n330), .A2(G214), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n205), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n330), .A2(G143), .A3(G214), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(KEYINPUT18), .A2(G131), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n479), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n483), .A2(KEYINPUT85), .A3(KEYINPUT18), .A4(G131), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OR2_X1    g302(.A1(new_n381), .A2(new_n203), .ZN(new_n489));
  AOI22_X1  g303(.A1(new_n484), .A2(new_n485), .B1(new_n489), .B2(new_n393), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  OR3_X1    g305(.A1(new_n387), .A2(new_n385), .A3(KEYINPUT87), .ZN(new_n492));
  OAI21_X1  g306(.A(KEYINPUT87), .B1(new_n387), .B2(new_n385), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n483), .A2(KEYINPUT17), .A3(G131), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n483), .B(G131), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n495), .B1(new_n496), .B2(KEYINPUT17), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n491), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  XNOR2_X1  g312(.A(G113), .B(G122), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n499), .B(new_n242), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n500), .B(new_n491), .C1(new_n494), .C2(new_n497), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(new_n296), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(G475), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n381), .B(KEYINPUT19), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n387), .B1(new_n203), .B2(new_n507), .ZN(new_n508));
  AOI22_X1  g322(.A1(new_n488), .A2(new_n490), .B1(new_n508), .B2(new_n496), .ZN(new_n509));
  OAI21_X1  g323(.A(KEYINPUT86), .B1(new_n509), .B2(new_n500), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n508), .A2(new_n496), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n491), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT86), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n512), .A2(new_n513), .A3(new_n501), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n510), .A2(new_n514), .A3(new_n503), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT20), .ZN(new_n516));
  NOR2_X1   g330(.A1(G475), .A2(G902), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n516), .B1(new_n515), .B2(new_n517), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n506), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR3_X1   g335(.A1(new_n187), .A2(new_n407), .A3(G953), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n424), .A2(G122), .ZN(new_n524));
  INV_X1    g338(.A(G122), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(G116), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n524), .A2(new_n526), .A3(new_n190), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n205), .A2(G128), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n209), .A2(G143), .ZN(new_n529));
  AND3_X1   g343(.A1(new_n528), .A2(new_n529), .A3(new_n219), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n219), .B1(new_n528), .B2(new_n529), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n527), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(KEYINPUT14), .B1(new_n525), .B2(G116), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n525), .A2(G116), .ZN(new_n534));
  OAI21_X1  g348(.A(KEYINPUT89), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT14), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n536), .B1(new_n424), .B2(G122), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT89), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n537), .A2(new_n538), .A3(new_n524), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT90), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n540), .B1(new_n524), .B2(KEYINPUT14), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n534), .A2(KEYINPUT90), .A3(new_n536), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n535), .A2(new_n539), .A3(new_n541), .A4(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n532), .B1(G107), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n528), .A2(new_n529), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT13), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n529), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n545), .A2(new_n547), .A3(G134), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n528), .B(new_n529), .C1(new_n546), .C2(new_n219), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT88), .ZN(new_n551));
  INV_X1    g365(.A(new_n527), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n190), .B1(new_n524), .B2(new_n526), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n524), .A2(new_n526), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(G107), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n556), .A2(KEYINPUT88), .A3(new_n527), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n550), .B1(new_n554), .B2(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n523), .B1(new_n544), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n543), .A2(G107), .ZN(new_n560));
  INV_X1    g374(.A(new_n532), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AND2_X1   g376(.A1(new_n548), .A2(new_n549), .ZN(new_n563));
  NOR3_X1   g377(.A1(new_n552), .A2(new_n553), .A3(new_n551), .ZN(new_n564));
  AOI21_X1  g378(.A(KEYINPUT88), .B1(new_n556), .B2(new_n527), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n562), .A2(new_n566), .A3(new_n522), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n559), .A2(new_n567), .A3(KEYINPUT91), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n562), .A2(new_n566), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT91), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n569), .A2(new_n570), .A3(new_n523), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n568), .A2(new_n296), .A3(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(G478), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n573), .A2(KEYINPUT15), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n572), .B(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n521), .A2(new_n575), .ZN(new_n576));
  AND3_X1   g390(.A1(new_n468), .A2(new_n478), .A3(new_n576), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n302), .A2(new_n370), .A3(new_n416), .A4(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n578), .B(G101), .ZN(G3));
  NAND2_X1  g393(.A1(new_n348), .A2(new_n296), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(KEYINPUT92), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT92), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n348), .A2(new_n582), .A3(new_n296), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n581), .A2(G472), .A3(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n354), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n353), .B1(new_n348), .B2(new_n349), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n588), .A2(new_n415), .ZN(new_n589));
  AND2_X1   g403(.A1(new_n589), .A2(new_n302), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT33), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n568), .A2(new_n591), .A3(new_n571), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n573), .A2(G902), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT93), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n591), .B1(new_n569), .B2(new_n523), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n594), .B1(new_n595), .B2(new_n567), .ZN(new_n596));
  AND4_X1   g410(.A1(new_n594), .A2(new_n559), .A3(new_n567), .A4(KEYINPUT33), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n592), .B(new_n593), .C1(new_n596), .C2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT94), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n595), .A2(new_n594), .A3(new_n567), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n559), .A2(new_n567), .A3(KEYINPUT33), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(KEYINPUT93), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n604), .A2(KEYINPUT94), .A3(new_n592), .A4(new_n593), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n600), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(KEYINPUT95), .B(G478), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n572), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT96), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT97), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n606), .A2(new_n610), .A3(KEYINPUT97), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n521), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n468), .A2(new_n478), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n590), .A2(new_n618), .ZN(new_n619));
  XOR2_X1   g433(.A(KEYINPUT34), .B(G104), .Z(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G6));
  INV_X1    g435(.A(new_n575), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n515), .A2(new_n517), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(KEYINPUT20), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n624), .A2(KEYINPUT98), .A3(new_n518), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n625), .B(new_n506), .C1(KEYINPUT98), .C2(new_n518), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n617), .A2(new_n622), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n590), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT35), .B(G107), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G9));
  AND2_X1   g444(.A1(new_n302), .A2(new_n577), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT36), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n399), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(new_n395), .B(new_n633), .Z(new_n634));
  AOI22_X1  g448(.A1(new_n406), .A2(new_n408), .B1(new_n413), .B2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n588), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n631), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT37), .B(G110), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G12));
  XOR2_X1   g453(.A(KEYINPUT99), .B(G900), .Z(new_n640));
  NAND2_X1  g454(.A1(new_n475), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n473), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n626), .A2(new_n622), .A3(new_n643), .ZN(new_n644));
  AND2_X1   g458(.A1(new_n644), .A2(new_n468), .ZN(new_n645));
  INV_X1    g459(.A(new_n635), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n645), .A2(new_n302), .A3(new_n370), .A4(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G128), .ZN(G30));
  INV_X1    g462(.A(new_n369), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n649), .B1(new_n587), .B2(new_n352), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n356), .A2(new_n334), .ZN(new_n651));
  INV_X1    g465(.A(new_n362), .ZN(new_n652));
  OAI211_X1 g466(.A(new_n651), .B(new_n296), .C1(new_n652), .C2(new_n334), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(G472), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n656), .A2(new_n646), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n642), .B(KEYINPUT39), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n302), .A2(new_n658), .ZN(new_n659));
  OR2_X1    g473(.A1(new_n659), .A2(KEYINPUT40), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(KEYINPUT40), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n464), .A2(new_n467), .ZN(new_n662));
  XNOR2_X1  g476(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n464), .A2(new_n467), .A3(new_n663), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n521), .A2(new_n575), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n667), .A2(new_n418), .A3(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n657), .A2(new_n660), .A3(new_n661), .A4(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G143), .ZN(G45));
  AND3_X1   g485(.A1(new_n606), .A2(KEYINPUT97), .A3(new_n610), .ZN(new_n672));
  AOI21_X1  g486(.A(KEYINPUT97), .B1(new_n606), .B2(new_n610), .ZN(new_n673));
  OAI211_X1 g487(.A(new_n521), .B(new_n642), .C1(new_n672), .C2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT101), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n615), .A2(KEYINPUT101), .A3(new_n521), .A4(new_n642), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n676), .A2(new_n677), .A3(new_n468), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(KEYINPUT102), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n297), .A2(new_n301), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n370), .A2(new_n680), .A3(new_n188), .A4(new_n646), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT102), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n676), .A2(new_n677), .A3(new_n683), .A4(new_n468), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n679), .A2(new_n682), .A3(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT103), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n681), .B1(KEYINPUT102), .B2(new_n678), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n688), .A2(KEYINPUT103), .A3(new_n684), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G146), .ZN(G48));
  AND2_X1   g505(.A1(new_n370), .A2(new_n416), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n295), .B1(new_n294), .B2(new_n296), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n693), .A2(new_n694), .A3(new_n189), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n692), .A2(new_n618), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(KEYINPUT41), .B(G113), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G15));
  NAND3_X1  g512(.A1(new_n692), .A2(new_n627), .A3(new_n695), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G116), .ZN(G18));
  AND3_X1   g514(.A1(new_n370), .A2(new_n577), .A3(new_n646), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n695), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G119), .ZN(G21));
  NAND2_X1  g517(.A1(new_n580), .A2(G472), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n652), .A2(KEYINPUT28), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n334), .B1(new_n705), .B2(new_n359), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n345), .A2(new_n347), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n349), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n704), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n709), .A2(new_n415), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n617), .A2(new_n668), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n695), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G122), .ZN(G24));
  NAND2_X1  g527(.A1(new_n695), .A2(new_n468), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n709), .A2(new_n635), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n676), .A2(new_n677), .A3(new_n715), .ZN(new_n716));
  OR2_X1    g530(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G125), .ZN(G27));
  AOI21_X1  g532(.A(KEYINPUT32), .B1(new_n348), .B2(new_n349), .ZN(new_n719));
  OAI21_X1  g533(.A(KEYINPUT104), .B1(new_n649), .B2(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n719), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT104), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n721), .A2(new_n722), .A3(new_n369), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n720), .A2(new_n723), .A3(new_n368), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n724), .A2(new_n676), .A3(new_n677), .A4(new_n416), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n464), .A2(new_n467), .A3(new_n417), .ZN(new_n726));
  AOI211_X1 g540(.A(new_n189), .B(new_n726), .C1(new_n297), .C2(new_n301), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  OAI21_X1  g542(.A(KEYINPUT42), .B1(new_n725), .B2(new_n728), .ZN(new_n729));
  AND2_X1   g543(.A1(new_n676), .A2(new_n677), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT42), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n730), .A2(new_n692), .A3(new_n731), .A4(new_n727), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(new_n230), .ZN(G33));
  NAND3_X1  g548(.A1(new_n692), .A2(new_n644), .A3(new_n727), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G134), .ZN(G36));
  INV_X1    g550(.A(new_n278), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n270), .A2(new_n273), .A3(new_n737), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n738), .B1(new_n737), .B2(new_n298), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT45), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n295), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n738), .B(KEYINPUT45), .C1(new_n737), .C2(new_n298), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(KEYINPUT105), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n299), .A2(new_n278), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT105), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n744), .A2(new_n745), .A3(KEYINPUT45), .A4(new_n738), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n741), .A2(new_n743), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(G469), .A2(G902), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT46), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n747), .A2(KEYINPUT46), .A3(new_n748), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n751), .A2(new_n297), .A3(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n753), .A2(new_n188), .A3(new_n658), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(KEYINPUT106), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n726), .B(KEYINPUT107), .ZN(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(new_n521), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n758), .B1(new_n672), .B2(new_n673), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(KEYINPUT43), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT43), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n615), .A2(new_n761), .A3(new_n758), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n760), .A2(new_n762), .A3(new_n588), .A4(new_n646), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n763), .A2(KEYINPUT44), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(KEYINPUT44), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n757), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n755), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G137), .ZN(G39));
  INV_X1    g582(.A(KEYINPUT47), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n693), .B1(new_n749), .B2(new_n750), .ZN(new_n770));
  AOI211_X1 g584(.A(new_n769), .B(new_n189), .C1(new_n770), .C2(new_n752), .ZN(new_n771));
  AOI21_X1  g585(.A(KEYINPUT47), .B1(new_n753), .B2(new_n188), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n730), .ZN(new_n775));
  NOR4_X1   g589(.A1(new_n775), .A2(new_n416), .A3(new_n370), .A4(new_n726), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G140), .ZN(G42));
  OR4_X1    g592(.A1(new_n415), .A2(new_n759), .A3(new_n189), .A4(new_n418), .ZN(new_n779));
  XOR2_X1   g593(.A(new_n779), .B(KEYINPUT108), .Z(new_n780));
  NOR2_X1   g594(.A1(new_n693), .A2(new_n694), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(KEYINPUT49), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n780), .A2(new_n656), .A3(new_n667), .A4(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n668), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n784), .A2(new_n468), .A3(new_n642), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n655), .A2(new_n302), .A3(new_n635), .A4(new_n785), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n786), .B(new_n647), .C1(new_n714), .C2(new_n716), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n787), .B1(new_n687), .B2(new_n689), .ZN(new_n788));
  OAI21_X1  g602(.A(KEYINPUT52), .B1(new_n788), .B2(KEYINPUT110), .ZN(new_n789));
  INV_X1    g603(.A(new_n787), .ZN(new_n790));
  AOI21_X1  g604(.A(KEYINPUT103), .B1(new_n688), .B2(new_n684), .ZN(new_n791));
  AND4_X1   g605(.A1(KEYINPUT103), .A2(new_n679), .A3(new_n682), .A4(new_n684), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n790), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT110), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n789), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n696), .A2(new_n637), .A3(new_n578), .A4(new_n712), .ZN(new_n798));
  INV_X1    g612(.A(new_n615), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n576), .B1(new_n799), .B2(new_n521), .ZN(new_n800));
  INV_X1    g614(.A(new_n617), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n589), .A2(new_n800), .A3(new_n302), .A4(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n699), .A2(new_n702), .A3(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n798), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT109), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n729), .A2(new_n732), .A3(new_n735), .ZN(new_n806));
  INV_X1    g620(.A(new_n709), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n676), .A2(new_n677), .A3(new_n807), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n626), .A2(new_n575), .A3(new_n643), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n370), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n811), .A2(new_n646), .A3(new_n727), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n804), .A2(new_n805), .A3(new_n806), .A4(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n370), .A2(new_n416), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n294), .A2(new_n296), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(G469), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n816), .A2(new_n188), .A3(new_n297), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  AOI22_X1  g632(.A1(new_n818), .A2(new_n627), .B1(new_n701), .B2(new_n695), .ZN(new_n819));
  AOI22_X1  g633(.A1(new_n818), .A2(new_n618), .B1(new_n631), .B2(new_n636), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n712), .A2(new_n578), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n819), .A2(new_n820), .A3(new_n821), .A4(new_n802), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n812), .A2(new_n729), .A3(new_n732), .A4(new_n735), .ZN(new_n823));
  OAI21_X1  g637(.A(KEYINPUT109), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(KEYINPUT53), .B1(new_n813), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n797), .A2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n793), .A2(new_n795), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n788), .A2(KEYINPUT52), .ZN(new_n829));
  AOI22_X1  g643(.A1(new_n828), .A2(new_n829), .B1(new_n813), .B2(new_n824), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n826), .B(KEYINPUT54), .C1(new_n827), .C2(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n760), .A2(new_n762), .A3(new_n710), .A4(new_n474), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n470), .B1(new_n714), .B2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n726), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n816), .A2(new_n188), .A3(new_n297), .A4(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n415), .A2(new_n473), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n836), .A2(new_n355), .A3(new_n369), .A4(new_n654), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n835), .A2(new_n837), .A3(new_n616), .ZN(new_n838));
  OR2_X1    g652(.A1(new_n833), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n760), .A2(new_n762), .A3(new_n474), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n724), .A2(new_n416), .ZN(new_n842));
  INV_X1    g656(.A(new_n835), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n844), .A2(KEYINPUT48), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n844), .A2(KEYINPUT48), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n839), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n832), .A2(new_n757), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n781), .A2(new_n189), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n850), .B1(new_n773), .B2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT51), .ZN(new_n853));
  INV_X1    g667(.A(new_n832), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n667), .A2(new_n418), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n817), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n854), .A2(KEYINPUT50), .A3(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT50), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n417), .B1(new_n665), .B2(new_n666), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n859), .A2(new_n816), .A3(new_n188), .A4(new_n297), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n858), .B1(new_n832), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n853), .B1(new_n857), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n799), .A2(new_n758), .ZN(new_n863));
  OR3_X1    g677(.A1(new_n835), .A2(new_n837), .A3(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n841), .A2(new_n715), .A3(new_n843), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT112), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(new_n715), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n840), .A2(new_n835), .A3(new_n868), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n835), .A2(new_n837), .A3(new_n863), .ZN(new_n870));
  OAI21_X1  g684(.A(KEYINPUT112), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n862), .A2(new_n867), .A3(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n848), .B1(new_n852), .B2(new_n872), .ZN(new_n873));
  XNOR2_X1  g687(.A(KEYINPUT111), .B(KEYINPUT51), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n747), .A2(KEYINPUT46), .A3(new_n748), .ZN(new_n876));
  AOI21_X1  g690(.A(KEYINPUT46), .B1(new_n747), .B2(new_n748), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n876), .A2(new_n877), .A3(new_n693), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n769), .B1(new_n878), .B2(new_n189), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n753), .A2(KEYINPUT47), .A3(new_n188), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n879), .A2(new_n880), .A3(new_n851), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(new_n849), .ZN(new_n882));
  AOI211_X1 g696(.A(new_n870), .B(new_n869), .C1(new_n857), .C2(new_n861), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n875), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n873), .A2(new_n884), .A3(KEYINPUT113), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT113), .ZN(new_n886));
  INV_X1    g700(.A(new_n883), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n874), .B1(new_n852), .B2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n833), .A2(new_n838), .ZN(new_n889));
  AND2_X1   g703(.A1(new_n844), .A2(KEYINPUT48), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n889), .B1(new_n890), .B2(new_n845), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n862), .A2(new_n867), .A3(new_n871), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n891), .B1(new_n892), .B2(new_n882), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n886), .B1(new_n888), .B2(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n885), .A2(new_n894), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n822), .A2(new_n823), .A3(new_n827), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n795), .B1(new_n793), .B2(new_n794), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n788), .A2(KEYINPUT110), .A3(KEYINPUT52), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT54), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n899), .B(new_n900), .C1(KEYINPUT53), .C2(new_n830), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n831), .A2(new_n895), .A3(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT114), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n831), .A2(new_n895), .A3(new_n901), .A4(KEYINPUT114), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n469), .A2(new_n276), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n783), .B1(new_n904), .B2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT115), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI211_X1 g724(.A(KEYINPUT115), .B(new_n783), .C1(new_n904), .C2(new_n907), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(G75));
  NOR2_X1   g726(.A1(new_n276), .A2(G952), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT56), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n899), .B1(new_n830), .B2(KEYINPUT53), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(G902), .ZN(new_n917));
  INV_X1    g731(.A(G210), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n915), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n455), .A2(new_n459), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT116), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n921), .B(KEYINPUT55), .Z(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT117), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(new_n457), .Z(new_n924));
  OAI21_X1  g738(.A(new_n914), .B1(new_n919), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n919), .A2(new_n924), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT118), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n919), .A2(KEYINPUT118), .A3(new_n924), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n925), .B1(new_n928), .B2(new_n929), .ZN(G51));
  NAND2_X1  g744(.A1(new_n916), .A2(KEYINPUT54), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(new_n901), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n748), .B(KEYINPUT57), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n294), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n747), .B(KEYINPUT119), .Z(new_n936));
  NAND3_X1  g750(.A1(new_n916), .A2(G902), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n913), .B1(new_n935), .B2(new_n937), .ZN(G54));
  NAND4_X1  g752(.A1(new_n916), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n939));
  INV_X1    g753(.A(new_n515), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n939), .A2(new_n940), .ZN(new_n942));
  NOR3_X1   g756(.A1(new_n941), .A2(new_n942), .A3(new_n913), .ZN(G60));
  AND2_X1   g757(.A1(new_n604), .A2(new_n592), .ZN(new_n944));
  NAND2_X1  g758(.A1(G478), .A2(G902), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(KEYINPUT59), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n913), .B1(new_n932), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n831), .A2(new_n901), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n949), .A2(new_n946), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n948), .B1(new_n950), .B2(new_n944), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT120), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OAI211_X1 g767(.A(new_n948), .B(KEYINPUT120), .C1(new_n944), .C2(new_n950), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(G63));
  NAND2_X1  g769(.A1(G217), .A2(G902), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT60), .Z(new_n957));
  NAND3_X1  g771(.A1(new_n916), .A2(new_n634), .A3(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n410), .B1(new_n916), .B2(new_n957), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n959), .A2(new_n913), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(KEYINPUT61), .B1(new_n958), .B2(KEYINPUT121), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n961), .B(new_n962), .Z(G66));
  NOR3_X1   g777(.A1(new_n476), .A2(new_n433), .A3(new_n276), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n964), .B1(new_n804), .B2(new_n276), .ZN(new_n965));
  INV_X1    g779(.A(new_n921), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n966), .B1(G898), .B2(new_n276), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n965), .B(new_n967), .ZN(G69));
  NAND2_X1  g782(.A1(new_n340), .A2(new_n341), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(new_n507), .Z(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  AND2_X1   g785(.A1(new_n767), .A2(new_n777), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n717), .A2(new_n647), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n973), .B1(new_n687), .B2(new_n689), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(new_n670), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(KEYINPUT62), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n692), .A2(new_n834), .A3(new_n800), .ZN(new_n977));
  OR2_X1    g791(.A1(new_n977), .A2(new_n659), .ZN(new_n978));
  AND3_X1   g792(.A1(new_n972), .A2(new_n976), .A3(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT122), .ZN(new_n980));
  OR3_X1    g794(.A1(new_n975), .A2(new_n980), .A3(KEYINPUT62), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n980), .B1(new_n975), .B2(KEYINPUT62), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  AND2_X1   g797(.A1(new_n979), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n971), .B1(new_n984), .B2(G953), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n755), .A2(new_n468), .A3(new_n784), .A4(new_n842), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n974), .A2(new_n806), .ZN(new_n987));
  INV_X1    g801(.A(new_n987), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n972), .A2(new_n276), .A3(new_n986), .A4(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n971), .B1(G900), .B2(G953), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n985), .A2(new_n991), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT123), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n993), .B1(new_n989), .B2(new_n990), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n276), .B1(G227), .B2(G900), .ZN(new_n995));
  OAI21_X1  g809(.A(KEYINPUT124), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(new_n996), .ZN(new_n997));
  NOR3_X1   g811(.A1(new_n994), .A2(KEYINPUT124), .A3(new_n995), .ZN(new_n998));
  NOR3_X1   g812(.A1(new_n992), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(new_n998), .ZN(new_n1000));
  AOI22_X1  g814(.A1(new_n1000), .A2(new_n996), .B1(new_n985), .B2(new_n991), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n999), .A2(new_n1001), .ZN(G72));
  NAND3_X1  g816(.A1(new_n979), .A2(new_n983), .A3(new_n804), .ZN(new_n1003));
  XNOR2_X1  g817(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1004));
  AND2_X1   g818(.A1(G472), .A2(G902), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n1004), .B(new_n1005), .Z(new_n1006));
  INV_X1    g820(.A(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1003), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g822(.A(new_n651), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  OR2_X1    g824(.A1(new_n830), .A2(new_n827), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n356), .A2(new_n334), .ZN(new_n1012));
  NOR3_X1   g826(.A1(new_n1009), .A2(new_n1006), .A3(new_n1012), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n1011), .A2(new_n826), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g828(.A(KEYINPUT126), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g830(.A1(new_n1011), .A2(KEYINPUT126), .A3(new_n826), .A4(new_n1013), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n972), .A2(new_n986), .A3(new_n988), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1007), .B1(new_n1018), .B2(new_n822), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n913), .B1(new_n1019), .B2(new_n1012), .ZN(new_n1020));
  NAND4_X1  g834(.A1(new_n1010), .A2(new_n1016), .A3(new_n1017), .A4(new_n1020), .ZN(new_n1021));
  INV_X1    g835(.A(KEYINPUT127), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  AND2_X1   g837(.A1(new_n1020), .A2(new_n1017), .ZN(new_n1024));
  NAND4_X1  g838(.A1(new_n1024), .A2(KEYINPUT127), .A3(new_n1010), .A4(new_n1016), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1023), .A2(new_n1025), .ZN(G57));
endmodule


