//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 1 1 0 0 0 0 1 0 0 1 1 0 1 0 0 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 0 0 1 0 1 1 0 0 0 0 1 1 1 1 1 0 1 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n779,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n858, new_n860, new_n861, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n984, new_n985, new_n986, new_n987;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G64gat), .B(G92gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n202), .B(new_n203), .Z(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G226gat), .A2(G233gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT25), .ZN(new_n208));
  NAND2_X1  g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT24), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g010(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  NOR3_X1   g013(.A1(KEYINPUT64), .A2(G183gat), .A3(G190gat), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n211), .B(new_n212), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  AND2_X1   g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218));
  OR2_X1    g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT23), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(G176gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n220), .A2(G169gat), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n221), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n208), .B1(new_n217), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT66), .ZN(new_n227));
  NAND2_X1  g026(.A1(G169gat), .A2(G176gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(G169gat), .A2(G176gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n228), .B1(new_n229), .B2(KEYINPUT23), .ZN(new_n230));
  AND2_X1   g029(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n231));
  NOR2_X1   g030(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n230), .B1(new_n233), .B2(new_n223), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT25), .B1(new_n234), .B2(new_n216), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT66), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n208), .B1(new_n229), .B2(KEYINPUT23), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n211), .A2(new_n212), .ZN(new_n239));
  NOR2_X1   g038(.A1(G183gat), .A2(G190gat), .ZN(new_n240));
  OAI211_X1 g039(.A(new_n221), .B(new_n238), .C1(new_n239), .C2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n227), .A2(new_n237), .A3(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(KEYINPUT27), .B(G183gat), .ZN(new_n243));
  INV_X1    g042(.A(G190gat), .ZN(new_n244));
  AOI21_X1  g043(.A(KEYINPUT28), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n243), .A2(KEYINPUT28), .A3(new_n244), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT26), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n228), .B1(new_n229), .B2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT68), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  OAI211_X1 g051(.A(KEYINPUT68), .B(new_n228), .C1(new_n229), .C2(new_n249), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n229), .A2(new_n249), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n252), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n248), .A2(new_n255), .A3(new_n209), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n242), .A2(KEYINPUT78), .A3(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT78), .B1(new_n242), .B2(new_n256), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n207), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  AND2_X1   g059(.A1(G197gat), .A2(G204gat), .ZN(new_n261));
  NOR2_X1   g060(.A1(G197gat), .A2(G204gat), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT22), .ZN(new_n264));
  NAND2_X1  g063(.A1(G211gat), .A2(G218gat), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n266), .A2(KEYINPUT77), .ZN(new_n267));
  XOR2_X1   g066(.A(G211gat), .B(G218gat), .Z(new_n268));
  XNOR2_X1  g067(.A(new_n267), .B(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n241), .B1(new_n235), .B2(new_n236), .ZN(new_n271));
  AOI211_X1 g070(.A(KEYINPUT66), .B(KEYINPUT25), .C1(new_n234), .C2(new_n216), .ZN(new_n272));
  OAI21_X1  g071(.A(KEYINPUT67), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT67), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n227), .A2(new_n274), .A3(new_n237), .A4(new_n241), .ZN(new_n275));
  INV_X1    g074(.A(new_n247), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n209), .B1(new_n276), .B2(new_n245), .ZN(new_n277));
  INV_X1    g076(.A(new_n255), .ZN(new_n278));
  OAI21_X1  g077(.A(KEYINPUT69), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT69), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n248), .A2(new_n255), .A3(new_n280), .A4(new_n209), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n273), .A2(new_n275), .A3(new_n282), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n207), .A2(KEYINPUT29), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AND3_X1   g084(.A1(new_n260), .A2(new_n270), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n242), .A2(new_n256), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT78), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n289), .A2(new_n257), .A3(new_n284), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n273), .A2(new_n275), .A3(new_n207), .A4(new_n282), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n270), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n205), .B1(new_n286), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n290), .A2(new_n291), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(new_n269), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n260), .A2(new_n270), .A3(new_n285), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n295), .A2(new_n296), .A3(new_n204), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n293), .A2(KEYINPUT30), .A3(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT30), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n295), .A2(new_n299), .A3(new_n296), .A4(new_n204), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(G225gat), .A2(G233gat), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT72), .ZN(new_n304));
  INV_X1    g103(.A(G127gat), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n305), .A2(KEYINPUT70), .A3(G134gat), .ZN(new_n306));
  INV_X1    g105(.A(G134gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(G127gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(KEYINPUT70), .B(KEYINPUT71), .ZN(new_n310));
  XNOR2_X1  g109(.A(G113gat), .B(G120gat), .ZN(new_n311));
  OAI22_X1  g110(.A1(new_n309), .A2(new_n310), .B1(new_n311), .B2(KEYINPUT1), .ZN(new_n312));
  AND2_X1   g111(.A1(new_n309), .A2(new_n310), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n304), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  XOR2_X1   g113(.A(G113gat), .B(G120gat), .Z(new_n315));
  INV_X1    g114(.A(KEYINPUT1), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT71), .ZN(new_n318));
  AND2_X1   g117(.A1(new_n318), .A2(KEYINPUT70), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n318), .A2(KEYINPUT70), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n308), .B(new_n306), .C1(new_n319), .C2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n309), .A2(new_n310), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n317), .A2(new_n321), .A3(new_n322), .A4(KEYINPUT72), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n314), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n308), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n307), .A2(G127gat), .ZN(new_n326));
  NOR3_X1   g125(.A1(new_n317), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n324), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(G141gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(G148gat), .ZN(new_n331));
  OR2_X1    g130(.A1(new_n331), .A2(KEYINPUT79), .ZN(new_n332));
  XNOR2_X1  g131(.A(G155gat), .B(G162gat), .ZN(new_n333));
  INV_X1    g132(.A(G148gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(G141gat), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n331), .A2(new_n335), .A3(KEYINPUT79), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n332), .A2(new_n333), .A3(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(KEYINPUT80), .B(G162gat), .ZN(new_n339));
  INV_X1    g138(.A(G155gat), .ZN(new_n340));
  OAI21_X1  g139(.A(KEYINPUT2), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n331), .A2(new_n335), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT2), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n333), .ZN(new_n345));
  AOI22_X1  g144(.A1(new_n338), .A2(new_n341), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT3), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n344), .A2(new_n345), .ZN(new_n349));
  INV_X1    g148(.A(new_n341), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n349), .B1(new_n350), .B2(new_n337), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(KEYINPUT3), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n329), .A2(new_n348), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n327), .B1(new_n314), .B2(new_n323), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT4), .ZN(new_n355));
  AND3_X1   g154(.A1(new_n354), .A2(new_n355), .A3(new_n346), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n355), .B1(new_n354), .B2(new_n346), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n303), .B(new_n353), .C1(new_n356), .C2(new_n357), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n358), .A2(KEYINPUT5), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n329), .A2(new_n351), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n354), .A2(new_n346), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n303), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT82), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT5), .ZN(new_n365));
  NOR3_X1   g164(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n303), .ZN(new_n367));
  AND3_X1   g166(.A1(new_n324), .A2(new_n328), .A3(new_n346), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n354), .A2(new_n346), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n367), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(KEYINPUT82), .B1(new_n370), .B2(KEYINPUT5), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n366), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n358), .A2(KEYINPUT81), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n362), .A2(KEYINPUT4), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n354), .A2(new_n355), .A3(new_n346), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT81), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n376), .A2(new_n377), .A3(new_n303), .A4(new_n353), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n373), .A2(new_n378), .ZN(new_n379));
  AND3_X1   g178(.A1(new_n372), .A2(KEYINPUT83), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT83), .B1(new_n372), .B2(new_n379), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n360), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(G1gat), .B(G29gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n383), .B(KEYINPUT0), .ZN(new_n384));
  XNOR2_X1  g183(.A(G57gat), .B(G85gat), .ZN(new_n385));
  XOR2_X1   g184(.A(new_n384), .B(new_n385), .Z(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n382), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT84), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT6), .ZN(new_n390));
  OAI211_X1 g189(.A(new_n360), .B(new_n386), .C1(new_n380), .C2(new_n381), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n388), .A2(new_n389), .A3(new_n390), .A4(new_n391), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n382), .B(new_n387), .C1(KEYINPUT84), .C2(KEYINPUT6), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n302), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT29), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n269), .B1(new_n395), .B2(new_n348), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n396), .B1(G228gat), .B2(G233gat), .ZN(new_n397));
  INV_X1    g196(.A(new_n266), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n268), .B1(new_n398), .B2(KEYINPUT85), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n399), .A2(KEYINPUT85), .A3(new_n398), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(new_n395), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n399), .B1(KEYINPUT85), .B2(new_n398), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n347), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(new_n351), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n397), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n269), .A2(new_n395), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n346), .B1(new_n406), .B2(new_n347), .ZN(new_n407));
  OAI211_X1 g206(.A(G228gat), .B(G233gat), .C1(new_n407), .C2(new_n396), .ZN(new_n408));
  XNOR2_X1  g207(.A(KEYINPUT31), .B(G50gat), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  AND3_X1   g209(.A1(new_n405), .A2(new_n408), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n410), .B1(new_n405), .B2(new_n408), .ZN(new_n412));
  XNOR2_X1  g211(.A(G78gat), .B(G106gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n413), .B(G22gat), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  OR3_X1    g214(.A1(new_n411), .A2(new_n412), .A3(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n415), .B1(new_n411), .B2(new_n412), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n283), .A2(new_n354), .ZN(new_n419));
  INV_X1    g218(.A(G227gat), .ZN(new_n420));
  INV_X1    g219(.A(G233gat), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n273), .A2(new_n275), .A3(new_n329), .A4(new_n282), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n419), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT33), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(KEYINPUT73), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT73), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n424), .A2(new_n428), .A3(new_n425), .ZN(new_n429));
  XOR2_X1   g228(.A(G15gat), .B(G43gat), .Z(new_n430));
  XNOR2_X1  g229(.A(new_n430), .B(KEYINPUT74), .ZN(new_n431));
  XNOR2_X1  g230(.A(G71gat), .B(G99gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n431), .B(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n433), .B1(new_n424), .B2(KEYINPUT32), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n427), .A2(new_n429), .A3(new_n434), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n424), .B(KEYINPUT32), .C1(new_n425), .C2(new_n433), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n422), .B1(new_n419), .B2(new_n423), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n437), .B(KEYINPUT34), .ZN(new_n438));
  AND3_X1   g237(.A1(new_n435), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n438), .B1(new_n435), .B2(new_n436), .ZN(new_n440));
  NOR3_X1   g239(.A1(new_n418), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n394), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT35), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n416), .A2(new_n443), .A3(new_n417), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT90), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n445), .B1(new_n439), .B2(new_n440), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n435), .A2(new_n436), .ZN(new_n447));
  INV_X1    g246(.A(new_n438), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n435), .A2(new_n436), .A3(new_n438), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n449), .A2(KEYINPUT90), .A3(new_n450), .ZN(new_n451));
  AOI211_X1 g250(.A(new_n302), .B(new_n444), .C1(new_n446), .C2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT83), .ZN(new_n453));
  AND2_X1   g252(.A1(new_n373), .A2(new_n378), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n364), .B1(new_n363), .B2(new_n365), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n370), .A2(KEYINPUT82), .A3(KEYINPUT5), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n453), .B1(new_n454), .B2(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n372), .A2(KEYINPUT83), .A3(new_n379), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n359), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT6), .B1(new_n460), .B2(new_n386), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n387), .B1(new_n460), .B2(KEYINPUT87), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT87), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n382), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n461), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n460), .A2(new_n386), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT6), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  AOI22_X1  g267(.A1(KEYINPUT35), .A2(new_n442), .B1(new_n452), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT76), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n470), .B1(new_n439), .B2(new_n440), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT75), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n472), .B1(new_n439), .B2(new_n440), .ZN(new_n473));
  AOI22_X1  g272(.A1(KEYINPUT75), .A2(new_n471), .B1(new_n473), .B2(KEYINPUT36), .ZN(new_n474));
  AND3_X1   g273(.A1(new_n471), .A2(KEYINPUT75), .A3(KEYINPUT36), .ZN(new_n475));
  INV_X1    g274(.A(new_n418), .ZN(new_n476));
  OAI22_X1  g275(.A1(new_n474), .A2(new_n475), .B1(new_n394), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT89), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT37), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n295), .A2(new_n479), .A3(new_n296), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n294), .A2(new_n270), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n260), .A2(new_n269), .A3(new_n285), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n481), .A2(KEYINPUT37), .A3(new_n482), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n204), .A2(KEYINPUT38), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n480), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(new_n297), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT88), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n479), .B1(new_n295), .B2(new_n296), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n487), .B1(new_n488), .B2(new_n204), .ZN(new_n489));
  OAI21_X1  g288(.A(KEYINPUT37), .B1(new_n286), .B2(new_n292), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n490), .A2(KEYINPUT88), .A3(new_n205), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n489), .A2(new_n491), .A3(new_n480), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n486), .B1(new_n492), .B2(KEYINPUT38), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n465), .A2(new_n467), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n376), .A2(new_n353), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(new_n367), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n361), .A2(new_n303), .A3(new_n362), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n496), .A2(KEYINPUT39), .A3(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT39), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n495), .A2(new_n499), .A3(new_n367), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n500), .A2(KEYINPUT86), .A3(new_n386), .ZN(new_n501));
  AOI21_X1  g300(.A(KEYINPUT86), .B1(new_n500), .B2(new_n386), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n498), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT40), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT40), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n505), .B(new_n498), .C1(new_n501), .C2(new_n502), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n301), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n382), .A2(new_n463), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n460), .A2(KEYINPUT87), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n508), .A2(new_n509), .A3(new_n387), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n418), .B1(new_n507), .B2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n478), .B1(new_n494), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n477), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n494), .A2(new_n511), .A3(new_n478), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n469), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(G43gat), .ZN(new_n516));
  OAI21_X1  g315(.A(KEYINPUT15), .B1(new_n516), .B2(G50gat), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n517), .B1(new_n516), .B2(G50gat), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT94), .ZN(new_n519));
  INV_X1    g318(.A(G29gat), .ZN(new_n520));
  INV_X1    g319(.A(G36gat), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(KEYINPUT94), .A2(G29gat), .A3(G36gat), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n518), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g323(.A1(G29gat), .A2(G36gat), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT14), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n525), .B1(KEYINPUT91), .B2(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(KEYINPUT91), .B(KEYINPUT14), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n527), .B1(new_n528), .B2(new_n525), .ZN(new_n529));
  XNOR2_X1  g328(.A(KEYINPUT92), .B(KEYINPUT15), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT93), .ZN(new_n531));
  INV_X1    g330(.A(G50gat), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n531), .B1(new_n532), .B2(G43gat), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n533), .B1(new_n516), .B2(G50gat), .ZN(new_n534));
  NOR3_X1   g333(.A1(new_n531), .A2(new_n532), .A3(G43gat), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n530), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n524), .A2(new_n529), .A3(new_n536), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n529), .B1(new_n520), .B2(new_n521), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(new_n518), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT17), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(G15gat), .B(G22gat), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT16), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n543), .B1(new_n544), .B2(G1gat), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n545), .B1(G1gat), .B2(new_n543), .ZN(new_n546));
  INV_X1    g345(.A(G8gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n542), .A2(new_n549), .ZN(new_n550));
  AND3_X1   g349(.A1(new_n540), .A2(KEYINPUT95), .A3(new_n541), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT95), .B1(new_n540), .B2(new_n541), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(G229gat), .A2(G233gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n549), .A2(new_n540), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT18), .ZN(new_n557));
  AOI21_X1  g356(.A(KEYINPUT98), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(G113gat), .B(G141gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(G197gat), .ZN(new_n560));
  XOR2_X1   g359(.A(KEYINPUT11), .B(G169gat), .Z(new_n561));
  XNOR2_X1  g360(.A(new_n560), .B(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(KEYINPUT12), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n558), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n556), .A2(new_n557), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT96), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n555), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n549), .A2(KEYINPUT96), .A3(new_n540), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n548), .A2(new_n539), .A3(new_n537), .ZN(new_n569));
  AND2_X1   g368(.A1(new_n569), .A2(KEYINPUT97), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n569), .A2(KEYINPUT97), .ZN(new_n571));
  OAI211_X1 g370(.A(new_n567), .B(new_n568), .C1(new_n570), .C2(new_n571), .ZN(new_n572));
  XOR2_X1   g371(.A(new_n554), .B(KEYINPUT13), .Z(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n553), .A2(KEYINPUT18), .A3(new_n554), .A4(new_n555), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n565), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n564), .A2(new_n576), .ZN(new_n577));
  AOI22_X1  g376(.A1(new_n556), .A2(new_n557), .B1(new_n572), .B2(new_n573), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n578), .B(new_n575), .C1(new_n558), .C2(new_n563), .ZN(new_n579));
  AND2_X1   g378(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n551), .A2(new_n552), .ZN(new_n581));
  NAND2_X1  g380(.A1(G85gat), .A2(G92gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT7), .ZN(new_n583));
  NAND2_X1  g382(.A1(G99gat), .A2(G106gat), .ZN(new_n584));
  INV_X1    g383(.A(G85gat), .ZN(new_n585));
  INV_X1    g384(.A(G92gat), .ZN(new_n586));
  AOI22_X1  g385(.A1(KEYINPUT8), .A2(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(KEYINPUT102), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT102), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n583), .A2(new_n590), .A3(new_n587), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G99gat), .B(G106gat), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n593), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n589), .A2(new_n595), .A3(new_n591), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NOR3_X1   g396(.A1(new_n581), .A2(new_n542), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n540), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT41), .ZN(new_n600));
  NAND2_X1  g399(.A1(G232gat), .A2(G233gat), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  XOR2_X1   g402(.A(G190gat), .B(G218gat), .Z(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  XOR2_X1   g404(.A(G134gat), .B(G162gat), .Z(new_n606));
  NAND2_X1  g405(.A1(new_n601), .A2(new_n600), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n605), .B(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G120gat), .B(G148gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(G176gat), .B(G204gat), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n610), .B(new_n611), .Z(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT104), .ZN(new_n613));
  OAI21_X1  g412(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n614), .B1(G57gat), .B2(G64gat), .ZN(new_n615));
  INV_X1    g414(.A(G71gat), .ZN(new_n616));
  INV_X1    g415(.A(G78gat), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(G71gat), .A2(G78gat), .ZN(new_n619));
  OR3_X1    g418(.A1(new_n615), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(KEYINPUT99), .A2(G57gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(G64gat), .ZN(new_n622));
  AND2_X1   g421(.A1(new_n619), .A2(KEYINPUT9), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n622), .B1(new_n618), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n597), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n594), .A2(new_n625), .A3(new_n596), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT10), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n597), .A2(KEYINPUT10), .A3(new_n626), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(G230gat), .A2(G233gat), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n633), .B1(new_n627), .B2(new_n628), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n613), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(KEYINPUT105), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT105), .ZN(new_n639));
  OAI211_X1 g438(.A(new_n639), .B(new_n613), .C1(new_n635), .C2(new_n636), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT103), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n630), .A2(new_n631), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n642), .B1(new_n643), .B2(new_n633), .ZN(new_n644));
  AOI211_X1 g443(.A(KEYINPUT103), .B(new_n634), .C1(new_n630), .C2(new_n631), .ZN(new_n645));
  INV_X1    g444(.A(new_n612), .ZN(new_n646));
  OR4_X1    g445(.A1(new_n644), .A2(new_n645), .A3(new_n636), .A4(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n641), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT21), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n625), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(G231gat), .A2(G233gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(G127gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(G183gat), .B(G211gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n548), .B1(new_n650), .B2(new_n625), .ZN(new_n657));
  XOR2_X1   g456(.A(KEYINPUT100), .B(KEYINPUT101), .Z(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(G155gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n659), .B(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  OR2_X1    g462(.A1(new_n656), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n656), .A2(new_n663), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n609), .A2(new_n649), .A3(new_n667), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n515), .A2(new_n580), .A3(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n391), .A2(new_n389), .A3(new_n390), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n670), .A2(new_n466), .ZN(new_n671));
  INV_X1    g470(.A(new_n393), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g473(.A(KEYINPUT106), .B(G1gat), .Z(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(G1324gat));
  INV_X1    g475(.A(KEYINPUT107), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT16), .B(G8gat), .Z(new_n678));
  NAND3_X1  g477(.A1(new_n669), .A2(new_n302), .A3(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT42), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n515), .A2(new_n580), .ZN(new_n682));
  INV_X1    g481(.A(new_n668), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(G8gat), .B1(new_n684), .B2(new_n301), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n685), .A2(new_n679), .ZN(new_n686));
  OAI211_X1 g485(.A(new_n677), .B(new_n681), .C1(new_n686), .C2(new_n680), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n680), .B1(new_n685), .B2(new_n679), .ZN(new_n688));
  INV_X1    g487(.A(new_n681), .ZN(new_n689));
  OAI21_X1  g488(.A(KEYINPUT107), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n687), .A2(new_n690), .ZN(G1325gat));
  INV_X1    g490(.A(new_n475), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n473), .A2(KEYINPUT36), .ZN(new_n693));
  AOI21_X1  g492(.A(KEYINPUT76), .B1(new_n449), .B2(new_n450), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n693), .B1(new_n472), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(G15gat), .B1(new_n684), .B2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(G15gat), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n446), .A2(new_n451), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n669), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n697), .A2(new_n700), .ZN(G1326gat));
  NAND2_X1  g500(.A1(new_n669), .A2(new_n418), .ZN(new_n702));
  XNOR2_X1  g501(.A(KEYINPUT43), .B(G22gat), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n702), .B(new_n703), .ZN(G1327gat));
  NAND2_X1  g503(.A1(new_n649), .A2(new_n666), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n705), .A2(new_n609), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(KEYINPUT108), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n682), .A2(new_n520), .A3(new_n673), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(KEYINPUT109), .B(KEYINPUT45), .ZN(new_n709));
  OR2_X1    g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n711), .B1(new_n515), .B2(new_n609), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n494), .A2(new_n511), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(KEYINPUT89), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n418), .B1(new_n673), .B2(new_n302), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n714), .A2(new_n514), .A3(new_n715), .A4(new_n696), .ZN(new_n716));
  INV_X1    g515(.A(new_n469), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n608), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n605), .B(new_n719), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n718), .A2(KEYINPUT44), .A3(new_n720), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n705), .A2(new_n580), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n712), .A2(new_n721), .A3(new_n673), .A4(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(G29gat), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n710), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT110), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n710), .A2(KEYINPUT110), .A3(new_n724), .A4(new_n725), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(G1328gat));
  NAND4_X1  g529(.A1(new_n682), .A2(new_n521), .A3(new_n302), .A4(new_n707), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(KEYINPUT46), .ZN(new_n732));
  AND2_X1   g531(.A1(new_n712), .A2(new_n721), .ZN(new_n733));
  AND3_X1   g532(.A1(new_n733), .A2(new_n302), .A3(new_n722), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n731), .A2(KEYINPUT46), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n735), .A2(KEYINPUT111), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n735), .A2(KEYINPUT111), .ZN(new_n737));
  OAI221_X1 g536(.A(new_n732), .B1(new_n734), .B2(new_n521), .C1(new_n736), .C2(new_n737), .ZN(G1329gat));
  NAND3_X1  g537(.A1(new_n682), .A2(new_n699), .A3(new_n707), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n516), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n696), .A2(new_n516), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n712), .A2(new_n721), .A3(new_n722), .A4(new_n741), .ZN(new_n742));
  XNOR2_X1  g541(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n740), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n744), .A2(KEYINPUT113), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n744), .A2(KEYINPUT113), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n740), .A2(new_n742), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(KEYINPUT47), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n745), .B1(new_n746), .B2(new_n748), .ZN(G1330gat));
  NAND4_X1  g548(.A1(new_n712), .A2(new_n721), .A3(new_n418), .A4(new_n722), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(G50gat), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n682), .A2(new_n532), .A3(new_n418), .A4(new_n707), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT48), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n753), .B(new_n754), .ZN(G1331gat));
  NAND2_X1  g554(.A1(new_n577), .A2(new_n579), .ZN(new_n756));
  NOR4_X1   g555(.A1(new_n720), .A2(new_n649), .A3(new_n756), .A4(new_n666), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n718), .A2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(new_n673), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g560(.A1(new_n758), .A2(new_n301), .ZN(new_n762));
  NOR2_X1   g561(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n763));
  AND2_X1   g562(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n762), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n765), .B1(new_n762), .B2(new_n763), .ZN(G1333gat));
  NOR2_X1   g565(.A1(new_n696), .A2(new_n616), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n759), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(KEYINPUT114), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT114), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n759), .A2(new_n770), .A3(new_n767), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(new_n699), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n616), .B1(new_n758), .B2(new_n773), .ZN(new_n774));
  XNOR2_X1  g573(.A(KEYINPUT115), .B(KEYINPUT50), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n772), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n775), .B1(new_n772), .B2(new_n774), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n776), .A2(new_n777), .ZN(G1334gat));
  NOR2_X1   g577(.A1(new_n758), .A2(new_n476), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(new_n617), .ZN(G1335gat));
  NOR3_X1   g579(.A1(new_n649), .A2(new_n667), .A3(new_n756), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n733), .A2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n673), .ZN(new_n783));
  OAI21_X1  g582(.A(G85gat), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n667), .A2(new_n756), .ZN(new_n785));
  INV_X1    g584(.A(new_n514), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n786), .A2(new_n477), .A3(new_n512), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n720), .B(new_n785), .C1(new_n787), .C2(new_n469), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT51), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n609), .B1(new_n716), .B2(new_n717), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n791), .A2(KEYINPUT51), .A3(new_n785), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n649), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n793), .A2(new_n585), .A3(new_n673), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n784), .A2(new_n794), .ZN(G1336gat));
  NAND4_X1  g594(.A1(new_n712), .A2(new_n721), .A3(new_n302), .A4(new_n781), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(G92gat), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n649), .A2(G92gat), .A3(new_n301), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n788), .A2(new_n789), .ZN(new_n799));
  AOI21_X1  g598(.A(KEYINPUT51), .B1(new_n791), .B2(new_n785), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n798), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n797), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(KEYINPUT52), .ZN(G1337gat));
  OAI21_X1  g602(.A(G99gat), .B1(new_n782), .B2(new_n696), .ZN(new_n804));
  INV_X1    g603(.A(G99gat), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n793), .A2(new_n805), .A3(new_n699), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(G1338gat));
  INV_X1    g606(.A(KEYINPUT117), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n476), .A2(G106gat), .ZN(new_n809));
  OAI211_X1 g608(.A(new_n648), .B(new_n809), .C1(new_n799), .C2(new_n800), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n712), .A2(new_n721), .A3(new_n418), .A4(new_n781), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(G106gat), .ZN(new_n812));
  XOR2_X1   g611(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n813));
  AND4_X1   g612(.A1(new_n808), .A2(new_n810), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  AOI22_X1  g613(.A1(new_n793), .A2(new_n809), .B1(new_n811), .B2(G106gat), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n808), .B1(new_n815), .B2(new_n813), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n810), .A2(new_n812), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(KEYINPUT53), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n814), .B1(new_n816), .B2(new_n818), .ZN(G1339gat));
  NAND3_X1  g618(.A1(new_n578), .A2(new_n563), .A3(new_n575), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n572), .A2(new_n573), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n554), .B1(new_n553), .B2(new_n555), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n562), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n824), .B1(new_n641), .B2(new_n647), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT54), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n643), .A2(new_n827), .A3(new_n633), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n646), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(KEYINPUT103), .B1(new_n632), .B2(new_n634), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n643), .A2(new_n642), .A3(new_n633), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n630), .A2(new_n631), .A3(new_n634), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(KEYINPUT54), .ZN(new_n835));
  OAI211_X1 g634(.A(KEYINPUT55), .B(new_n830), .C1(new_n833), .C2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT55), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n644), .A2(new_n645), .A3(new_n835), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n837), .B1(new_n838), .B2(new_n829), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n756), .A2(new_n647), .A3(new_n836), .A4(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n720), .B1(new_n826), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n839), .A2(new_n836), .A3(new_n647), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n609), .A2(new_n842), .A3(new_n824), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n666), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n668), .A2(new_n756), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n418), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n847), .A2(new_n673), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n439), .A2(new_n440), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n848), .A2(new_n301), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(G113gat), .B1(new_n850), .B2(new_n756), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n848), .A2(new_n301), .A3(new_n699), .ZN(new_n852));
  INV_X1    g651(.A(G113gat), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n852), .A2(new_n853), .A3(new_n580), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n851), .A2(new_n854), .ZN(G1340gat));
  AOI21_X1  g654(.A(G120gat), .B1(new_n850), .B2(new_n648), .ZN(new_n856));
  INV_X1    g655(.A(G120gat), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n852), .A2(new_n857), .A3(new_n649), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n856), .A2(new_n858), .ZN(G1341gat));
  NAND3_X1  g658(.A1(new_n850), .A2(new_n305), .A3(new_n667), .ZN(new_n860));
  OAI21_X1  g659(.A(G127gat), .B1(new_n852), .B2(new_n666), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(G1342gat));
  NOR2_X1   g661(.A1(new_n609), .A2(new_n302), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n848), .A2(new_n307), .A3(new_n849), .A4(new_n863), .ZN(new_n864));
  OR2_X1    g663(.A1(new_n864), .A2(KEYINPUT118), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(KEYINPUT118), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n865), .A2(KEYINPUT56), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(G134gat), .B1(new_n852), .B2(new_n609), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(KEYINPUT56), .B1(new_n865), .B2(new_n866), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n869), .A2(new_n870), .ZN(G1343gat));
  INV_X1    g670(.A(KEYINPUT58), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n476), .B1(new_n844), .B2(new_n846), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n783), .B1(new_n695), .B2(new_n692), .ZN(new_n874));
  AND3_X1   g673(.A1(new_n873), .A2(new_n301), .A3(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n875), .A2(new_n330), .A3(new_n756), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n874), .A2(new_n301), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT57), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n877), .B1(new_n878), .B2(new_n873), .ZN(new_n879));
  INV_X1    g678(.A(new_n843), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n580), .B1(KEYINPUT119), .B2(new_n842), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT119), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n839), .A2(new_n836), .A3(new_n882), .A4(new_n647), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n825), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n880), .B1(new_n884), .B2(new_n720), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n845), .B1(new_n885), .B2(new_n666), .ZN(new_n886));
  OAI21_X1  g685(.A(KEYINPUT57), .B1(new_n886), .B2(new_n476), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n879), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n756), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT120), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(G141gat), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n889), .A2(new_n890), .ZN(new_n893));
  OAI211_X1 g692(.A(new_n872), .B(new_n876), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n889), .A2(G141gat), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(new_n876), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(KEYINPUT58), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n894), .A2(new_n897), .ZN(G1344gat));
  INV_X1    g697(.A(KEYINPUT122), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n875), .A2(new_n334), .A3(new_n648), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT121), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n873), .A2(KEYINPUT57), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n842), .A2(KEYINPUT119), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n903), .A2(new_n756), .A3(new_n883), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n720), .B1(new_n904), .B2(new_n826), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n666), .B1(new_n905), .B2(new_n843), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n476), .B1(new_n906), .B2(new_n846), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n902), .B1(new_n907), .B2(KEYINPUT57), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n874), .A2(new_n301), .A3(new_n648), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n334), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT59), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n901), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n878), .B1(new_n886), .B2(new_n476), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n909), .B1(new_n914), .B2(new_n902), .ZN(new_n915));
  OAI211_X1 g714(.A(KEYINPUT121), .B(KEYINPUT59), .C1(new_n915), .C2(new_n334), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n913), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n888), .A2(new_n648), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n334), .A2(KEYINPUT59), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI211_X1 g719(.A(new_n899), .B(new_n900), .C1(new_n917), .C2(new_n920), .ZN(new_n921));
  AOI22_X1  g720(.A1(new_n913), .A2(new_n916), .B1(new_n918), .B2(new_n919), .ZN(new_n922));
  INV_X1    g721(.A(new_n900), .ZN(new_n923));
  OAI21_X1  g722(.A(KEYINPUT122), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n921), .A2(new_n924), .ZN(G1345gat));
  AOI21_X1  g724(.A(G155gat), .B1(new_n875), .B2(new_n667), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n667), .A2(G155gat), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n927), .B(KEYINPUT123), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n926), .B1(new_n888), .B2(new_n928), .ZN(G1346gat));
  NAND4_X1  g728(.A1(new_n873), .A2(new_n339), .A3(new_n863), .A4(new_n874), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n888), .A2(KEYINPUT124), .A3(new_n720), .ZN(new_n931));
  INV_X1    g730(.A(new_n339), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g732(.A(KEYINPUT124), .B1(new_n888), .B2(new_n720), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n930), .B1(new_n933), .B2(new_n934), .ZN(G1347gat));
  NAND2_X1  g734(.A1(new_n844), .A2(new_n846), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n673), .A2(new_n301), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n936), .A2(new_n441), .A3(new_n937), .ZN(new_n938));
  INV_X1    g737(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g738(.A(G169gat), .B1(new_n939), .B2(new_n756), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n847), .A2(new_n699), .A3(new_n937), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT125), .ZN(new_n942));
  OR2_X1    g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n941), .A2(new_n942), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AND2_X1   g744(.A1(new_n756), .A2(G169gat), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n940), .B1(new_n945), .B2(new_n946), .ZN(G1348gat));
  AOI21_X1  g746(.A(G176gat), .B1(new_n939), .B2(new_n648), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n649), .A2(new_n233), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n948), .B1(new_n945), .B2(new_n949), .ZN(G1349gat));
  NAND3_X1  g749(.A1(new_n943), .A2(new_n667), .A3(new_n944), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(G183gat), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n939), .A2(new_n243), .A3(new_n667), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n954), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g754(.A1(new_n939), .A2(new_n244), .A3(new_n720), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT61), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n945), .A2(new_n720), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n957), .B1(new_n958), .B2(G190gat), .ZN(new_n959));
  AOI211_X1 g758(.A(KEYINPUT61), .B(new_n244), .C1(new_n945), .C2(new_n720), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n956), .B1(new_n959), .B2(new_n960), .ZN(G1351gat));
  NAND2_X1  g760(.A1(new_n696), .A2(new_n937), .ZN(new_n962));
  INV_X1    g761(.A(new_n962), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(new_n873), .ZN(new_n964));
  INV_X1    g763(.A(new_n964), .ZN(new_n965));
  AOI21_X1  g764(.A(G197gat), .B1(new_n965), .B2(new_n756), .ZN(new_n966));
  XNOR2_X1  g765(.A(new_n962), .B(KEYINPUT126), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n908), .A2(new_n967), .ZN(new_n968));
  INV_X1    g767(.A(new_n968), .ZN(new_n969));
  AND2_X1   g768(.A1(new_n756), .A2(G197gat), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n966), .B1(new_n969), .B2(new_n970), .ZN(G1352gat));
  OAI21_X1  g770(.A(G204gat), .B1(new_n968), .B2(new_n649), .ZN(new_n972));
  NOR4_X1   g771(.A1(new_n673), .A2(G204gat), .A3(new_n301), .A4(new_n649), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n873), .A2(new_n696), .A3(new_n973), .ZN(new_n974));
  XOR2_X1   g773(.A(new_n974), .B(KEYINPUT62), .Z(new_n975));
  NAND2_X1  g774(.A1(new_n972), .A2(new_n975), .ZN(G1353gat));
  INV_X1    g775(.A(G211gat), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n963), .A2(new_n667), .ZN(new_n978));
  INV_X1    g777(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n977), .B1(new_n908), .B2(new_n979), .ZN(new_n980));
  XNOR2_X1  g779(.A(new_n980), .B(KEYINPUT63), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n965), .A2(new_n977), .A3(new_n667), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n981), .A2(new_n982), .ZN(G1354gat));
  INV_X1    g782(.A(G218gat), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n984), .B1(new_n964), .B2(new_n609), .ZN(new_n985));
  XNOR2_X1  g784(.A(new_n985), .B(KEYINPUT127), .ZN(new_n986));
  NOR3_X1   g785(.A1(new_n968), .A2(new_n984), .A3(new_n609), .ZN(new_n987));
  NOR2_X1   g786(.A1(new_n986), .A2(new_n987), .ZN(G1355gat));
endmodule


