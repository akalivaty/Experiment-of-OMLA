

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584;

  XOR2_X1 U322 ( .A(n442), .B(n441), .Z(n525) );
  NOR2_X1 U323 ( .A1(n380), .A2(n574), .ZN(n382) );
  XNOR2_X1 U324 ( .A(n483), .B(KEYINPUT99), .ZN(n484) );
  XOR2_X1 U325 ( .A(KEYINPUT121), .B(n444), .Z(n562) );
  XOR2_X1 U326 ( .A(n355), .B(n354), .Z(n561) );
  AND2_X1 U327 ( .A1(G228GAT), .A2(G233GAT), .ZN(n290) );
  AND2_X1 U328 ( .A1(n544), .A2(n547), .ZN(n341) );
  XNOR2_X1 U329 ( .A(n410), .B(n290), .ZN(n411) );
  INV_X1 U330 ( .A(KEYINPUT110), .ZN(n381) );
  XNOR2_X1 U331 ( .A(n346), .B(n329), .ZN(n330) );
  XNOR2_X1 U332 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U333 ( .A(n415), .B(KEYINPUT24), .ZN(n416) );
  XNOR2_X1 U334 ( .A(n422), .B(n330), .ZN(n335) );
  XNOR2_X1 U335 ( .A(n417), .B(n416), .ZN(n420) );
  NOR2_X1 U336 ( .A1(n540), .A2(n518), .ZN(n524) );
  XOR2_X1 U337 ( .A(n561), .B(KEYINPUT36), .Z(n582) );
  NOR2_X1 U338 ( .A1(n443), .A2(n454), .ZN(n444) );
  XNOR2_X1 U339 ( .A(n485), .B(n484), .ZN(n512) );
  XOR2_X1 U340 ( .A(KEYINPUT41), .B(n574), .Z(n547) );
  XNOR2_X1 U341 ( .A(n447), .B(G176GAT), .ZN(n448) );
  XNOR2_X1 U342 ( .A(n449), .B(n448), .ZN(G1349GAT) );
  XOR2_X1 U343 ( .A(G169GAT), .B(G8GAT), .Z(n309) );
  XOR2_X1 U344 ( .A(G36GAT), .B(G190GAT), .Z(n353) );
  XNOR2_X1 U345 ( .A(n309), .B(n353), .ZN(n304) );
  XOR2_X1 U346 ( .A(KEYINPUT90), .B(KEYINPUT88), .Z(n292) );
  NAND2_X1 U347 ( .A1(G226GAT), .A2(G233GAT), .ZN(n291) );
  XNOR2_X1 U348 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U349 ( .A(n293), .B(KEYINPUT89), .Z(n299) );
  XOR2_X1 U350 ( .A(G183GAT), .B(KEYINPUT18), .Z(n295) );
  XNOR2_X1 U351 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n294) );
  XNOR2_X1 U352 ( .A(n295), .B(n294), .ZN(n433) );
  XOR2_X1 U353 ( .A(G211GAT), .B(KEYINPUT21), .Z(n297) );
  XNOR2_X1 U354 ( .A(G197GAT), .B(G218GAT), .ZN(n296) );
  XNOR2_X1 U355 ( .A(n297), .B(n296), .ZN(n412) );
  XNOR2_X1 U356 ( .A(n433), .B(n412), .ZN(n298) );
  XNOR2_X1 U357 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U358 ( .A(G176GAT), .B(G64GAT), .Z(n331) );
  XOR2_X1 U359 ( .A(n300), .B(n331), .Z(n302) );
  XNOR2_X1 U360 ( .A(G204GAT), .B(G92GAT), .ZN(n301) );
  XNOR2_X1 U361 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U362 ( .A(n304), .B(n303), .Z(n515) );
  INV_X1 U363 ( .A(n515), .ZN(n387) );
  XOR2_X1 U364 ( .A(G1GAT), .B(G197GAT), .Z(n306) );
  XNOR2_X1 U365 ( .A(G113GAT), .B(G15GAT), .ZN(n305) );
  XNOR2_X1 U366 ( .A(n306), .B(n305), .ZN(n322) );
  XOR2_X1 U367 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n308) );
  XNOR2_X1 U368 ( .A(KEYINPUT67), .B(KEYINPUT66), .ZN(n307) );
  XNOR2_X1 U369 ( .A(n308), .B(n307), .ZN(n313) );
  XOR2_X1 U370 ( .A(G50GAT), .B(G36GAT), .Z(n311) );
  XOR2_X1 U371 ( .A(G141GAT), .B(G22GAT), .Z(n418) );
  XNOR2_X1 U372 ( .A(n418), .B(n309), .ZN(n310) );
  XNOR2_X1 U373 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U374 ( .A(n313), .B(n312), .Z(n315) );
  NAND2_X1 U375 ( .A1(G229GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U376 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U377 ( .A(n316), .B(KEYINPUT68), .Z(n320) );
  XOR2_X1 U378 ( .A(G29GAT), .B(G43GAT), .Z(n318) );
  XNOR2_X1 U379 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n317) );
  XNOR2_X1 U380 ( .A(n318), .B(n317), .ZN(n345) );
  XNOR2_X1 U381 ( .A(n345), .B(KEYINPUT69), .ZN(n319) );
  XNOR2_X1 U382 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U383 ( .A(n322), .B(n321), .ZN(n571) );
  INV_X1 U384 ( .A(n571), .ZN(n544) );
  XNOR2_X1 U385 ( .A(G148GAT), .B(KEYINPUT71), .ZN(n323) );
  XNOR2_X1 U386 ( .A(n323), .B(KEYINPUT72), .ZN(n324) );
  XOR2_X1 U387 ( .A(n324), .B(G204GAT), .Z(n326) );
  XNOR2_X1 U388 ( .A(G78GAT), .B(G106GAT), .ZN(n325) );
  XNOR2_X1 U389 ( .A(n326), .B(n325), .ZN(n422) );
  XOR2_X1 U390 ( .A(KEYINPUT73), .B(G92GAT), .Z(n328) );
  XNOR2_X1 U391 ( .A(G99GAT), .B(G85GAT), .ZN(n327) );
  XNOR2_X1 U392 ( .A(n328), .B(n327), .ZN(n346) );
  XOR2_X1 U393 ( .A(KEYINPUT75), .B(KEYINPUT31), .Z(n329) );
  XOR2_X1 U394 ( .A(G57GAT), .B(KEYINPUT13), .Z(n362) );
  XOR2_X1 U395 ( .A(n362), .B(n331), .Z(n333) );
  NAND2_X1 U396 ( .A1(G230GAT), .A2(G233GAT), .ZN(n332) );
  XOR2_X1 U397 ( .A(n333), .B(n332), .Z(n334) );
  XNOR2_X1 U398 ( .A(n335), .B(n334), .ZN(n340) );
  XOR2_X1 U399 ( .A(G120GAT), .B(G71GAT), .Z(n429) );
  XOR2_X1 U400 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n337) );
  XNOR2_X1 U401 ( .A(KEYINPUT70), .B(KEYINPUT74), .ZN(n336) );
  XNOR2_X1 U402 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U403 ( .A(n429), .B(n338), .ZN(n339) );
  XNOR2_X1 U404 ( .A(n340), .B(n339), .ZN(n574) );
  XNOR2_X1 U405 ( .A(n341), .B(KEYINPUT46), .ZN(n356) );
  XOR2_X1 U406 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n343) );
  NAND2_X1 U407 ( .A1(G232GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U408 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U409 ( .A(n344), .B(KEYINPUT9), .Z(n348) );
  XNOR2_X1 U410 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U411 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U412 ( .A(KEYINPUT64), .B(G218GAT), .Z(n350) );
  XNOR2_X1 U413 ( .A(G134GAT), .B(G106GAT), .ZN(n349) );
  XNOR2_X1 U414 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U415 ( .A(n352), .B(n351), .Z(n355) );
  XOR2_X1 U416 ( .A(G50GAT), .B(G162GAT), .Z(n410) );
  XNOR2_X1 U417 ( .A(n410), .B(n353), .ZN(n354) );
  NOR2_X1 U418 ( .A1(n356), .A2(n561), .ZN(n375) );
  XOR2_X1 U419 ( .A(G211GAT), .B(G78GAT), .Z(n358) );
  XNOR2_X1 U420 ( .A(G1GAT), .B(G8GAT), .ZN(n357) );
  XNOR2_X1 U421 ( .A(n358), .B(n357), .ZN(n374) );
  XOR2_X1 U422 ( .A(KEYINPUT79), .B(KEYINPUT78), .Z(n360) );
  NAND2_X1 U423 ( .A1(G231GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U424 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U425 ( .A(KEYINPUT12), .B(n361), .ZN(n372) );
  XOR2_X1 U426 ( .A(G15GAT), .B(G127GAT), .Z(n428) );
  XOR2_X1 U427 ( .A(n362), .B(n428), .Z(n364) );
  XNOR2_X1 U428 ( .A(G183GAT), .B(G71GAT), .ZN(n363) );
  XNOR2_X1 U429 ( .A(n364), .B(n363), .ZN(n368) );
  XOR2_X1 U430 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n366) );
  XNOR2_X1 U431 ( .A(G64GAT), .B(KEYINPUT77), .ZN(n365) );
  XNOR2_X1 U432 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U433 ( .A(n368), .B(n367), .Z(n370) );
  XNOR2_X1 U434 ( .A(G22GAT), .B(G155GAT), .ZN(n369) );
  XNOR2_X1 U435 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U436 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U437 ( .A(n374), .B(n373), .Z(n531) );
  NAND2_X1 U438 ( .A1(n375), .A2(n531), .ZN(n377) );
  XOR2_X1 U439 ( .A(KEYINPUT47), .B(KEYINPUT109), .Z(n376) );
  XNOR2_X1 U440 ( .A(n377), .B(n376), .ZN(n385) );
  NOR2_X1 U441 ( .A1(n531), .A2(n582), .ZN(n379) );
  XNOR2_X1 U442 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n378) );
  XNOR2_X1 U443 ( .A(n379), .B(n378), .ZN(n380) );
  NOR2_X1 U444 ( .A1(n544), .A2(n383), .ZN(n384) );
  NOR2_X1 U445 ( .A1(n385), .A2(n384), .ZN(n386) );
  XNOR2_X1 U446 ( .A(n386), .B(KEYINPUT48), .ZN(n541) );
  NOR2_X1 U447 ( .A1(n387), .A2(n541), .ZN(n388) );
  XNOR2_X1 U448 ( .A(n388), .B(KEYINPUT54), .ZN(n567) );
  XOR2_X1 U449 ( .A(KEYINPUT87), .B(G148GAT), .Z(n390) );
  XNOR2_X1 U450 ( .A(G141GAT), .B(G127GAT), .ZN(n389) );
  XNOR2_X1 U451 ( .A(n390), .B(n389), .ZN(n394) );
  XOR2_X1 U452 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n392) );
  XNOR2_X1 U453 ( .A(KEYINPUT4), .B(KEYINPUT5), .ZN(n391) );
  XNOR2_X1 U454 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U455 ( .A(n394), .B(n393), .Z(n399) );
  XOR2_X1 U456 ( .A(KEYINPUT86), .B(G57GAT), .Z(n396) );
  NAND2_X1 U457 ( .A1(G225GAT), .A2(G233GAT), .ZN(n395) );
  XNOR2_X1 U458 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U459 ( .A(G1GAT), .B(n397), .ZN(n398) );
  XNOR2_X1 U460 ( .A(n399), .B(n398), .ZN(n404) );
  XOR2_X1 U461 ( .A(G85GAT), .B(G162GAT), .Z(n402) );
  XNOR2_X1 U462 ( .A(G155GAT), .B(KEYINPUT2), .ZN(n400) );
  XNOR2_X1 U463 ( .A(n400), .B(KEYINPUT3), .ZN(n414) );
  XNOR2_X1 U464 ( .A(G29GAT), .B(n414), .ZN(n401) );
  XNOR2_X1 U465 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U466 ( .A(n404), .B(n403), .Z(n409) );
  XOR2_X1 U467 ( .A(KEYINPUT0), .B(G134GAT), .Z(n406) );
  XNOR2_X1 U468 ( .A(KEYINPUT80), .B(KEYINPUT81), .ZN(n405) );
  XNOR2_X1 U469 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U470 ( .A(G113GAT), .B(n407), .ZN(n441) );
  XOR2_X1 U471 ( .A(n441), .B(G120GAT), .Z(n408) );
  XOR2_X1 U472 ( .A(n409), .B(n408), .Z(n568) );
  XNOR2_X1 U473 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U474 ( .A(n413), .B(KEYINPUT22), .Z(n417) );
  XNOR2_X1 U475 ( .A(KEYINPUT85), .B(n414), .ZN(n415) );
  XOR2_X1 U476 ( .A(n418), .B(KEYINPUT23), .Z(n419) );
  XNOR2_X1 U477 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U478 ( .A(n422), .B(n421), .ZN(n460) );
  AND2_X1 U479 ( .A1(n568), .A2(n460), .ZN(n423) );
  NAND2_X1 U480 ( .A1(n567), .A2(n423), .ZN(n425) );
  XOR2_X1 U481 ( .A(KEYINPUT55), .B(KEYINPUT120), .Z(n424) );
  XNOR2_X1 U482 ( .A(n425), .B(n424), .ZN(n443) );
  XOR2_X1 U483 ( .A(KEYINPUT83), .B(KEYINPUT82), .Z(n427) );
  XNOR2_X1 U484 ( .A(G169GAT), .B(G176GAT), .ZN(n426) );
  XNOR2_X1 U485 ( .A(n427), .B(n426), .ZN(n440) );
  XOR2_X1 U486 ( .A(KEYINPUT84), .B(G190GAT), .Z(n431) );
  XNOR2_X1 U487 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U488 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U489 ( .A(n432), .B(G99GAT), .Z(n438) );
  XOR2_X1 U490 ( .A(n433), .B(KEYINPUT20), .Z(n435) );
  NAND2_X1 U491 ( .A1(G227GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U492 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U493 ( .A(G43GAT), .B(n436), .ZN(n437) );
  XNOR2_X1 U494 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U495 ( .A(n440), .B(n439), .ZN(n442) );
  INV_X1 U496 ( .A(n525), .ZN(n454) );
  NAND2_X1 U497 ( .A1(n562), .A2(n544), .ZN(n446) );
  XNOR2_X1 U498 ( .A(G169GAT), .B(KEYINPUT122), .ZN(n445) );
  XNOR2_X1 U499 ( .A(n446), .B(n445), .ZN(G1348GAT) );
  NAND2_X1 U500 ( .A1(n562), .A2(n547), .ZN(n449) );
  XOR2_X1 U501 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n447) );
  XOR2_X1 U502 ( .A(KEYINPUT34), .B(KEYINPUT96), .Z(n472) );
  NOR2_X1 U503 ( .A1(n574), .A2(n571), .ZN(n450) );
  XOR2_X1 U504 ( .A(KEYINPUT76), .B(n450), .Z(n486) );
  NOR2_X1 U505 ( .A1(n531), .A2(n561), .ZN(n451) );
  XNOR2_X1 U506 ( .A(n451), .B(KEYINPUT16), .ZN(n469) );
  INV_X1 U507 ( .A(n568), .ZN(n513) );
  XNOR2_X1 U508 ( .A(n515), .B(KEYINPUT27), .ZN(n459) );
  NAND2_X1 U509 ( .A1(n513), .A2(n459), .ZN(n540) );
  INV_X1 U510 ( .A(KEYINPUT28), .ZN(n452) );
  XNOR2_X1 U511 ( .A(n452), .B(n460), .ZN(n518) );
  INV_X1 U512 ( .A(KEYINPUT91), .ZN(n453) );
  XNOR2_X1 U513 ( .A(n524), .B(n453), .ZN(n455) );
  NAND2_X1 U514 ( .A1(n455), .A2(n454), .ZN(n456) );
  XNOR2_X1 U515 ( .A(n456), .B(KEYINPUT92), .ZN(n468) );
  NOR2_X1 U516 ( .A1(n525), .A2(n460), .ZN(n457) );
  XOR2_X1 U517 ( .A(KEYINPUT93), .B(n457), .Z(n458) );
  XNOR2_X1 U518 ( .A(KEYINPUT26), .B(n458), .ZN(n569) );
  NAND2_X1 U519 ( .A1(n569), .A2(n459), .ZN(n465) );
  NAND2_X1 U520 ( .A1(n515), .A2(n525), .ZN(n461) );
  NAND2_X1 U521 ( .A1(n461), .A2(n460), .ZN(n462) );
  XNOR2_X1 U522 ( .A(n462), .B(KEYINPUT94), .ZN(n463) );
  XOR2_X1 U523 ( .A(KEYINPUT25), .B(n463), .Z(n464) );
  NAND2_X1 U524 ( .A1(n465), .A2(n464), .ZN(n466) );
  NAND2_X1 U525 ( .A1(n466), .A2(n568), .ZN(n467) );
  NAND2_X1 U526 ( .A1(n468), .A2(n467), .ZN(n481) );
  NAND2_X1 U527 ( .A1(n469), .A2(n481), .ZN(n470) );
  XOR2_X1 U528 ( .A(KEYINPUT95), .B(n470), .Z(n498) );
  NOR2_X1 U529 ( .A1(n486), .A2(n498), .ZN(n479) );
  NAND2_X1 U530 ( .A1(n479), .A2(n513), .ZN(n471) );
  XNOR2_X1 U531 ( .A(n472), .B(n471), .ZN(n473) );
  XOR2_X1 U532 ( .A(G1GAT), .B(n473), .Z(G1324GAT) );
  XOR2_X1 U533 ( .A(G8GAT), .B(KEYINPUT97), .Z(n475) );
  NAND2_X1 U534 ( .A1(n479), .A2(n515), .ZN(n474) );
  XNOR2_X1 U535 ( .A(n475), .B(n474), .ZN(G1325GAT) );
  XOR2_X1 U536 ( .A(KEYINPUT98), .B(KEYINPUT35), .Z(n477) );
  NAND2_X1 U537 ( .A1(n479), .A2(n525), .ZN(n476) );
  XNOR2_X1 U538 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U539 ( .A(G15GAT), .B(n478), .ZN(G1326GAT) );
  NAND2_X1 U540 ( .A1(n518), .A2(n479), .ZN(n480) );
  XNOR2_X1 U541 ( .A(n480), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U542 ( .A(G29GAT), .B(KEYINPUT39), .Z(n490) );
  NAND2_X1 U543 ( .A1(n531), .A2(n481), .ZN(n482) );
  NOR2_X1 U544 ( .A1(n482), .A2(n582), .ZN(n485) );
  INV_X1 U545 ( .A(KEYINPUT37), .ZN(n483) );
  OR2_X1 U546 ( .A1(n512), .A2(n486), .ZN(n488) );
  INV_X1 U547 ( .A(KEYINPUT38), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n488), .B(n487), .ZN(n495) );
  NAND2_X1 U549 ( .A1(n513), .A2(n495), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n490), .B(n489), .ZN(G1328GAT) );
  NAND2_X1 U551 ( .A1(n495), .A2(n515), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n491), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U553 ( .A1(n495), .A2(n525), .ZN(n493) );
  XOR2_X1 U554 ( .A(KEYINPUT100), .B(KEYINPUT40), .Z(n492) );
  XNOR2_X1 U555 ( .A(n493), .B(n492), .ZN(n494) );
  XOR2_X1 U556 ( .A(G43GAT), .B(n494), .Z(G1330GAT) );
  XOR2_X1 U557 ( .A(G50GAT), .B(KEYINPUT101), .Z(n497) );
  NAND2_X1 U558 ( .A1(n495), .A2(n518), .ZN(n496) );
  XNOR2_X1 U559 ( .A(n497), .B(n496), .ZN(G1331GAT) );
  XNOR2_X1 U560 ( .A(KEYINPUT102), .B(KEYINPUT42), .ZN(n502) );
  XOR2_X1 U561 ( .A(G57GAT), .B(KEYINPUT103), .Z(n500) );
  NAND2_X1 U562 ( .A1(n547), .A2(n571), .ZN(n511) );
  NOR2_X1 U563 ( .A1(n498), .A2(n511), .ZN(n506) );
  NAND2_X1 U564 ( .A1(n506), .A2(n513), .ZN(n499) );
  XNOR2_X1 U565 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U566 ( .A(n502), .B(n501), .ZN(G1332GAT) );
  NAND2_X1 U567 ( .A1(n515), .A2(n506), .ZN(n503) );
  XNOR2_X1 U568 ( .A(n503), .B(KEYINPUT104), .ZN(n504) );
  XNOR2_X1 U569 ( .A(G64GAT), .B(n504), .ZN(G1333GAT) );
  NAND2_X1 U570 ( .A1(n506), .A2(n525), .ZN(n505) );
  XNOR2_X1 U571 ( .A(n505), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U572 ( .A(KEYINPUT106), .B(KEYINPUT43), .Z(n508) );
  NAND2_X1 U573 ( .A1(n506), .A2(n518), .ZN(n507) );
  XNOR2_X1 U574 ( .A(n508), .B(n507), .ZN(n510) );
  XOR2_X1 U575 ( .A(G78GAT), .B(KEYINPUT105), .Z(n509) );
  XNOR2_X1 U576 ( .A(n510), .B(n509), .ZN(G1335GAT) );
  NOR2_X1 U577 ( .A1(n512), .A2(n511), .ZN(n519) );
  NAND2_X1 U578 ( .A1(n513), .A2(n519), .ZN(n514) );
  XNOR2_X1 U579 ( .A(G85GAT), .B(n514), .ZN(G1336GAT) );
  NAND2_X1 U580 ( .A1(n515), .A2(n519), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n516), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U582 ( .A1(n519), .A2(n525), .ZN(n517) );
  XNOR2_X1 U583 ( .A(n517), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U584 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n523) );
  XOR2_X1 U585 ( .A(KEYINPUT108), .B(KEYINPUT107), .Z(n521) );
  NAND2_X1 U586 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U587 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U588 ( .A(n523), .B(n522), .ZN(G1339GAT) );
  NAND2_X1 U589 ( .A1(n525), .A2(n524), .ZN(n526) );
  NOR2_X1 U590 ( .A1(n541), .A2(n526), .ZN(n536) );
  NAND2_X1 U591 ( .A1(n536), .A2(n544), .ZN(n527) );
  XNOR2_X1 U592 ( .A(n527), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT111), .B(KEYINPUT49), .Z(n529) );
  NAND2_X1 U594 ( .A1(n536), .A2(n547), .ZN(n528) );
  XNOR2_X1 U595 ( .A(n529), .B(n528), .ZN(n530) );
  XOR2_X1 U596 ( .A(G120GAT), .B(n530), .Z(G1341GAT) );
  XNOR2_X1 U597 ( .A(G127GAT), .B(KEYINPUT112), .ZN(n535) );
  XOR2_X1 U598 ( .A(KEYINPUT50), .B(KEYINPUT113), .Z(n533) );
  INV_X1 U599 ( .A(n531), .ZN(n579) );
  NAND2_X1 U600 ( .A1(n536), .A2(n579), .ZN(n532) );
  XNOR2_X1 U601 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n535), .B(n534), .ZN(G1342GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT114), .B(KEYINPUT51), .Z(n538) );
  NAND2_X1 U604 ( .A1(n536), .A2(n561), .ZN(n537) );
  XNOR2_X1 U605 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U606 ( .A(G134GAT), .B(n539), .ZN(G1343GAT) );
  NOR2_X1 U607 ( .A1(n541), .A2(n540), .ZN(n542) );
  NAND2_X1 U608 ( .A1(n569), .A2(n542), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n543), .B(KEYINPUT115), .ZN(n554) );
  NAND2_X1 U610 ( .A1(n554), .A2(n544), .ZN(n545) );
  XNOR2_X1 U611 ( .A(n545), .B(KEYINPUT116), .ZN(n546) );
  XNOR2_X1 U612 ( .A(G141GAT), .B(n546), .ZN(G1344GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT53), .B(KEYINPUT117), .Z(n549) );
  NAND2_X1 U614 ( .A1(n554), .A2(n547), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n549), .B(n548), .ZN(n551) );
  XOR2_X1 U616 ( .A(G148GAT), .B(KEYINPUT52), .Z(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(G1345GAT) );
  NAND2_X1 U618 ( .A1(n579), .A2(n554), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n552), .B(KEYINPUT118), .ZN(n553) );
  XNOR2_X1 U620 ( .A(G155GAT), .B(n553), .ZN(G1346GAT) );
  XOR2_X1 U621 ( .A(G162GAT), .B(KEYINPUT119), .Z(n556) );
  NAND2_X1 U622 ( .A1(n554), .A2(n561), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(G1347GAT) );
  XOR2_X1 U624 ( .A(G183GAT), .B(KEYINPUT123), .Z(n558) );
  NAND2_X1 U625 ( .A1(n562), .A2(n579), .ZN(n557) );
  XNOR2_X1 U626 ( .A(n558), .B(n557), .ZN(G1350GAT) );
  XNOR2_X1 U627 ( .A(G190GAT), .B(KEYINPUT125), .ZN(n559) );
  XNOR2_X1 U628 ( .A(n559), .B(KEYINPUT124), .ZN(n560) );
  XOR2_X1 U629 ( .A(KEYINPUT58), .B(n560), .Z(n564) );
  NAND2_X1 U630 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(G1351GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT60), .B(KEYINPUT126), .Z(n566) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n565) );
  XNOR2_X1 U634 ( .A(n566), .B(n565), .ZN(n573) );
  AND2_X1 U635 ( .A1(n568), .A2(n567), .ZN(n570) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n581) );
  NOR2_X1 U637 ( .A1(n571), .A2(n581), .ZN(n572) );
  XOR2_X1 U638 ( .A(n573), .B(n572), .Z(G1352GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT61), .B(KEYINPUT127), .Z(n576) );
  INV_X1 U640 ( .A(n581), .ZN(n578) );
  NAND2_X1 U641 ( .A1(n578), .A2(n574), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n577) );
  XOR2_X1 U643 ( .A(G204GAT), .B(n577), .Z(G1353GAT) );
  NAND2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n580), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U647 ( .A(KEYINPUT62), .B(n583), .Z(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

