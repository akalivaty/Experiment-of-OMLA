//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 1 1 1 0 0 1 1 0 1 0 1 1 1 0 0 0 0 0 1 0 0 1 0 0 1 0 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n738, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n861, new_n862, new_n863,
    new_n864, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT84), .ZN(new_n203));
  XNOR2_X1  g002(.A(G197gat), .B(G204gat), .ZN(new_n204));
  INV_X1    g003(.A(G211gat), .ZN(new_n205));
  INV_X1    g004(.A(G218gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n204), .B1(KEYINPUT22), .B2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G211gat), .B(G218gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT77), .ZN(new_n212));
  AND2_X1   g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G155gat), .ZN(new_n217));
  OR2_X1    g016(.A1(KEYINPUT76), .A2(G162gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(KEYINPUT76), .A2(G162gat), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT2), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n216), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  AND2_X1   g021(.A1(G141gat), .A2(G148gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(G141gat), .A2(G148gat), .ZN(new_n224));
  OAI21_X1  g023(.A(KEYINPUT75), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G141gat), .ZN(new_n226));
  INV_X1    g025(.A(G148gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT75), .ZN(new_n229));
  NAND2_X1  g028(.A1(G141gat), .A2(G148gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  AND2_X1   g030(.A1(new_n225), .A2(new_n231), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n212), .B1(new_n222), .B2(new_n232), .ZN(new_n233));
  AND2_X1   g032(.A1(KEYINPUT76), .A2(G162gat), .ZN(new_n234));
  NOR2_X1   g033(.A1(KEYINPUT76), .A2(G162gat), .ZN(new_n235));
  OAI21_X1  g034(.A(G155gat), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n215), .B1(new_n236), .B2(KEYINPUT2), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n225), .A2(new_n231), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n237), .A2(KEYINPUT77), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n233), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT74), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n216), .A2(new_n242), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n228), .B(new_n230), .C1(new_n213), .C2(new_n221), .ZN(new_n244));
  OR2_X1    g043(.A1(new_n213), .A2(new_n242), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n243), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n240), .A2(new_n241), .A3(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT29), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n211), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n241), .B1(new_n210), .B2(KEYINPUT29), .ZN(new_n250));
  AND3_X1   g049(.A1(new_n237), .A2(KEYINPUT77), .A3(new_n238), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT77), .B1(new_n237), .B2(new_n238), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n246), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n250), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n203), .B1(new_n249), .B2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(G22gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n254), .A2(KEYINPUT85), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT85), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n250), .A2(new_n259), .A3(new_n253), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n258), .A2(G228gat), .A3(G233gat), .A4(new_n260), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n256), .B(new_n257), .C1(new_n261), .C2(new_n249), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT86), .ZN(new_n263));
  XNOR2_X1  g062(.A(KEYINPUT83), .B(KEYINPUT31), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n264), .B(G50gat), .ZN(new_n265));
  XOR2_X1   g064(.A(G78gat), .B(G106gat), .Z(new_n266));
  XNOR2_X1  g065(.A(new_n265), .B(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n263), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n256), .B1(new_n261), .B2(new_n249), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(G22gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(new_n262), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n263), .A2(new_n270), .A3(new_n262), .A4(new_n267), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n274), .A2(KEYINPUT35), .ZN(new_n275));
  NAND2_X1  g074(.A1(G227gat), .A2(G233gat), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(G169gat), .A2(G176gat), .ZN(new_n278));
  INV_X1    g077(.A(G169gat), .ZN(new_n279));
  INV_X1    g078(.A(G176gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT23), .ZN(new_n282));
  OAI211_X1 g081(.A(KEYINPUT25), .B(new_n278), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n284));
  MUX2_X1   g083(.A(G183gat), .B(new_n284), .S(G190gat), .Z(new_n285));
  OR2_X1    g084(.A1(KEYINPUT66), .A2(KEYINPUT24), .ZN(new_n286));
  NAND2_X1  g085(.A1(G183gat), .A2(G190gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(KEYINPUT66), .A2(KEYINPUT24), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n283), .B1(new_n285), .B2(new_n289), .ZN(new_n290));
  AND2_X1   g089(.A1(KEYINPUT64), .A2(KEYINPUT23), .ZN(new_n291));
  NOR2_X1   g090(.A1(KEYINPUT64), .A2(KEYINPUT23), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n281), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT65), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT65), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n281), .B(new_n295), .C1(new_n291), .C2(new_n292), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n290), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n278), .B1(new_n281), .B2(new_n282), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT24), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n287), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n299), .B1(new_n285), .B2(new_n301), .ZN(new_n302));
  AND2_X1   g101(.A1(new_n297), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n298), .B1(new_n303), .B2(KEYINPUT25), .ZN(new_n304));
  XOR2_X1   g103(.A(G127gat), .B(G134gat), .Z(new_n305));
  INV_X1    g104(.A(KEYINPUT1), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n306), .B1(G113gat), .B2(G120gat), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  XOR2_X1   g107(.A(KEYINPUT68), .B(G120gat), .Z(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(G113gat), .ZN(new_n310));
  INV_X1    g109(.A(G113gat), .ZN(new_n311));
  INV_X1    g110(.A(G120gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  OR2_X1    g112(.A1(new_n313), .A2(new_n307), .ZN(new_n314));
  AOI22_X1  g113(.A1(new_n308), .A2(new_n310), .B1(new_n314), .B2(new_n305), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT26), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n287), .B1(new_n281), .B2(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(KEYINPUT26), .B1(new_n279), .B2(new_n280), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n318), .B1(new_n278), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(G183gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT27), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT27), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(G183gat), .ZN(new_n324));
  AND3_X1   g123(.A1(new_n322), .A2(new_n324), .A3(KEYINPUT67), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT67), .B1(new_n322), .B2(new_n324), .ZN(new_n326));
  INV_X1    g125(.A(G190gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(KEYINPUT28), .ZN(new_n328));
  NOR3_X1   g127(.A1(new_n325), .A2(new_n326), .A3(new_n328), .ZN(new_n329));
  AND2_X1   g128(.A1(new_n322), .A2(new_n324), .ZN(new_n330));
  AOI21_X1  g129(.A(KEYINPUT28), .B1(new_n330), .B2(new_n327), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n320), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n304), .A2(new_n316), .A3(new_n332), .ZN(new_n333));
  AND2_X1   g132(.A1(new_n290), .A2(new_n297), .ZN(new_n334));
  AOI21_X1  g133(.A(KEYINPUT25), .B1(new_n297), .B2(new_n302), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n332), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(new_n315), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n277), .B1(new_n333), .B2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT69), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(KEYINPUT34), .ZN(new_n340));
  AND2_X1   g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n338), .A2(new_n342), .ZN(new_n343));
  OR2_X1    g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(G15gat), .B(G43gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(G71gat), .B(G99gat), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n345), .B(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n333), .A2(new_n337), .A3(new_n277), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT33), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n348), .A2(KEYINPUT32), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n348), .B(KEYINPUT32), .C1(new_n349), .C2(new_n347), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  OR3_X1    g153(.A1(new_n344), .A2(new_n354), .A3(KEYINPUT70), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n344), .A2(new_n354), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n341), .A2(new_n343), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n357), .A2(new_n352), .A3(new_n353), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n356), .A2(new_n358), .A3(KEYINPUT70), .ZN(new_n359));
  AND3_X1   g158(.A1(new_n355), .A2(new_n359), .A3(KEYINPUT89), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT89), .B1(new_n355), .B2(new_n359), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n275), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n363), .A2(new_n247), .A3(new_n316), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n246), .B(new_n315), .C1(new_n251), .C2(new_n252), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT4), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT4), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n240), .A2(new_n367), .A3(new_n246), .A4(new_n315), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(G225gat), .A2(G233gat), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n364), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n253), .A2(new_n316), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT78), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n372), .A2(new_n373), .A3(new_n365), .ZN(new_n374));
  INV_X1    g173(.A(new_n370), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n253), .A2(KEYINPUT78), .A3(new_n316), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n371), .A2(new_n377), .A3(KEYINPUT5), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(KEYINPUT79), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT79), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n371), .A2(new_n377), .A3(new_n380), .A4(KEYINPUT5), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT81), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n366), .A2(new_n383), .A3(new_n368), .ZN(new_n384));
  INV_X1    g183(.A(new_n253), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n385), .A2(KEYINPUT81), .A3(new_n367), .A4(new_n315), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n384), .A2(new_n364), .A3(new_n386), .ZN(new_n387));
  NOR3_X1   g186(.A1(new_n387), .A2(KEYINPUT5), .A3(new_n375), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n382), .A2(new_n389), .ZN(new_n390));
  XOR2_X1   g189(.A(G1gat), .B(G29gat), .Z(new_n391));
  XNOR2_X1  g190(.A(G57gat), .B(G85gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n391), .B(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n394));
  XOR2_X1   g193(.A(new_n393), .B(new_n394), .Z(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n390), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n388), .B1(new_n379), .B2(new_n381), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT6), .B1(new_n398), .B2(new_n395), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n390), .A2(KEYINPUT6), .A3(new_n396), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  XOR2_X1   g201(.A(G8gat), .B(G36gat), .Z(new_n403));
  XNOR2_X1  g202(.A(new_n403), .B(KEYINPUT72), .ZN(new_n404));
  XNOR2_X1  g203(.A(G64gat), .B(G92gat), .ZN(new_n405));
  XOR2_X1   g204(.A(new_n404), .B(new_n405), .Z(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT71), .ZN(new_n408));
  NAND2_X1  g207(.A1(G226gat), .A2(G233gat), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n410), .B1(new_n336), .B2(new_n248), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n409), .B1(new_n304), .B2(new_n332), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n408), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT29), .B1(new_n304), .B2(new_n332), .ZN(new_n414));
  OAI21_X1  g213(.A(KEYINPUT71), .B1(new_n414), .B2(new_n410), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n413), .A2(new_n211), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n336), .A2(new_n410), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n417), .B1(new_n414), .B2(new_n410), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(new_n210), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n407), .B1(new_n416), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT30), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n416), .A2(new_n419), .A3(new_n407), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n420), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n416), .A2(KEYINPUT30), .A3(new_n419), .A4(new_n407), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT73), .ZN(new_n425));
  AND2_X1   g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n424), .A2(new_n425), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n423), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n402), .A2(new_n429), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n362), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n274), .ZN(new_n432));
  AND3_X1   g231(.A1(new_n432), .A2(new_n358), .A3(new_n356), .ZN(new_n433));
  AOI21_X1  g232(.A(KEYINPUT82), .B1(new_n402), .B2(new_n429), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT82), .ZN(new_n435));
  AOI211_X1 g234(.A(new_n435), .B(new_n428), .C1(new_n400), .C2(new_n401), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n433), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n431), .B1(new_n437), .B2(KEYINPUT35), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT37), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n416), .A2(new_n439), .A3(new_n419), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(KEYINPUT88), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT88), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n416), .A2(new_n442), .A3(new_n439), .A4(new_n419), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n416), .A2(new_n419), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n407), .B1(new_n445), .B2(KEYINPUT37), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(KEYINPUT38), .ZN(new_n448));
  INV_X1    g247(.A(new_n422), .ZN(new_n449));
  OR2_X1    g248(.A1(new_n407), .A2(KEYINPUT38), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n413), .A2(new_n210), .A3(new_n415), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n439), .B1(new_n418), .B2(new_n211), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT87), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT87), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n451), .A2(new_n452), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n450), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n449), .B1(new_n457), .B2(new_n444), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n448), .A2(new_n400), .A3(new_n458), .A4(new_n401), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT40), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n387), .A2(new_n375), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT39), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n374), .A2(new_n376), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n462), .B1(new_n463), .B2(new_n370), .ZN(new_n464));
  AND2_X1   g263(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n387), .A2(new_n462), .A3(new_n375), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(new_n395), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n460), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n461), .A2(new_n464), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n469), .A2(KEYINPUT40), .A3(new_n395), .A4(new_n466), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n398), .A2(new_n395), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n274), .B1(new_n473), .B2(new_n428), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n356), .A2(KEYINPUT36), .A3(new_n358), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n355), .A2(new_n359), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n476), .B1(new_n477), .B2(KEYINPUT36), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n434), .A2(new_n436), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n479), .B1(new_n274), .B2(new_n480), .ZN(new_n481));
  OR2_X1    g280(.A1(new_n438), .A2(new_n481), .ZN(new_n482));
  OR2_X1    g281(.A1(G43gat), .A2(G50gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(G43gat), .A2(G50gat), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n483), .A2(KEYINPUT90), .A3(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT90), .ZN(new_n486));
  AND2_X1   g285(.A1(G43gat), .A2(G50gat), .ZN(new_n487));
  NOR2_X1   g286(.A1(G43gat), .A2(G50gat), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n485), .A2(new_n489), .A3(KEYINPUT15), .ZN(new_n490));
  INV_X1    g289(.A(G29gat), .ZN(new_n491));
  INV_X1    g290(.A(G36gat), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n487), .A2(new_n488), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT15), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n491), .A2(new_n492), .A3(KEYINPUT14), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT14), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n498), .B1(G29gat), .B2(G36gat), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n497), .A2(new_n499), .A3(KEYINPUT91), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n497), .A2(new_n499), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT91), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n490), .A2(new_n496), .A3(new_n500), .A4(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(G43gat), .B(G50gat), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n495), .B1(new_n505), .B2(new_n486), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n506), .B(new_n485), .C1(new_n501), .C2(new_n493), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT92), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT17), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n504), .A2(new_n507), .A3(KEYINPUT92), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(G15gat), .B(G22gat), .ZN(new_n514));
  INV_X1    g313(.A(G1gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(KEYINPUT16), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(KEYINPUT94), .ZN(new_n518));
  INV_X1    g317(.A(G8gat), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT94), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n514), .A2(new_n520), .A3(new_n516), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n518), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(KEYINPUT93), .A2(G8gat), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n523), .B1(new_n514), .B2(new_n516), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n524), .B1(G1gat), .B2(new_n514), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n514), .A2(G1gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(new_n523), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n522), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n504), .A2(new_n507), .A3(KEYINPUT17), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n513), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  AND3_X1   g329(.A1(new_n504), .A2(new_n507), .A3(KEYINPUT92), .ZN(new_n531));
  AOI21_X1  g330(.A(KEYINPUT92), .B1(new_n504), .B2(new_n507), .ZN(new_n532));
  NOR3_X1   g331(.A1(new_n531), .A2(new_n532), .A3(new_n528), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(G229gat), .A2(G233gat), .ZN(new_n535));
  XOR2_X1   g334(.A(new_n535), .B(KEYINPUT95), .Z(new_n536));
  NAND3_X1  g335(.A1(new_n530), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT97), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT18), .ZN(new_n539));
  AND3_X1   g338(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n538), .B1(new_n537), .B2(new_n539), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n530), .A2(new_n534), .A3(KEYINPUT18), .A4(new_n536), .ZN(new_n543));
  XOR2_X1   g342(.A(new_n536), .B(KEYINPUT13), .Z(new_n544));
  AND3_X1   g343(.A1(new_n522), .A2(new_n525), .A3(new_n527), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n545), .B1(new_n510), .B2(new_n512), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n544), .B1(new_n533), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT96), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT96), .ZN(new_n549));
  OAI211_X1 g348(.A(new_n549), .B(new_n544), .C1(new_n533), .C2(new_n546), .ZN(new_n550));
  XNOR2_X1  g349(.A(G113gat), .B(G141gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(G197gat), .ZN(new_n552));
  XOR2_X1   g351(.A(KEYINPUT11), .B(G169gat), .Z(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(KEYINPUT12), .ZN(new_n555));
  AND4_X1   g354(.A1(new_n543), .A2(new_n548), .A3(new_n550), .A4(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n537), .A2(new_n539), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n557), .A2(new_n543), .A3(new_n548), .A4(new_n550), .ZN(new_n558));
  INV_X1    g357(.A(new_n555), .ZN(new_n559));
  AOI22_X1  g358(.A1(new_n542), .A2(new_n556), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(G71gat), .ZN(new_n562));
  INV_X1    g361(.A(G78gat), .ZN(new_n563));
  OAI21_X1  g362(.A(KEYINPUT98), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G57gat), .B(G64gat), .ZN(new_n565));
  AOI21_X1  g364(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G71gat), .B(G78gat), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n566), .ZN(new_n571));
  OR2_X1    g370(.A1(G57gat), .A2(G64gat), .ZN(new_n572));
  NAND2_X1  g371(.A1(G57gat), .A2(G64gat), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n574), .A2(new_n568), .A3(new_n564), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n570), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(KEYINPUT21), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n528), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(KEYINPUT101), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n576), .A2(KEYINPUT21), .ZN(new_n580));
  XNOR2_X1  g379(.A(KEYINPUT100), .B(KEYINPUT19), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n579), .B(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(G127gat), .B(G155gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(KEYINPUT20), .ZN(new_n585));
  NAND2_X1  g384(.A1(G231gat), .A2(G233gat), .ZN(new_n586));
  XOR2_X1   g385(.A(new_n586), .B(KEYINPUT99), .Z(new_n587));
  XNOR2_X1  g386(.A(new_n585), .B(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G183gat), .B(G211gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n583), .B(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G134gat), .B(G162gat), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n531), .A2(new_n532), .ZN(new_n593));
  NAND3_X1  g392(.A1(KEYINPUT103), .A2(G85gat), .A3(G92gat), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(KEYINPUT7), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT7), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n596), .A2(KEYINPUT103), .A3(G85gat), .A4(G92gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G99gat), .B(G106gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(G99gat), .A2(G106gat), .ZN(new_n600));
  INV_X1    g399(.A(G85gat), .ZN(new_n601));
  INV_X1    g400(.A(G92gat), .ZN(new_n602));
  AOI22_X1  g401(.A1(KEYINPUT8), .A2(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  AND3_X1   g402(.A1(new_n598), .A2(new_n599), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n599), .B1(new_n598), .B2(new_n603), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AND2_X1   g405(.A1(G232gat), .A2(G233gat), .ZN(new_n607));
  AOI22_X1  g406(.A1(new_n593), .A2(new_n606), .B1(KEYINPUT41), .B2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n606), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n513), .A2(new_n529), .A3(new_n609), .ZN(new_n610));
  AND2_X1   g409(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g410(.A(G190gat), .B(G218gat), .Z(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT104), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT105), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n592), .B1(new_n611), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n613), .A2(new_n614), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n607), .A2(KEYINPUT41), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(KEYINPUT102), .ZN(new_n619));
  XOR2_X1   g418(.A(new_n617), .B(new_n619), .Z(new_n620));
  AOI21_X1  g419(.A(new_n615), .B1(new_n608), .B2(new_n610), .ZN(new_n621));
  INV_X1    g420(.A(new_n592), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n616), .A2(new_n620), .A3(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n620), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n621), .A2(new_n622), .ZN(new_n626));
  AOI211_X1 g425(.A(new_n615), .B(new_n592), .C1(new_n608), .C2(new_n610), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n625), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n598), .A2(new_n599), .A3(new_n603), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n598), .A2(new_n603), .ZN(new_n631));
  INV_X1    g430(.A(new_n599), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n567), .A2(new_n569), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n568), .B1(new_n574), .B2(new_n564), .ZN(new_n635));
  OAI211_X1 g434(.A(new_n630), .B(new_n633), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  OAI211_X1 g435(.A(new_n570), .B(new_n575), .C1(new_n604), .C2(new_n605), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(G230gat), .A2(G233gat), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(G120gat), .B(G148gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(G176gat), .B(G204gat), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n642), .B(new_n643), .Z(new_n644));
  NAND2_X1  g443(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT10), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n636), .A2(new_n646), .A3(new_n637), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n606), .A2(new_n576), .A3(KEYINPUT10), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT106), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n640), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n647), .A2(KEYINPUT106), .A3(new_n648), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n645), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n639), .B(KEYINPUT107), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n654), .B1(new_n647), .B2(new_n648), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n644), .B1(new_n656), .B2(new_n641), .ZN(new_n657));
  OAI21_X1  g456(.A(KEYINPUT108), .B1(new_n653), .B2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT108), .ZN(new_n659));
  INV_X1    g458(.A(new_n644), .ZN(new_n660));
  INV_X1    g459(.A(new_n641), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n660), .B1(new_n661), .B2(new_n655), .ZN(new_n662));
  AND3_X1   g461(.A1(new_n647), .A2(KEYINPUT106), .A3(new_n648), .ZN(new_n663));
  AOI21_X1  g462(.A(KEYINPUT106), .B1(new_n647), .B2(new_n648), .ZN(new_n664));
  NOR3_X1   g463(.A1(new_n663), .A2(new_n664), .A3(new_n640), .ZN(new_n665));
  OAI211_X1 g464(.A(new_n659), .B(new_n662), .C1(new_n665), .C2(new_n645), .ZN(new_n666));
  AND2_X1   g465(.A1(new_n658), .A2(new_n666), .ZN(new_n667));
  NOR3_X1   g466(.A1(new_n591), .A2(new_n629), .A3(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n482), .A2(new_n561), .A3(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n669), .A2(new_n402), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(new_n515), .ZN(G1324gat));
  XNOR2_X1  g470(.A(KEYINPUT16), .B(G8gat), .ZN(new_n672));
  OR3_X1    g471(.A1(new_n669), .A2(new_n429), .A3(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(G8gat), .B1(new_n669), .B2(new_n429), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  MUX2_X1   g474(.A(new_n673), .B(new_n675), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g475(.A(G15gat), .B1(new_n669), .B2(new_n478), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n360), .A2(new_n361), .ZN(new_n678));
  OR2_X1    g477(.A1(new_n678), .A2(G15gat), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n677), .B1(new_n669), .B2(new_n679), .ZN(G1326gat));
  NOR2_X1   g479(.A1(new_n669), .A2(new_n432), .ZN(new_n681));
  XOR2_X1   g480(.A(KEYINPUT43), .B(G22gat), .Z(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(G1327gat));
  INV_X1    g482(.A(new_n667), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n684), .A2(new_n591), .A3(new_n629), .ZN(new_n685));
  XOR2_X1   g484(.A(new_n685), .B(KEYINPUT109), .Z(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  OAI211_X1 g486(.A(new_n561), .B(new_n687), .C1(new_n438), .C2(new_n481), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n688), .A2(G29gat), .A3(new_n402), .ZN(new_n689));
  XOR2_X1   g488(.A(new_n689), .B(KEYINPUT45), .Z(new_n690));
  OAI21_X1  g489(.A(new_n629), .B1(new_n438), .B2(new_n481), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT44), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  OAI211_X1 g492(.A(KEYINPUT44), .B(new_n629), .C1(new_n438), .C2(new_n481), .ZN(new_n694));
  INV_X1    g493(.A(new_n591), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n695), .A2(new_n560), .A3(new_n667), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n693), .A2(new_n694), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(G29gat), .B1(new_n697), .B2(new_n402), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n690), .A2(new_n698), .ZN(G1328gat));
  NOR3_X1   g498(.A1(new_n688), .A2(G36gat), .A3(new_n429), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT46), .ZN(new_n701));
  OAI21_X1  g500(.A(G36gat), .B1(new_n697), .B2(new_n429), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(G1329gat));
  OR2_X1    g502(.A1(new_n678), .A2(G43gat), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n688), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT110), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n705), .B(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(G43gat), .B1(new_n697), .B2(new_n478), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT47), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n707), .A2(KEYINPUT47), .A3(new_n708), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(G1330gat));
  OAI21_X1  g512(.A(G50gat), .B1(new_n697), .B2(new_n432), .ZN(new_n714));
  OR3_X1    g513(.A1(new_n688), .A2(G50gat), .A3(new_n432), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT48), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n716), .B(new_n717), .ZN(G1331gat));
  NOR3_X1   g517(.A1(new_n561), .A2(new_n591), .A3(new_n629), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n482), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(new_n667), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n721), .A2(new_n402), .ZN(new_n722));
  XOR2_X1   g521(.A(new_n722), .B(G57gat), .Z(G1332gat));
  NOR2_X1   g522(.A1(new_n429), .A2(new_n684), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n720), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n725), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n726));
  XOR2_X1   g525(.A(KEYINPUT49), .B(G64gat), .Z(new_n727));
  OAI21_X1  g526(.A(new_n726), .B1(new_n725), .B2(new_n727), .ZN(G1333gat));
  OAI21_X1  g527(.A(G71gat), .B1(new_n721), .B2(new_n478), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n678), .A2(G71gat), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n720), .A2(new_n667), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g531(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n729), .A2(new_n731), .A3(new_n733), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(G1334gat));
  NOR2_X1   g536(.A1(new_n721), .A2(new_n432), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(new_n563), .ZN(G1335gat));
  NOR2_X1   g538(.A1(new_n561), .A2(new_n695), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n482), .A2(new_n629), .A3(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT51), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n482), .A2(KEYINPUT51), .A3(new_n629), .A4(new_n740), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n743), .A2(KEYINPUT113), .A3(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT113), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n741), .A2(new_n746), .A3(new_n742), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n402), .A2(G85gat), .A3(new_n684), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n745), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  NOR3_X1   g548(.A1(new_n561), .A2(new_n695), .A3(new_n684), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n693), .A2(new_n694), .A3(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT112), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n402), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n693), .A2(KEYINPUT112), .A3(new_n694), .A4(new_n750), .ZN(new_n755));
  AND3_X1   g554(.A1(new_n753), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n749), .B1(new_n756), .B2(new_n601), .ZN(G1336gat));
  NAND2_X1  g556(.A1(new_n724), .A2(new_n602), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n745), .A2(new_n747), .A3(new_n759), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n693), .A2(new_n428), .A3(new_n694), .A4(new_n750), .ZN(new_n761));
  AOI21_X1  g560(.A(KEYINPUT52), .B1(new_n761), .B2(G92gat), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n758), .B(KEYINPUT114), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n764), .B1(new_n743), .B2(new_n744), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n753), .A2(new_n428), .A3(new_n755), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n765), .B1(new_n766), .B2(G92gat), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT52), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n763), .B1(new_n767), .B2(new_n768), .ZN(G1337gat));
  INV_X1    g568(.A(new_n478), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n753), .A2(new_n770), .A3(new_n755), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(G99gat), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n678), .A2(G99gat), .A3(new_n684), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n745), .A2(new_n747), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n774), .ZN(G1338gat));
  NOR3_X1   g574(.A1(new_n432), .A2(G106gat), .A3(new_n684), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n745), .A2(new_n747), .A3(new_n776), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n693), .A2(new_n274), .A3(new_n694), .A4(new_n750), .ZN(new_n778));
  AOI21_X1  g577(.A(KEYINPUT53), .B1(new_n778), .B2(G106gat), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(new_n776), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n781), .B1(new_n743), .B2(new_n744), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n753), .A2(new_n274), .A3(new_n755), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n782), .B1(new_n783), .B2(G106gat), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT53), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n780), .B1(new_n784), .B2(new_n785), .ZN(G1339gat));
  NOR2_X1   g585(.A1(new_n560), .A2(G113gat), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n719), .A2(new_n684), .ZN(new_n788));
  INV_X1    g587(.A(new_n541), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n556), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n536), .B1(new_n530), .B2(new_n534), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n533), .A2(new_n546), .A3(new_n544), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n554), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n791), .A2(new_n667), .A3(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n660), .B1(new_n656), .B2(KEYINPUT54), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT55), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n647), .A2(new_n648), .A3(new_n654), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(KEYINPUT54), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n665), .A2(KEYINPUT115), .A3(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT115), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n651), .A2(new_n652), .ZN(new_n803));
  INV_X1    g602(.A(new_n800), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n802), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n798), .B1(new_n801), .B2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(new_n653), .ZN(new_n807));
  OAI21_X1  g606(.A(KEYINPUT115), .B1(new_n665), .B2(new_n800), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n803), .A2(new_n802), .A3(new_n804), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n796), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  OAI211_X1 g609(.A(new_n806), .B(new_n807), .C1(new_n810), .C2(KEYINPUT55), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n795), .B1(new_n811), .B2(new_n560), .ZN(new_n812));
  INV_X1    g611(.A(new_n629), .ZN(new_n813));
  AND3_X1   g612(.A1(new_n629), .A2(new_n791), .A3(new_n794), .ZN(new_n814));
  INV_X1    g613(.A(new_n811), .ZN(new_n815));
  AOI22_X1  g614(.A1(new_n812), .A2(new_n813), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n591), .B1(new_n816), .B2(KEYINPUT116), .ZN(new_n817));
  INV_X1    g616(.A(new_n796), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n818), .B1(new_n801), .B2(new_n805), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n797), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n808), .A2(new_n809), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n653), .B1(new_n821), .B2(new_n798), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n558), .A2(new_n559), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n548), .A2(new_n543), .A3(new_n550), .A4(new_n555), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n824), .A2(new_n540), .A3(new_n541), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n820), .B(new_n822), .C1(new_n823), .C2(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n629), .B1(new_n826), .B2(new_n795), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT116), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n629), .A2(new_n791), .A3(new_n794), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n829), .A2(new_n811), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n827), .A2(new_n828), .A3(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n788), .B1(new_n817), .B2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT117), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n828), .B1(new_n827), .B2(new_n830), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n812), .A2(new_n813), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n814), .A2(new_n815), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n836), .A2(KEYINPUT116), .A3(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n835), .A2(new_n838), .A3(new_n591), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n839), .A2(KEYINPUT117), .A3(new_n788), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n834), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n841), .A2(new_n402), .ZN(new_n842));
  AND3_X1   g641(.A1(new_n842), .A2(KEYINPUT120), .A3(new_n433), .ZN(new_n843));
  AOI21_X1  g642(.A(KEYINPUT120), .B1(new_n842), .B2(new_n433), .ZN(new_n844));
  OAI211_X1 g643(.A(new_n429), .B(new_n787), .C1(new_n843), .C2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n754), .A2(new_n429), .ZN(new_n846));
  OR2_X1    g645(.A1(new_n846), .A2(new_n678), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n834), .A2(new_n432), .A3(new_n840), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT118), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n834), .A2(KEYINPUT118), .A3(new_n432), .A4(new_n840), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n847), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n311), .B1(new_n852), .B2(new_n561), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n853), .A2(KEYINPUT119), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n853), .A2(KEYINPUT119), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n845), .B1(new_n854), .B2(new_n855), .ZN(G1340gat));
  NOR2_X1   g655(.A1(new_n684), .A2(new_n309), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n429), .B(new_n857), .C1(new_n843), .C2(new_n844), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n852), .A2(new_n667), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n858), .B1(new_n859), .B2(new_n312), .ZN(G1341gat));
  NOR2_X1   g659(.A1(new_n591), .A2(G127gat), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n429), .B(new_n861), .C1(new_n843), .C2(new_n844), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n852), .A2(new_n695), .ZN(new_n863));
  INV_X1    g662(.A(G127gat), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n862), .B1(new_n863), .B2(new_n864), .ZN(G1342gat));
  NOR3_X1   g664(.A1(new_n428), .A2(G134gat), .A3(new_n813), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n866), .B1(new_n843), .B2(new_n844), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(KEYINPUT56), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT56), .ZN(new_n869));
  OAI211_X1 g668(.A(new_n869), .B(new_n866), .C1(new_n843), .C2(new_n844), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n852), .A2(new_n629), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(G134gat), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n868), .A2(new_n870), .A3(new_n872), .ZN(G1343gat));
  INV_X1    g672(.A(KEYINPUT58), .ZN(new_n874));
  AND3_X1   g673(.A1(new_n839), .A2(KEYINPUT117), .A3(new_n788), .ZN(new_n875));
  AOI21_X1  g674(.A(KEYINPUT117), .B1(new_n839), .B2(new_n788), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT57), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n877), .A2(new_n878), .A3(new_n274), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n816), .A2(KEYINPUT121), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n591), .B1(new_n836), .B2(KEYINPUT121), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n788), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n878), .B1(new_n882), .B2(new_n274), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n883), .A2(new_n770), .A3(new_n846), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n879), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(G141gat), .B1(new_n885), .B2(new_n560), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n874), .B1(new_n886), .B2(KEYINPUT122), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n770), .A2(new_n432), .ZN(new_n888));
  INV_X1    g687(.A(new_n888), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n889), .A2(new_n428), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n842), .A2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n561), .A2(new_n226), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n886), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n887), .A2(new_n894), .ZN(new_n895));
  OAI221_X1 g694(.A(new_n886), .B1(KEYINPUT122), .B2(new_n874), .C1(new_n892), .C2(new_n893), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(G1344gat));
  NAND3_X1  g696(.A1(new_n891), .A2(new_n227), .A3(new_n667), .ZN(new_n898));
  INV_X1    g697(.A(new_n885), .ZN(new_n899));
  AOI211_X1 g698(.A(KEYINPUT59), .B(new_n227), .C1(new_n899), .C2(new_n667), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT59), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n591), .B1(new_n827), .B2(new_n830), .ZN(new_n902));
  AOI211_X1 g701(.A(KEYINPUT57), .B(new_n432), .C1(new_n902), .C2(new_n788), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n877), .A2(new_n274), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n903), .B1(new_n904), .B2(KEYINPUT57), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n846), .A2(new_n770), .A3(new_n684), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n901), .B1(new_n907), .B2(G148gat), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n898), .B1(new_n900), .B2(new_n908), .ZN(G1345gat));
  NAND3_X1  g708(.A1(new_n891), .A2(new_n217), .A3(new_n695), .ZN(new_n910));
  OAI21_X1  g709(.A(G155gat), .B1(new_n885), .B2(new_n591), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT123), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n912), .B(new_n913), .ZN(G1346gat));
  NAND4_X1  g713(.A1(new_n891), .A2(new_n218), .A3(new_n219), .A4(new_n629), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n899), .A2(KEYINPUT124), .A3(new_n629), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n916), .B1(new_n235), .B2(new_n234), .ZN(new_n917));
  AOI21_X1  g716(.A(KEYINPUT124), .B1(new_n899), .B2(new_n629), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n915), .B1(new_n917), .B2(new_n918), .ZN(G1347gat));
  NOR2_X1   g718(.A1(new_n841), .A2(new_n754), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n920), .A2(new_n433), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n560), .A2(G169gat), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n921), .A2(new_n428), .A3(new_n922), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n754), .A2(new_n429), .ZN(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n926), .A2(new_n678), .ZN(new_n927));
  INV_X1    g726(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n928), .B1(new_n850), .B2(new_n851), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n279), .B1(new_n929), .B2(new_n561), .ZN(new_n930));
  OAI21_X1  g729(.A(KEYINPUT125), .B1(new_n924), .B2(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT125), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n929), .A2(new_n561), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n923), .B(new_n932), .C1(new_n933), .C2(new_n279), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n931), .A2(new_n934), .ZN(G1348gat));
  NAND3_X1  g734(.A1(new_n921), .A2(new_n280), .A3(new_n724), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n929), .A2(new_n667), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n936), .B1(new_n937), .B2(new_n280), .ZN(G1349gat));
  INV_X1    g737(.A(KEYINPUT126), .ZN(new_n939));
  OR2_X1    g738(.A1(new_n939), .A2(KEYINPUT60), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(KEYINPUT60), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n321), .B1(new_n929), .B2(new_n695), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n591), .A2(new_n326), .A3(new_n325), .ZN(new_n943));
  AND4_X1   g742(.A1(new_n433), .A2(new_n920), .A3(new_n428), .A4(new_n943), .ZN(new_n944));
  OAI211_X1 g743(.A(new_n940), .B(new_n941), .C1(new_n942), .C2(new_n944), .ZN(new_n945));
  AOI21_X1  g744(.A(KEYINPUT118), .B1(new_n877), .B2(new_n432), .ZN(new_n946));
  INV_X1    g745(.A(new_n851), .ZN(new_n947));
  OAI211_X1 g746(.A(new_n695), .B(new_n927), .C1(new_n946), .C2(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(G183gat), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n921), .A2(new_n428), .A3(new_n943), .ZN(new_n950));
  NAND4_X1  g749(.A1(new_n949), .A2(new_n939), .A3(new_n950), .A4(KEYINPUT60), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n945), .A2(new_n951), .ZN(G1350gat));
  NAND4_X1  g751(.A1(new_n921), .A2(new_n327), .A3(new_n428), .A4(new_n629), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT61), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n929), .A2(new_n629), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n954), .B1(new_n955), .B2(G190gat), .ZN(new_n956));
  AOI211_X1 g755(.A(KEYINPUT61), .B(new_n327), .C1(new_n929), .C2(new_n629), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n953), .B1(new_n956), .B2(new_n957), .ZN(G1351gat));
  NOR2_X1   g757(.A1(new_n889), .A2(new_n429), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n920), .A2(new_n959), .ZN(new_n960));
  INV_X1    g759(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g760(.A(G197gat), .B1(new_n961), .B2(new_n561), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n925), .A2(new_n478), .ZN(new_n963));
  AOI211_X1 g762(.A(new_n903), .B(new_n963), .C1(new_n904), .C2(KEYINPUT57), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n561), .A2(G197gat), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n962), .B1(new_n964), .B2(new_n965), .ZN(G1352gat));
  NAND2_X1  g765(.A1(new_n964), .A2(new_n667), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n967), .A2(G204gat), .ZN(new_n968));
  OR2_X1    g767(.A1(new_n684), .A2(G204gat), .ZN(new_n969));
  OAI21_X1  g768(.A(KEYINPUT62), .B1(new_n960), .B2(new_n969), .ZN(new_n970));
  OR3_X1    g769(.A1(new_n960), .A2(KEYINPUT62), .A3(new_n969), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n968), .A2(new_n970), .A3(new_n971), .ZN(G1353gat));
  NAND3_X1  g771(.A1(new_n961), .A2(new_n205), .A3(new_n695), .ZN(new_n973));
  INV_X1    g772(.A(new_n963), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n905), .A2(new_n695), .A3(new_n974), .ZN(new_n975));
  AND3_X1   g774(.A1(new_n975), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n976));
  AOI21_X1  g775(.A(KEYINPUT63), .B1(new_n975), .B2(G211gat), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n973), .B1(new_n976), .B2(new_n977), .ZN(G1354gat));
  INV_X1    g777(.A(KEYINPUT127), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n206), .B1(new_n964), .B2(new_n629), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n629), .A2(new_n206), .ZN(new_n981));
  NOR2_X1   g780(.A1(new_n960), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n979), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n904), .A2(KEYINPUT57), .ZN(new_n984));
  INV_X1    g783(.A(new_n903), .ZN(new_n985));
  NAND4_X1  g784(.A1(new_n984), .A2(new_n629), .A3(new_n985), .A4(new_n974), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n986), .A2(G218gat), .ZN(new_n987));
  OAI211_X1 g786(.A(new_n987), .B(KEYINPUT127), .C1(new_n960), .C2(new_n981), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n983), .A2(new_n988), .ZN(G1355gat));
endmodule


