//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 0 1 0 1 1 1 1 0 0 0 1 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 0 1 0 0 1 1 0 0 1 0 1 0 0 1 0 1 1 1 0 0 0 0 1 0 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:52 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G221), .ZN(new_n189));
  XOR2_X1   g003(.A(KEYINPUT9), .B(G234), .Z(new_n190));
  INV_X1    g004(.A(G902), .ZN(new_n191));
  AOI21_X1  g005(.A(new_n189), .B1(new_n190), .B2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT77), .B(G101), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT3), .ZN(new_n195));
  INV_X1    g009(.A(G107), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n195), .A2(new_n196), .A3(G104), .ZN(new_n197));
  INV_X1    g011(.A(G104), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(G107), .ZN(new_n199));
  AOI21_X1  g013(.A(KEYINPUT3), .B1(new_n198), .B2(G107), .ZN(new_n200));
  OAI211_X1 g014(.A(new_n194), .B(new_n197), .C1(new_n199), .C2(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(G104), .B(G107), .ZN(new_n202));
  INV_X1    g016(.A(G101), .ZN(new_n203));
  OAI21_X1  g017(.A(KEYINPUT78), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT78), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n196), .A2(G104), .ZN(new_n206));
  OAI211_X1 g020(.A(new_n205), .B(G101), .C1(new_n199), .C2(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n201), .A2(new_n204), .A3(new_n207), .ZN(new_n208));
  AND2_X1   g022(.A1(KEYINPUT64), .A2(G146), .ZN(new_n209));
  NOR2_X1   g023(.A1(KEYINPUT64), .A2(G146), .ZN(new_n210));
  OAI21_X1  g024(.A(G143), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT1), .ZN(new_n212));
  INV_X1    g026(.A(G146), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n213), .A2(G143), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n211), .A2(new_n212), .A3(G128), .A4(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G143), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n217), .A2(G146), .ZN(new_n218));
  OAI21_X1  g032(.A(G128), .B1(new_n218), .B2(new_n212), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT64), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(new_n213), .ZN(new_n221));
  NAND2_X1  g035(.A1(KEYINPUT64), .A2(G146), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n217), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n219), .B1(new_n223), .B2(new_n214), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n208), .B1(new_n216), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n216), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n227), .B1(new_n223), .B2(new_n212), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n211), .A2(KEYINPUT68), .A3(KEYINPUT1), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n228), .A2(G128), .A3(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n218), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n221), .A2(new_n222), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n231), .B1(new_n232), .B2(G143), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n226), .B1(new_n230), .B2(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n225), .B1(new_n234), .B2(new_n208), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT11), .ZN(new_n236));
  INV_X1    g050(.A(G134), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n236), .B1(new_n237), .B2(G137), .ZN(new_n238));
  INV_X1    g052(.A(G137), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n239), .A2(KEYINPUT11), .A3(G134), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n237), .A2(G137), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n238), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n242), .B(G131), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  OAI21_X1  g058(.A(KEYINPUT12), .B1(new_n235), .B2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT12), .ZN(new_n246));
  INV_X1    g060(.A(new_n233), .ZN(new_n247));
  INV_X1    g061(.A(G128), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n211), .A2(KEYINPUT1), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n248), .B1(new_n249), .B2(new_n227), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n247), .B1(new_n250), .B2(new_n229), .ZN(new_n251));
  AND3_X1   g065(.A1(new_n201), .A2(new_n204), .A3(new_n207), .ZN(new_n252));
  NOR3_X1   g066(.A1(new_n251), .A2(new_n226), .A3(new_n252), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n246), .B(new_n243), .C1(new_n253), .C2(new_n225), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT10), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n208), .A2(new_n255), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n256), .B1(new_n251), .B2(new_n226), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n214), .B1(new_n232), .B2(G143), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n258), .A2(KEYINPUT65), .A3(KEYINPUT0), .A4(G128), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n211), .A2(KEYINPUT0), .A3(G128), .A4(new_n215), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT65), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n197), .B1(new_n200), .B2(new_n199), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G101), .ZN(new_n265));
  OR2_X1    g079(.A1(new_n265), .A2(KEYINPUT4), .ZN(new_n266));
  XOR2_X1   g080(.A(KEYINPUT0), .B(G128), .Z(new_n267));
  NAND2_X1  g081(.A1(new_n233), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n265), .A2(KEYINPUT4), .A3(new_n201), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n263), .A2(new_n266), .A3(new_n268), .A4(new_n269), .ZN(new_n270));
  AND2_X1   g084(.A1(new_n224), .A2(new_n216), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n255), .B1(new_n271), .B2(new_n208), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n257), .A2(new_n244), .A3(new_n270), .A4(new_n272), .ZN(new_n273));
  XNOR2_X1  g087(.A(G110), .B(G140), .ZN(new_n274));
  INV_X1    g088(.A(G953), .ZN(new_n275));
  AND2_X1   g089(.A1(new_n275), .A2(G227), .ZN(new_n276));
  XOR2_X1   g090(.A(new_n274), .B(new_n276), .Z(new_n277));
  NAND4_X1  g091(.A1(new_n245), .A2(new_n254), .A3(new_n273), .A4(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT80), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n257), .A2(new_n270), .A3(new_n272), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n243), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n273), .ZN(new_n282));
  INV_X1    g096(.A(new_n277), .ZN(new_n283));
  AOI22_X1  g097(.A1(new_n278), .A2(new_n279), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  AND2_X1   g098(.A1(new_n273), .A2(new_n277), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n285), .A2(KEYINPUT80), .A3(new_n254), .A4(new_n245), .ZN(new_n286));
  AOI211_X1 g100(.A(G469), .B(G902), .C1(new_n284), .C2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n285), .A2(KEYINPUT79), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n273), .A2(new_n277), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT79), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n288), .A2(new_n281), .A3(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n245), .A2(new_n254), .A3(new_n273), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n283), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n292), .A2(G469), .A3(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G469), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n296), .A2(new_n191), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n193), .B1(new_n287), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(G210), .B1(G237), .B2(G902), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(G116), .B(G119), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  XNOR2_X1  g118(.A(KEYINPUT2), .B(G113), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  XOR2_X1   g120(.A(KEYINPUT81), .B(KEYINPUT5), .Z(new_n307));
  OR2_X1    g121(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G113), .ZN(new_n309));
  INV_X1    g123(.A(G116), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n310), .A2(G119), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n309), .B1(new_n307), .B2(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n306), .B1(new_n308), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(new_n252), .ZN(new_n314));
  XOR2_X1   g128(.A(new_n303), .B(new_n305), .Z(new_n315));
  NAND3_X1  g129(.A1(new_n266), .A2(new_n315), .A3(new_n269), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(G110), .B(G122), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n317), .A2(new_n319), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n321), .A2(KEYINPUT6), .A3(new_n322), .ZN(new_n323));
  OR2_X1    g137(.A1(new_n323), .A2(KEYINPUT82), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n322), .A2(KEYINPUT6), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n323), .B1(new_n325), .B2(KEYINPUT82), .ZN(new_n326));
  AND2_X1   g140(.A1(new_n260), .A2(new_n261), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n260), .A2(new_n261), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n268), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G125), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n230), .A2(new_n233), .ZN(new_n331));
  INV_X1    g145(.A(G125), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n331), .A2(new_n332), .A3(new_n216), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT83), .B(G224), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n335), .A2(G953), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n334), .B(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n324), .A2(new_n326), .A3(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n318), .B(KEYINPUT8), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n303), .A2(KEYINPUT5), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n306), .B1(new_n312), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n339), .B1(new_n341), .B2(new_n208), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n342), .B1(new_n208), .B2(new_n313), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n333), .A2(KEYINPUT84), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT84), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n234), .A2(new_n345), .A3(new_n332), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n344), .A2(new_n330), .A3(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n336), .ZN(new_n348));
  AND2_X1   g162(.A1(new_n348), .A2(KEYINPUT7), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n343), .B1(new_n347), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n330), .A2(new_n349), .A3(new_n333), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT85), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n330), .A2(KEYINPUT85), .A3(new_n333), .A4(new_n349), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n351), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n320), .B1(new_n357), .B2(KEYINPUT86), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT86), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n351), .A2(new_n356), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(G902), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n338), .B1(new_n361), .B2(KEYINPUT87), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT87), .ZN(new_n363));
  AOI211_X1 g177(.A(new_n363), .B(G902), .C1(new_n358), .C2(new_n360), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n302), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n357), .A2(KEYINPUT86), .ZN(new_n366));
  AND3_X1   g180(.A1(new_n366), .A2(new_n360), .A3(new_n321), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n363), .B1(new_n367), .B2(G902), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n361), .A2(KEYINPUT87), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n368), .A2(new_n301), .A3(new_n369), .A4(new_n338), .ZN(new_n370));
  AOI211_X1 g184(.A(new_n188), .B(new_n300), .C1(new_n365), .C2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n190), .A2(G217), .A3(new_n275), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(G122), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G116), .ZN(new_n375));
  OAI21_X1  g189(.A(KEYINPUT92), .B1(new_n374), .B2(G116), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT92), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n377), .A2(new_n310), .A3(G122), .ZN(new_n378));
  AND2_X1   g192(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT14), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n379), .A2(new_n380), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n375), .B(new_n381), .C1(new_n382), .C2(KEYINPUT93), .ZN(new_n383));
  AND2_X1   g197(.A1(new_n382), .A2(KEYINPUT93), .ZN(new_n384));
  OAI21_X1  g198(.A(G107), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n379), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(new_n375), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n387), .A2(G107), .ZN(new_n388));
  XNOR2_X1  g202(.A(G128), .B(G143), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n389), .B(G134), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n385), .A2(new_n391), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n387), .B(G107), .ZN(new_n393));
  AOI21_X1  g207(.A(KEYINPUT13), .B1(new_n248), .B2(G143), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n394), .A2(new_n237), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n395), .B(new_n389), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n373), .B1(new_n392), .B2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n392), .A2(new_n397), .A3(new_n373), .ZN(new_n400));
  AOI21_X1  g214(.A(G902), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(G478), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n402), .A2(KEYINPUT15), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n401), .A2(KEYINPUT94), .A3(new_n404), .ZN(new_n405));
  AND3_X1   g219(.A1(new_n392), .A2(new_n397), .A3(new_n373), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n191), .B1(new_n406), .B2(new_n398), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT94), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n403), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n407), .A2(new_n408), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n405), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(KEYINPUT95), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT95), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n405), .B(new_n413), .C1(new_n409), .C2(new_n410), .ZN(new_n414));
  AND2_X1   g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  XNOR2_X1  g229(.A(KEYINPUT96), .B(G952), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n416), .A2(G953), .ZN(new_n417));
  NAND2_X1  g231(.A1(G234), .A2(G237), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  XOR2_X1   g233(.A(KEYINPUT21), .B(G898), .Z(new_n420));
  NAND3_X1  g234(.A1(new_n418), .A2(G902), .A3(G953), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n419), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT17), .ZN(new_n424));
  NOR2_X1   g238(.A1(G237), .A2(G953), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(G214), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n426), .A2(new_n217), .ZN(new_n427));
  AOI21_X1  g241(.A(G143), .B1(new_n425), .B2(G214), .ZN(new_n428));
  OAI21_X1  g242(.A(G131), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT88), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI211_X1 g245(.A(KEYINPUT88), .B(G131), .C1(new_n427), .C2(new_n428), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n424), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(G140), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(G125), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT16), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT74), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n332), .A2(G140), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT74), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n440), .B1(new_n436), .B2(new_n442), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n213), .B(new_n438), .C1(new_n443), .C2(new_n437), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n438), .B1(new_n443), .B2(new_n437), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(G146), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n434), .A2(KEYINPUT91), .A3(new_n444), .A4(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT91), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n446), .A2(new_n444), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n448), .B1(new_n449), .B2(new_n433), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n427), .A2(new_n428), .ZN(new_n451));
  INV_X1    g265(.A(G131), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n431), .A2(new_n432), .A3(new_n453), .ZN(new_n454));
  OR2_X1    g268(.A1(new_n454), .A2(KEYINPUT17), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n447), .A2(new_n450), .A3(new_n455), .ZN(new_n456));
  XNOR2_X1  g270(.A(G113), .B(G122), .ZN(new_n457));
  XNOR2_X1  g271(.A(KEYINPUT89), .B(G104), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n457), .B(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n232), .A2(new_n436), .A3(new_n441), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n460), .B1(new_n443), .B2(new_n213), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT18), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n451), .B1(new_n462), .B2(new_n452), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n461), .B(new_n463), .C1(new_n462), .C2(new_n429), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n456), .A2(new_n459), .A3(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n459), .B1(new_n456), .B2(new_n464), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n191), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(G475), .ZN(new_n469));
  INV_X1    g283(.A(new_n232), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT19), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n436), .A2(new_n441), .A3(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n472), .B1(new_n443), .B2(new_n471), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n454), .B(new_n446), .C1(new_n470), .C2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n464), .ZN(new_n475));
  INV_X1    g289(.A(new_n459), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(KEYINPUT90), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT90), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n475), .A2(new_n479), .A3(new_n476), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n465), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT20), .ZN(new_n482));
  NOR2_X1   g296(.A1(G475), .A2(G902), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n482), .B1(new_n481), .B2(new_n483), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n469), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NOR3_X1   g301(.A1(new_n415), .A2(new_n423), .A3(new_n487), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n268), .B(new_n243), .C1(new_n327), .C2(new_n328), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT66), .ZN(new_n490));
  OR2_X1    g304(.A1(new_n242), .A2(G131), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n239), .A2(G134), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n452), .B1(new_n492), .B2(new_n241), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT67), .ZN(new_n494));
  OR2_X1    g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n493), .A2(new_n494), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n491), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n498), .B1(new_n251), .B2(new_n226), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT66), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n263), .A2(new_n500), .A3(new_n268), .A4(new_n243), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n490), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT30), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(KEYINPUT69), .B1(new_n234), .B2(new_n497), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT69), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n498), .B(new_n506), .C1(new_n251), .C2(new_n226), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n505), .A2(new_n507), .A3(KEYINPUT30), .A4(new_n489), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n504), .A2(new_n315), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n315), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n505), .A2(new_n507), .A3(new_n510), .A4(new_n489), .ZN(new_n511));
  XNOR2_X1  g325(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n425), .A2(G210), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n512), .B(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT26), .B(G101), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n514), .B(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n509), .A2(new_n511), .A3(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT31), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(KEYINPUT71), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT28), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n502), .A2(new_n315), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n522), .B1(new_n523), .B2(new_n511), .ZN(new_n524));
  AND2_X1   g338(.A1(new_n489), .A2(new_n510), .ZN(new_n525));
  AOI21_X1  g339(.A(KEYINPUT28), .B1(new_n525), .B2(new_n499), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n516), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  XOR2_X1   g341(.A(KEYINPUT71), .B(KEYINPUT31), .Z(new_n528));
  NAND4_X1  g342(.A1(new_n509), .A2(new_n511), .A3(new_n517), .A4(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n521), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(G472), .A2(G902), .ZN(new_n531));
  AND3_X1   g345(.A1(new_n530), .A2(KEYINPUT32), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(KEYINPUT32), .B1(new_n530), .B2(new_n531), .ZN(new_n533));
  INV_X1    g347(.A(G472), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n509), .A2(new_n511), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n516), .ZN(new_n536));
  INV_X1    g350(.A(new_n234), .ZN(new_n537));
  AOI22_X1  g351(.A1(new_n537), .A2(new_n498), .B1(new_n489), .B2(KEYINPUT66), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n510), .B1(new_n538), .B2(new_n501), .ZN(new_n539));
  INV_X1    g353(.A(new_n511), .ZN(new_n540));
  OAI21_X1  g354(.A(KEYINPUT28), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n526), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n541), .A2(new_n542), .A3(new_n517), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT29), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n536), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n505), .A2(new_n507), .A3(new_n489), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n315), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n511), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n526), .B1(new_n548), .B2(KEYINPUT28), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n516), .A2(new_n544), .ZN(new_n550));
  AOI21_X1  g364(.A(G902), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n534), .B1(new_n545), .B2(new_n551), .ZN(new_n552));
  NOR3_X1   g366(.A1(new_n532), .A2(new_n533), .A3(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(G234), .ZN(new_n554));
  OAI21_X1  g368(.A(G217), .B1(new_n554), .B2(G902), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n555), .B(KEYINPUT72), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT25), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n248), .A2(G119), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n559), .B(KEYINPUT23), .ZN(new_n560));
  INV_X1    g374(.A(G110), .ZN(new_n561));
  OR2_X1    g375(.A1(new_n248), .A2(G119), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT75), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(KEYINPUT24), .B(G110), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(KEYINPUT73), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n562), .A2(new_n559), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n565), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n563), .A2(new_n564), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n460), .B(new_n446), .C1(new_n570), .C2(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n567), .A2(new_n568), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n561), .B1(new_n560), .B2(new_n562), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n449), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(KEYINPUT22), .B(G137), .ZN(new_n578));
  NOR3_X1   g392(.A1(new_n189), .A2(new_n554), .A3(G953), .ZN(new_n579));
  XOR2_X1   g393(.A(new_n578), .B(new_n579), .Z(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n572), .A2(new_n576), .A3(new_n580), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n558), .B1(new_n584), .B2(G902), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n582), .A2(KEYINPUT25), .A3(new_n191), .A4(new_n583), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n557), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n555), .A2(new_n191), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  OAI21_X1  g405(.A(KEYINPUT76), .B1(new_n553), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n530), .A2(new_n531), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT32), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n545), .A2(new_n551), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(G472), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n530), .A2(KEYINPUT32), .A3(new_n531), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n595), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT76), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n599), .A2(new_n600), .A3(new_n590), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n371), .A2(new_n488), .A3(new_n592), .A4(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(KEYINPUT97), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(new_n194), .ZN(G3));
  AOI211_X1 g418(.A(new_n188), .B(new_n423), .C1(new_n365), .C2(new_n370), .ZN(new_n605));
  AOI21_X1  g419(.A(KEYINPUT99), .B1(new_n399), .B2(new_n400), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n606), .A2(KEYINPUT33), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT33), .ZN(new_n608));
  AOI211_X1 g422(.A(KEYINPUT99), .B(new_n608), .C1(new_n399), .C2(new_n400), .ZN(new_n609));
  OR2_X1    g423(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n402), .A2(G902), .ZN(new_n611));
  AOI22_X1  g425(.A1(new_n610), .A2(new_n611), .B1(new_n402), .B2(new_n407), .ZN(new_n612));
  INV_X1    g426(.A(G475), .ZN(new_n613));
  INV_X1    g427(.A(new_n467), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n465), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n613), .B1(new_n615), .B2(new_n191), .ZN(new_n616));
  INV_X1    g430(.A(new_n486), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n616), .B1(new_n617), .B2(new_n484), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n612), .A2(new_n618), .ZN(new_n619));
  OAI211_X1 g433(.A(new_n590), .B(new_n193), .C1(new_n287), .C2(new_n299), .ZN(new_n620));
  NAND2_X1  g434(.A1(KEYINPUT98), .A2(G472), .ZN(new_n621));
  AND3_X1   g435(.A1(new_n530), .A2(new_n191), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n621), .B1(new_n530), .B2(new_n191), .ZN(new_n623));
  NOR3_X1   g437(.A1(new_n620), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n605), .A2(new_n619), .A3(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT34), .B(G104), .Z(new_n626));
  XOR2_X1   g440(.A(new_n626), .B(KEYINPUT100), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n625), .B(new_n627), .ZN(G6));
  AOI21_X1  g442(.A(new_n188), .B1(new_n365), .B2(new_n370), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT101), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n630), .B1(new_n485), .B2(new_n486), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n617), .A2(KEYINPUT101), .A3(new_n484), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n412), .A2(new_n414), .A3(new_n469), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AND3_X1   g449(.A1(new_n629), .A2(new_n422), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n624), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT35), .B(G107), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G9));
  NOR2_X1   g453(.A1(new_n622), .A2(new_n623), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n581), .A2(KEYINPUT36), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n577), .B(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n643), .A2(new_n588), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n587), .A2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n371), .A2(new_n488), .A3(new_n640), .A4(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT37), .B(G110), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G12));
  NOR2_X1   g463(.A1(new_n532), .A2(new_n533), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n645), .B1(new_n650), .B2(new_n597), .ZN(new_n651));
  INV_X1    g465(.A(new_n300), .ZN(new_n652));
  OR2_X1    g466(.A1(new_n421), .A2(G900), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n419), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n631), .A2(new_n632), .A3(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n655), .A2(new_n634), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n629), .A2(new_n651), .A3(new_n652), .A4(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G128), .ZN(G30));
  AND2_X1   g472(.A1(new_n415), .A2(new_n487), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n659), .A2(new_n187), .A3(new_n645), .ZN(new_n660));
  XOR2_X1   g474(.A(new_n654), .B(KEYINPUT39), .Z(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n652), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n660), .B1(KEYINPUT40), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n365), .A2(new_n370), .ZN(new_n665));
  XNOR2_X1  g479(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n516), .B1(new_n509), .B2(new_n511), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n191), .B1(new_n548), .B2(new_n517), .ZN(new_n669));
  OAI21_X1  g483(.A(G472), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n650), .A2(new_n670), .ZN(new_n671));
  OR2_X1    g485(.A1(new_n663), .A2(KEYINPUT40), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n664), .A2(new_n667), .A3(new_n671), .A4(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G143), .ZN(G45));
  OAI21_X1  g488(.A(new_n611), .B1(new_n607), .B2(new_n609), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n675), .B1(G478), .B2(new_n401), .ZN(new_n676));
  AND3_X1   g490(.A1(new_n487), .A2(new_n676), .A3(new_n654), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n629), .A2(new_n651), .A3(new_n652), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G146), .ZN(G48));
  AOI21_X1  g493(.A(new_n591), .B1(new_n650), .B2(new_n597), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n278), .A2(new_n279), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n282), .A2(new_n283), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n681), .A2(new_n286), .A3(new_n682), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n296), .B1(new_n683), .B2(new_n191), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n287), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g499(.A(KEYINPUT103), .B1(new_n685), .B2(new_n193), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT103), .ZN(new_n687));
  NOR4_X1   g501(.A1(new_n287), .A2(new_n684), .A3(new_n687), .A4(new_n192), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n605), .A2(new_n680), .A3(new_n619), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(KEYINPUT41), .B(G113), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G15));
  AND3_X1   g506(.A1(new_n629), .A2(new_n680), .A3(new_n689), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n636), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G116), .ZN(G18));
  AND2_X1   g509(.A1(new_n488), .A2(new_n599), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n696), .A2(new_n629), .A3(new_n646), .A4(new_n689), .ZN(new_n697));
  XOR2_X1   g511(.A(KEYINPUT104), .B(G119), .Z(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G21));
  NAND2_X1  g513(.A1(new_n530), .A2(new_n191), .ZN(new_n700));
  OAI211_X1 g514(.A(new_n521), .B(new_n529), .C1(new_n517), .C2(new_n549), .ZN(new_n701));
  AOI22_X1  g515(.A1(new_n700), .A2(G472), .B1(new_n531), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n590), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n605), .A2(new_n659), .A3(new_n689), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G122), .ZN(G24));
  NAND3_X1  g520(.A1(new_n487), .A2(new_n676), .A3(new_n654), .ZN(new_n707));
  AND2_X1   g521(.A1(new_n701), .A2(new_n531), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n534), .B1(new_n530), .B2(new_n191), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n707), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n629), .A2(new_n646), .A3(new_n710), .A4(new_n689), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G125), .ZN(G27));
  AND3_X1   g526(.A1(new_n365), .A2(new_n187), .A3(new_n370), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n713), .A2(new_n652), .A3(new_n680), .A4(new_n677), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT42), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n365), .A2(new_n370), .A3(new_n652), .A4(new_n187), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n599), .A2(new_n590), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n719), .A2(KEYINPUT42), .A3(new_n677), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G131), .ZN(G33));
  INV_X1    g536(.A(new_n656), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n717), .A2(new_n723), .A3(new_n718), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(new_n237), .ZN(G36));
  AND2_X1   g539(.A1(new_n292), .A2(new_n294), .ZN(new_n726));
  AND2_X1   g540(.A1(new_n726), .A2(KEYINPUT45), .ZN(new_n727));
  OAI21_X1  g541(.A(G469), .B1(new_n726), .B2(KEYINPUT45), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n729), .A2(new_n297), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT105), .ZN(new_n731));
  OR3_X1    g545(.A1(new_n730), .A2(new_n731), .A3(KEYINPUT46), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n731), .B1(new_n730), .B2(KEYINPUT46), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n287), .B1(new_n730), .B2(KEYINPUT46), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n732), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n735), .A2(new_n193), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n662), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n618), .A2(new_n676), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(KEYINPUT43), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n740), .A2(new_n645), .ZN(new_n741));
  INV_X1    g555(.A(new_n640), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT44), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT106), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n743), .A2(new_n744), .ZN(new_n747));
  INV_X1    g561(.A(new_n713), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OAI211_X1 g563(.A(KEYINPUT106), .B(new_n713), .C1(new_n743), .C2(new_n744), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n738), .A2(new_n745), .A3(new_n749), .A4(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(KEYINPUT107), .B(G137), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n751), .B(new_n752), .ZN(G39));
  NOR2_X1   g567(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n754));
  AND2_X1   g568(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n755));
  OAI211_X1 g569(.A(new_n735), .B(new_n193), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n735), .A2(new_n193), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n757), .B1(KEYINPUT108), .B2(KEYINPUT47), .ZN(new_n758));
  NOR4_X1   g572(.A1(new_n748), .A2(new_n599), .A3(new_n590), .A4(new_n707), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n756), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G140), .ZN(G42));
  AND2_X1   g575(.A1(new_n713), .A2(new_n689), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n740), .A2(new_n419), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n762), .A2(new_n763), .A3(new_n680), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(KEYINPUT48), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n765), .A2(KEYINPUT48), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n740), .A2(new_n419), .A3(new_n703), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n768), .A2(new_n629), .A3(new_n689), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(new_n417), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n671), .A2(new_n419), .A3(new_n591), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n762), .A2(new_n771), .ZN(new_n772));
  AOI211_X1 g586(.A(new_n767), .B(new_n770), .C1(new_n619), .C2(new_n772), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n763), .A2(new_n188), .A3(new_n689), .A4(new_n704), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n774), .A2(new_n667), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(KEYINPUT50), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n772), .A2(new_n618), .A3(new_n612), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n762), .A2(new_n763), .A3(new_n646), .A4(new_n702), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n776), .A2(KEYINPUT51), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n768), .A2(new_n713), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n758), .A2(new_n756), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n685), .A2(new_n192), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n766), .B(new_n773), .C1(new_n780), .C2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n783), .B(KEYINPUT114), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT113), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n788), .B1(new_n758), .B2(new_n756), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n758), .A2(new_n788), .A3(new_n756), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n787), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g606(.A(KEYINPUT115), .B1(new_n792), .B2(new_n781), .ZN(new_n793));
  INV_X1    g607(.A(new_n791), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n786), .B1(new_n794), .B2(new_n789), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT115), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n795), .A2(new_n796), .A3(new_n713), .A4(new_n768), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n776), .A2(new_n779), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n793), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT51), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n785), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n654), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n587), .A2(new_n644), .A3(new_n802), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n803), .B(new_n193), .C1(new_n287), .C2(new_n299), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n804), .B1(new_n650), .B2(new_n670), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n629), .A2(new_n805), .A3(new_n659), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n657), .A2(new_n678), .A3(new_n711), .A4(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(KEYINPUT52), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT111), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n371), .B(new_n651), .C1(new_n656), .C2(new_n677), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT52), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n810), .A2(new_n811), .A3(new_n711), .A4(new_n806), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n808), .A2(new_n809), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n809), .B1(new_n808), .B2(new_n812), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT53), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT110), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n665), .A2(new_n488), .A3(new_n187), .A4(new_n652), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n592), .A2(new_n601), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n640), .A2(new_n646), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n818), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g635(.A(KEYINPUT109), .B1(new_n612), .B2(new_n618), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT109), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n487), .A2(new_n676), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n629), .A2(new_n825), .A3(new_n422), .A4(new_n624), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n618), .A2(new_n411), .ZN(new_n827));
  INV_X1    g641(.A(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n629), .A2(new_n422), .A3(new_n624), .A4(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n817), .B1(new_n821), .B2(new_n830), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n605), .B(new_n624), .C1(new_n825), .C2(new_n828), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n832), .A2(new_n602), .A3(new_n647), .A4(KEYINPUT110), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  AND4_X1   g648(.A1(new_n690), .A2(new_n694), .A3(new_n697), .A4(new_n705), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n616), .A2(new_n411), .ZN(new_n836));
  AND4_X1   g650(.A1(new_n632), .A2(new_n631), .A3(new_n836), .A4(new_n654), .ZN(new_n837));
  AOI22_X1  g651(.A1(new_n837), .A2(new_n599), .B1(new_n677), .B2(new_n702), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n838), .A2(new_n717), .A3(new_n645), .ZN(new_n839));
  AOI211_X1 g653(.A(new_n724), .B(new_n839), .C1(new_n716), .C2(new_n720), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n834), .A2(new_n835), .A3(new_n840), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n815), .A2(new_n816), .A3(new_n841), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n834), .A2(new_n835), .A3(new_n840), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n808), .A2(new_n812), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(KEYINPUT53), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(KEYINPUT54), .B1(new_n842), .B2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT112), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n816), .B1(new_n815), .B2(new_n841), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT54), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n843), .A2(KEYINPUT53), .A3(new_n845), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n847), .A2(new_n848), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n844), .A2(KEYINPUT111), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n808), .A2(new_n809), .A3(new_n812), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(KEYINPUT53), .B1(new_n856), .B2(new_n843), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n841), .A2(new_n816), .A3(new_n844), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n857), .A2(KEYINPUT54), .A3(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n856), .A2(new_n843), .A3(KEYINPUT53), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n816), .B1(new_n841), .B2(new_n844), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n850), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(KEYINPUT112), .B1(new_n859), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n801), .A2(new_n853), .A3(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n864), .B1(G952), .B2(G953), .ZN(new_n865));
  NOR4_X1   g679(.A1(new_n739), .A2(new_n188), .A3(new_n192), .A4(new_n591), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT49), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n866), .B1(new_n867), .B2(new_n685), .ZN(new_n868));
  INV_X1    g682(.A(new_n685), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n869), .A2(KEYINPUT49), .ZN(new_n870));
  OR4_X1    g684(.A1(new_n667), .A2(new_n868), .A3(new_n671), .A4(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n865), .A2(new_n871), .ZN(G75));
  NAND2_X1  g686(.A1(new_n324), .A2(new_n326), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n873), .B(new_n337), .ZN(new_n874));
  XOR2_X1   g688(.A(new_n874), .B(KEYINPUT55), .Z(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT56), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n857), .A2(new_n858), .ZN(new_n879));
  OAI21_X1  g693(.A(KEYINPUT116), .B1(new_n879), .B2(new_n191), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n191), .B1(new_n849), .B2(new_n851), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT116), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n878), .B1(new_n884), .B2(new_n302), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n275), .A2(G952), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT56), .B1(new_n881), .B2(G210), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n887), .B1(new_n888), .B2(new_n876), .ZN(new_n889));
  OAI21_X1  g703(.A(KEYINPUT117), .B1(new_n885), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n881), .A2(G210), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(new_n877), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n886), .B1(new_n892), .B2(new_n875), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT117), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n301), .B1(new_n880), .B2(new_n883), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n893), .B(new_n894), .C1(new_n895), .C2(new_n878), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n890), .A2(new_n896), .ZN(G51));
  XNOR2_X1  g711(.A(new_n297), .B(KEYINPUT57), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n850), .B1(new_n849), .B2(new_n851), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n898), .B1(new_n859), .B2(new_n899), .ZN(new_n900));
  OR2_X1    g714(.A1(new_n900), .A2(KEYINPUT118), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(KEYINPUT118), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n683), .B(KEYINPUT119), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n729), .B(KEYINPUT120), .Z(new_n905));
  NAND2_X1  g719(.A1(new_n884), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n886), .B1(new_n904), .B2(new_n906), .ZN(G54));
  INV_X1    g721(.A(KEYINPUT121), .ZN(new_n908));
  INV_X1    g722(.A(new_n481), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n881), .B(KEYINPUT116), .ZN(new_n910));
  NAND2_X1  g724(.A1(KEYINPUT58), .A2(G475), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n908), .B(new_n909), .C1(new_n910), .C2(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n911), .B1(new_n880), .B2(new_n883), .ZN(new_n913));
  OAI21_X1  g727(.A(KEYINPUT121), .B1(new_n913), .B2(new_n481), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n886), .B1(new_n913), .B2(new_n481), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n912), .A2(new_n914), .A3(new_n915), .ZN(G60));
  NAND2_X1  g730(.A1(G478), .A2(G902), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT59), .Z(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n610), .B(new_n919), .C1(new_n859), .C2(new_n899), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n887), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT122), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n918), .B1(new_n863), .B2(new_n853), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n922), .B1(new_n923), .B2(new_n610), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n859), .A2(new_n862), .A3(KEYINPUT112), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n848), .B1(new_n847), .B2(new_n852), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n919), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(new_n610), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n927), .A2(KEYINPUT122), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n921), .B1(new_n924), .B2(new_n929), .ZN(G63));
  NAND2_X1  g744(.A1(G217), .A2(G902), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT60), .Z(new_n932));
  OAI21_X1  g746(.A(new_n932), .B1(new_n857), .B2(new_n858), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n887), .B1(new_n933), .B2(new_n643), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n934), .B1(new_n584), .B2(new_n933), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT61), .ZN(G66));
  INV_X1    g750(.A(new_n335), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n275), .B1(new_n937), .B2(new_n420), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n834), .A2(new_n835), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n938), .B1(new_n939), .B2(new_n275), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n873), .B1(G898), .B2(new_n275), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n940), .B(new_n941), .Z(G69));
  NAND2_X1  g756(.A1(new_n810), .A2(new_n711), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n629), .A2(new_n680), .A3(new_n659), .ZN(new_n944));
  OR4_X1    g758(.A1(KEYINPUT126), .A2(new_n757), .A3(new_n661), .A4(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(KEYINPUT126), .B1(new_n737), .B2(new_n944), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n943), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n947), .A2(new_n751), .A3(new_n760), .ZN(new_n948));
  INV_X1    g762(.A(new_n724), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n721), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(KEYINPUT127), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n751), .A2(new_n760), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT127), .ZN(new_n953));
  INV_X1    g767(.A(new_n950), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n952), .A2(new_n953), .A3(new_n954), .A4(new_n947), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n951), .A2(new_n955), .A3(new_n275), .ZN(new_n956));
  NAND2_X1  g770(.A1(G900), .A2(G953), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n504), .A2(new_n508), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(new_n473), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n956), .A2(new_n957), .A3(new_n959), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n959), .B(KEYINPUT123), .Z(new_n961));
  NAND2_X1  g775(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n673), .A2(new_n711), .A3(new_n810), .A4(new_n962), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n963), .B1(KEYINPUT124), .B2(KEYINPUT62), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n822), .A2(new_n824), .A3(new_n827), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n652), .B(new_n662), .C1(new_n965), .C2(KEYINPUT125), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n966), .B1(KEYINPUT125), .B2(new_n965), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n713), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n952), .B(new_n964), .C1(new_n819), .C2(new_n968), .ZN(new_n969));
  NOR3_X1   g783(.A1(new_n963), .A2(KEYINPUT124), .A3(KEYINPUT62), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n961), .B1(new_n971), .B2(G953), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n960), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n275), .B1(G227), .B2(G900), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n974), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n960), .A2(new_n972), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n975), .A2(new_n977), .ZN(G72));
  NAND2_X1  g792(.A1(G472), .A2(G902), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT63), .Z(new_n980));
  INV_X1    g794(.A(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(new_n939), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n981), .B1(new_n971), .B2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(new_n668), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n887), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n842), .A2(new_n846), .ZN(new_n986));
  AOI211_X1 g800(.A(new_n981), .B(new_n986), .C1(new_n518), .C2(new_n536), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n509), .A2(new_n511), .A3(new_n516), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n951), .A2(new_n955), .A3(new_n982), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n988), .B1(new_n989), .B2(new_n980), .ZN(new_n990));
  NOR3_X1   g804(.A1(new_n985), .A2(new_n987), .A3(new_n990), .ZN(G57));
endmodule


