//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 0 0 0 1 0 0 0 1 0 0 1 0 0 1 0 1 1 0 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 0 1 1 1 0 1 0 1 1 0 1 1 1 0 1 1 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:24 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n743, new_n744, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(G143), .ZN(new_n188));
  OAI21_X1  g002(.A(KEYINPUT1), .B1(new_n188), .B2(G146), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n188), .A2(G146), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G143), .ZN(new_n192));
  OAI211_X1 g006(.A(G128), .B(new_n189), .C1(new_n190), .C2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n188), .A2(G146), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  OAI211_X1 g010(.A(new_n194), .B(new_n195), .C1(KEYINPUT1), .C2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n193), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G125), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(G143), .B(G146), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(KEYINPUT0), .A3(G128), .ZN(new_n203));
  XNOR2_X1  g017(.A(KEYINPUT0), .B(G128), .ZN(new_n204));
  OAI211_X1 g018(.A(new_n203), .B(G125), .C1(new_n202), .C2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G953), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G224), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(KEYINPUT7), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n201), .A2(new_n205), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT92), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT92), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n201), .A2(new_n211), .A3(new_n205), .A4(new_n208), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n201), .A2(new_n205), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT93), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT7), .B1(new_n207), .B2(new_n214), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n215), .B1(new_n214), .B2(new_n207), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  AND3_X1   g031(.A1(new_n210), .A2(new_n212), .A3(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G107), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G104), .ZN(new_n220));
  INV_X1    g034(.A(G104), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G107), .ZN(new_n222));
  AND3_X1   g036(.A1(new_n220), .A2(new_n222), .A3(KEYINPUT83), .ZN(new_n223));
  OAI21_X1  g037(.A(G101), .B1(new_n222), .B2(KEYINPUT83), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT81), .ZN(new_n227));
  OAI22_X1  g041(.A1(new_n227), .A2(KEYINPUT3), .B1(new_n219), .B2(G104), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n229));
  OAI22_X1  g043(.A1(KEYINPUT81), .A2(new_n229), .B1(new_n221), .B2(G107), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n227), .A2(new_n219), .A3(KEYINPUT3), .A4(G104), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n228), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G101), .ZN(new_n233));
  AOI21_X1  g047(.A(KEYINPUT82), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n230), .A2(new_n231), .ZN(new_n235));
  AOI22_X1  g049(.A1(KEYINPUT81), .A2(new_n229), .B1(new_n221), .B2(G107), .ZN(new_n236));
  AND4_X1   g050(.A1(KEYINPUT82), .A2(new_n235), .A3(new_n233), .A4(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n226), .B1(new_n234), .B2(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(G116), .B(G119), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT2), .B(G113), .ZN(new_n241));
  OR2_X1    g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n239), .A2(KEYINPUT5), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(KEYINPUT90), .ZN(new_n244));
  INV_X1    g058(.A(G116), .ZN(new_n245));
  NOR3_X1   g059(.A1(new_n245), .A2(KEYINPUT5), .A3(G119), .ZN(new_n246));
  INV_X1    g060(.A(G113), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n244), .A2(new_n248), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n243), .A2(KEYINPUT90), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n242), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  OR2_X1    g065(.A1(new_n251), .A2(KEYINPUT91), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(KEYINPUT91), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n238), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n241), .ZN(new_n255));
  AOI22_X1  g069(.A1(new_n248), .A2(new_n243), .B1(new_n239), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n238), .A2(new_n256), .ZN(new_n257));
  XNOR2_X1  g071(.A(G110), .B(G122), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n258), .B(KEYINPUT8), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n218), .B1(new_n254), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n235), .A2(new_n236), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n262), .B1(new_n263), .B2(G101), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n264), .B1(new_n234), .B2(new_n237), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n240), .A2(new_n241), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n242), .A2(new_n266), .ZN(new_n267));
  NOR3_X1   g081(.A1(new_n232), .A2(KEYINPUT4), .A3(new_n233), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n265), .A2(new_n267), .A3(new_n269), .ZN(new_n270));
  AND4_X1   g084(.A1(new_n227), .A2(new_n219), .A3(KEYINPUT3), .A4(G104), .ZN(new_n271));
  AOI22_X1  g085(.A1(new_n227), .A2(KEYINPUT3), .B1(new_n219), .B2(G104), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n233), .B(new_n236), .C1(new_n271), .C2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT82), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n235), .A2(KEYINPUT82), .A3(new_n233), .A4(new_n236), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n225), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(new_n256), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n270), .A2(new_n278), .A3(new_n258), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n187), .B1(new_n261), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT89), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n213), .B(new_n207), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n270), .A2(new_n278), .ZN(new_n285));
  INV_X1    g099(.A(new_n258), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(KEYINPUT88), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  AOI22_X1  g102(.A1(new_n279), .A2(KEYINPUT6), .B1(new_n285), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n275), .A2(new_n276), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n268), .B1(new_n290), .B2(new_n264), .ZN(new_n291));
  AOI22_X1  g105(.A1(new_n291), .A2(new_n267), .B1(new_n277), .B2(new_n256), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT6), .ZN(new_n293));
  NOR3_X1   g107(.A1(new_n292), .A2(new_n293), .A3(new_n287), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n283), .B(new_n284), .C1(new_n289), .C2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n285), .A2(KEYINPUT6), .A3(new_n288), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n293), .B1(new_n292), .B2(new_n258), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n292), .A2(new_n287), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n283), .B1(new_n300), .B2(new_n284), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n282), .B1(new_n296), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(G210), .B1(G237), .B2(G902), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n284), .B1(new_n289), .B2(new_n294), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT89), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n295), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n308), .A2(new_n303), .A3(new_n282), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n305), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(G214), .B1(G237), .B2(G902), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G221), .ZN(new_n313));
  XNOR2_X1  g127(.A(KEYINPUT9), .B(G234), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n313), .B1(new_n315), .B2(new_n187), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n316), .B(KEYINPUT80), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT11), .ZN(new_n319));
  INV_X1    g133(.A(G134), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  OR2_X1    g135(.A1(KEYINPUT65), .A2(G137), .ZN(new_n322));
  NAND2_X1  g136(.A1(KEYINPUT65), .A2(G137), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n320), .A2(KEYINPUT64), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT64), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G134), .ZN(new_n327));
  AOI21_X1  g141(.A(G137), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n324), .B1(new_n328), .B2(KEYINPUT11), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  XNOR2_X1  g144(.A(KEYINPUT64), .B(G134), .ZN(new_n331));
  AOI21_X1  g145(.A(G131), .B1(new_n331), .B2(G137), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n325), .A2(new_n327), .A3(G137), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n324), .B(new_n333), .C1(new_n328), .C2(KEYINPUT11), .ZN(new_n334));
  AOI22_X1  g148(.A1(new_n330), .A2(new_n332), .B1(new_n334), .B2(G131), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n203), .B1(new_n202), .B2(new_n204), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n291), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT10), .ZN(new_n339));
  AOI211_X1 g153(.A(KEYINPUT84), .B(new_n339), .C1(new_n277), .C2(new_n199), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n199), .B(new_n226), .C1(new_n234), .C2(new_n237), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT84), .ZN(new_n342));
  AOI21_X1  g156(.A(KEYINPUT10), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n335), .B(new_n338), .C1(new_n340), .C2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n238), .A2(new_n198), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n341), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT12), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n334), .A2(G131), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n332), .B(new_n324), .C1(KEYINPUT11), .C2(new_n328), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n346), .A2(KEYINPUT85), .A3(new_n347), .A4(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n199), .B1(new_n290), .B2(new_n226), .ZN(new_n352));
  AOI211_X1 g166(.A(new_n198), .B(new_n225), .C1(new_n275), .C2(new_n276), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n350), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  OR2_X1    g168(.A1(new_n347), .A2(KEYINPUT85), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n347), .A2(KEYINPUT85), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n344), .A2(new_n351), .A3(new_n357), .ZN(new_n358));
  XNOR2_X1  g172(.A(G110), .B(G140), .ZN(new_n359));
  AND2_X1   g173(.A1(new_n206), .A2(G227), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n359), .B(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT86), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n338), .B1(new_n340), .B2(new_n343), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n350), .ZN(new_n365));
  INV_X1    g179(.A(new_n361), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n365), .A2(new_n344), .A3(new_n366), .ZN(new_n367));
  AND3_X1   g181(.A1(new_n362), .A2(new_n363), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n363), .B1(new_n362), .B2(new_n367), .ZN(new_n369));
  INV_X1    g183(.A(G469), .ZN(new_n370));
  NOR3_X1   g184(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n366), .B1(new_n365), .B2(new_n344), .ZN(new_n372));
  AND4_X1   g186(.A1(new_n344), .A2(new_n357), .A3(new_n351), .A4(new_n366), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n370), .B(new_n187), .C1(new_n372), .C2(new_n373), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n370), .A2(new_n187), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n318), .B1(new_n371), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(KEYINPUT87), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT87), .ZN(new_n380));
  OAI211_X1 g194(.A(new_n380), .B(new_n318), .C1(new_n371), .C2(new_n377), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n312), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  NOR2_X1   g196(.A1(G472), .A2(G902), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT32), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT30), .ZN(new_n387));
  INV_X1    g201(.A(G131), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n333), .A2(new_n388), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n197), .B(new_n193), .C1(new_n329), .C2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n323), .ZN(new_n391));
  NOR2_X1   g205(.A1(KEYINPUT65), .A2(G137), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n320), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT66), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n325), .A2(new_n327), .ZN(new_n395));
  INV_X1    g209(.A(G137), .ZN(new_n396));
  AOI22_X1  g210(.A1(new_n393), .A2(new_n394), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  OAI211_X1 g211(.A(KEYINPUT66), .B(new_n320), .C1(new_n391), .C2(new_n392), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n388), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n390), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n336), .B1(new_n348), .B2(new_n349), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n387), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(KEYINPUT67), .B1(new_n390), .B2(new_n399), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n393), .A2(new_n394), .ZN(new_n404));
  INV_X1    g218(.A(new_n328), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n404), .A2(new_n405), .A3(new_n398), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G131), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT67), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n407), .A2(new_n408), .A3(new_n349), .A4(new_n199), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n403), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(KEYINPUT30), .B1(new_n335), .B2(new_n336), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n402), .B(new_n267), .C1(new_n410), .C2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT68), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n401), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n415), .A2(new_n403), .A3(new_n409), .A4(KEYINPUT30), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n416), .A2(KEYINPUT68), .A3(new_n267), .A4(new_n402), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n267), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n415), .A2(new_n403), .A3(new_n409), .A4(new_n419), .ZN(new_n420));
  OR2_X1    g234(.A1(KEYINPUT69), .A2(G237), .ZN(new_n421));
  NAND2_X1  g235(.A1(KEYINPUT69), .A2(G237), .ZN(new_n422));
  AOI21_X1  g236(.A(G953), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(G210), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n424), .B(KEYINPUT27), .ZN(new_n425));
  XNOR2_X1  g239(.A(KEYINPUT26), .B(G101), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n425), .B(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n420), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n418), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT31), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n418), .A2(KEYINPUT31), .A3(new_n429), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n427), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n267), .B1(new_n400), .B2(new_n401), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n420), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(KEYINPUT28), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n438), .A2(KEYINPUT70), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n400), .A2(new_n401), .ZN(new_n440));
  AOI21_X1  g254(.A(KEYINPUT28), .B1(new_n440), .B2(new_n419), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT28), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n443), .B1(new_n420), .B2(new_n436), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT70), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n442), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n435), .B1(new_n439), .B2(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(KEYINPUT71), .B1(new_n434), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(KEYINPUT31), .B1(new_n418), .B2(new_n429), .ZN(new_n449));
  AOI211_X1 g263(.A(new_n431), .B(new_n428), .C1(new_n414), .C2(new_n417), .ZN(new_n450));
  OAI211_X1 g264(.A(KEYINPUT71), .B(new_n447), .C1(new_n449), .C2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n386), .B1(new_n448), .B2(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n267), .B1(new_n410), .B2(new_n401), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n420), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n441), .B1(new_n455), .B2(KEYINPUT28), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT29), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n435), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(G902), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n418), .A2(new_n420), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT72), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n460), .A2(new_n461), .A3(new_n435), .ZN(new_n462));
  INV_X1    g276(.A(new_n420), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n463), .B1(new_n414), .B2(new_n417), .ZN(new_n464));
  OAI21_X1  g278(.A(KEYINPUT72), .B1(new_n464), .B2(new_n427), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n441), .B1(new_n438), .B2(KEYINPUT70), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n467), .B1(KEYINPUT70), .B2(new_n438), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n457), .B1(new_n468), .B2(new_n435), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n459), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(G472), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n447), .B1(new_n449), .B2(new_n450), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT71), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n384), .B1(new_n474), .B2(new_n451), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n453), .B(new_n471), .C1(KEYINPUT32), .C2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(G234), .ZN(new_n477));
  OAI21_X1  g291(.A(G217), .B1(new_n477), .B2(G902), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n478), .B(KEYINPUT73), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(KEYINPUT24), .B(G110), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT75), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n481), .B(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(G119), .ZN(new_n484));
  OR3_X1    g298(.A1(new_n484), .A2(KEYINPUT74), .A3(G128), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(G128), .ZN(new_n486));
  OAI21_X1  g300(.A(KEYINPUT74), .B1(new_n484), .B2(G128), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT23), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n489), .B1(new_n484), .B2(G128), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n196), .A2(KEYINPUT23), .A3(G119), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(new_n491), .A3(new_n486), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  XOR2_X1   g307(.A(KEYINPUT77), .B(G110), .Z(new_n494));
  AOI22_X1  g308(.A1(new_n483), .A2(new_n488), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(G140), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(G125), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n200), .A2(G140), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n497), .A2(new_n498), .A3(KEYINPUT16), .ZN(new_n499));
  OR3_X1    g313(.A1(new_n200), .A2(KEYINPUT16), .A3(G140), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n499), .A2(new_n500), .A3(G146), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n497), .A2(new_n498), .A3(new_n191), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OR2_X1    g317(.A1(new_n495), .A2(new_n503), .ZN(new_n504));
  OR2_X1    g318(.A1(new_n492), .A2(KEYINPUT76), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n492), .A2(KEYINPUT76), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n505), .A2(new_n506), .A3(G110), .ZN(new_n507));
  AOI21_X1  g321(.A(G146), .B1(new_n499), .B2(new_n500), .ZN(new_n508));
  INV_X1    g322(.A(new_n501), .ZN(new_n509));
  OAI221_X1 g323(.A(new_n507), .B1(new_n508), .B2(new_n509), .C1(new_n483), .C2(new_n488), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n504), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(KEYINPUT78), .ZN(new_n512));
  XNOR2_X1  g326(.A(KEYINPUT22), .B(G137), .ZN(new_n513));
  NOR3_X1   g327(.A1(new_n313), .A2(new_n477), .A3(G953), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n513), .B(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT78), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n504), .A2(new_n510), .A3(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n512), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT79), .ZN(new_n519));
  OR2_X1    g333(.A1(new_n511), .A2(new_n515), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT79), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n512), .A2(new_n521), .A3(new_n515), .A4(new_n517), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n519), .A2(new_n187), .A3(new_n520), .A4(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n480), .B1(new_n523), .B2(KEYINPUT25), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n523), .A2(KEYINPUT25), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n519), .A2(new_n520), .A3(new_n522), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n480), .A2(G902), .ZN(new_n529));
  AOI22_X1  g343(.A1(new_n525), .A2(new_n526), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(G143), .B1(new_n423), .B2(G214), .ZN(new_n531));
  INV_X1    g345(.A(new_n422), .ZN(new_n532));
  NOR2_X1   g346(.A1(KEYINPUT69), .A2(G237), .ZN(new_n533));
  OAI211_X1 g347(.A(G214), .B(new_n206), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n534), .A2(new_n188), .ZN(new_n535));
  OAI211_X1 g349(.A(KEYINPUT18), .B(G131), .C1(new_n531), .C2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n497), .A2(new_n498), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT94), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n497), .A2(new_n498), .A3(KEYINPUT94), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n539), .A2(G146), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(new_n502), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n423), .A2(G143), .A3(G214), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n534), .A2(new_n188), .ZN(new_n544));
  NAND2_X1  g358(.A1(KEYINPUT18), .A2(G131), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n536), .A2(new_n542), .A3(new_n546), .ZN(new_n547));
  AND3_X1   g361(.A1(new_n543), .A2(new_n544), .A3(new_n388), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n388), .B1(new_n543), .B2(new_n544), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n548), .A2(new_n549), .A3(KEYINPUT17), .ZN(new_n550));
  OAI211_X1 g364(.A(KEYINPUT17), .B(G131), .C1(new_n531), .C2(new_n535), .ZN(new_n551));
  OAI21_X1  g365(.A(KEYINPUT97), .B1(new_n509), .B2(new_n508), .ZN(new_n552));
  INV_X1    g366(.A(new_n508), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT97), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n553), .A2(new_n554), .A3(new_n501), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n551), .A2(new_n552), .A3(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n547), .B1(new_n550), .B2(new_n556), .ZN(new_n557));
  XOR2_X1   g371(.A(KEYINPUT95), .B(G104), .Z(new_n558));
  XNOR2_X1  g372(.A(G113), .B(G122), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n558), .B(new_n559), .ZN(new_n560));
  AND2_X1   g374(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n560), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n562), .B(new_n547), .C1(new_n550), .C2(new_n556), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n187), .B1(new_n561), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(G475), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT20), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n539), .A2(KEYINPUT19), .A3(new_n540), .ZN(new_n568));
  OR2_X1    g382(.A1(new_n537), .A2(KEYINPUT19), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n568), .A2(new_n191), .A3(new_n569), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n501), .B(new_n570), .C1(new_n548), .C2(new_n549), .ZN(new_n571));
  AOI211_X1 g385(.A(KEYINPUT96), .B(new_n562), .C1(new_n571), .C2(new_n547), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT96), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n571), .A2(new_n547), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n573), .B1(new_n574), .B2(new_n560), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n572), .B1(new_n575), .B2(new_n563), .ZN(new_n576));
  NOR2_X1   g390(.A1(G475), .A2(G902), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n567), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n574), .A2(new_n560), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n579), .A2(new_n563), .A3(KEYINPUT96), .ZN(new_n580));
  INV_X1    g394(.A(new_n572), .ZN(new_n581));
  AND4_X1   g395(.A1(new_n567), .A2(new_n580), .A3(new_n581), .A4(new_n577), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n566), .B1(new_n578), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n245), .A2(KEYINPUT14), .A3(G122), .ZN(new_n584));
  XOR2_X1   g398(.A(G116), .B(G122), .Z(new_n585));
  OAI211_X1 g399(.A(G107), .B(new_n584), .C1(new_n585), .C2(KEYINPUT14), .ZN(new_n586));
  XNOR2_X1  g400(.A(G116), .B(G122), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(new_n219), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n188), .A2(G128), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n196), .A2(G143), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n331), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n331), .B1(new_n589), .B2(new_n590), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n586), .B(new_n588), .C1(new_n592), .C2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n585), .A2(G107), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n588), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT13), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n589), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n590), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n589), .A2(new_n597), .ZN(new_n600));
  OAI21_X1  g414(.A(G134), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n596), .A2(new_n601), .A3(new_n591), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n594), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n315), .A2(G217), .A3(new_n206), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT98), .ZN(new_n606));
  INV_X1    g420(.A(new_n604), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n594), .A2(new_n602), .A3(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n605), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n603), .A2(KEYINPUT98), .A3(new_n604), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n609), .A2(KEYINPUT99), .A3(new_n187), .A4(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(G478), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n612), .A2(KEYINPUT15), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n611), .B(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(G234), .A2(G237), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n615), .A2(G952), .A3(new_n206), .ZN(new_n616));
  XNOR2_X1  g430(.A(KEYINPUT21), .B(G898), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n615), .A2(G902), .A3(G953), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n616), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(KEYINPUT100), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NOR3_X1   g436(.A1(new_n583), .A2(new_n614), .A3(new_n622), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n382), .A2(new_n476), .A3(new_n530), .A4(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(G101), .ZN(G3));
  INV_X1    g439(.A(new_n530), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n626), .B1(new_n379), .B2(new_n381), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n474), .A2(new_n451), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n187), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n475), .B1(new_n629), .B2(G472), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(new_n631), .B(KEYINPUT101), .Z(new_n632));
  NAND3_X1  g446(.A1(new_n305), .A2(KEYINPUT102), .A3(new_n309), .ZN(new_n633));
  INV_X1    g447(.A(new_n311), .ZN(new_n634));
  AOI211_X1 g448(.A(new_n304), .B(new_n281), .C1(new_n307), .C2(new_n295), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT102), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n634), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n609), .A2(new_n187), .A3(new_n610), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n612), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n609), .A2(new_n610), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT33), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g456(.A(KEYINPUT103), .B1(new_n603), .B2(new_n604), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(new_n608), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n642), .B1(new_n644), .B2(new_n641), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n612), .A2(G902), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n639), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n583), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n650), .A2(new_n622), .ZN(new_n651));
  AND3_X1   g465(.A1(new_n633), .A2(new_n637), .A3(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n632), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT34), .B(G104), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G6));
  OAI211_X1 g470(.A(new_n614), .B(new_n566), .C1(new_n578), .C2(new_n582), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n657), .A2(new_n622), .ZN(new_n658));
  AND3_X1   g472(.A1(new_n633), .A2(new_n637), .A3(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n632), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(KEYINPUT104), .ZN(new_n662));
  XNOR2_X1  g476(.A(KEYINPUT35), .B(G107), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G9));
  NAND2_X1  g478(.A1(new_n379), .A2(new_n381), .ZN(new_n665));
  INV_X1    g479(.A(new_n312), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n512), .A2(new_n517), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n515), .A2(KEYINPUT36), .ZN(new_n668));
  XOR2_X1   g482(.A(new_n667), .B(new_n668), .Z(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n529), .ZN(new_n670));
  INV_X1    g484(.A(new_n526), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n670), .B1(new_n671), .B2(new_n524), .ZN(new_n672));
  AND2_X1   g486(.A1(new_n672), .A2(new_n623), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n630), .A2(new_n665), .A3(new_n666), .A4(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT37), .B(G110), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G12));
  OR2_X1    g490(.A1(new_n619), .A2(G900), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n616), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n657), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n453), .A2(new_n471), .ZN(new_n681));
  AOI21_X1  g495(.A(KEYINPUT32), .B1(new_n628), .B2(new_n383), .ZN(new_n682));
  OAI211_X1 g496(.A(new_n672), .B(new_n680), .C1(new_n681), .C2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n633), .A2(new_n637), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n381), .ZN(new_n686));
  AND2_X1   g500(.A1(new_n374), .A2(new_n376), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n362), .A2(new_n367), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(KEYINPUT86), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n362), .A2(new_n363), .A3(new_n367), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n689), .A2(G469), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n687), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n380), .B1(new_n692), .B2(new_n318), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n685), .B1(new_n686), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g508(.A(KEYINPUT105), .B1(new_n683), .B2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n672), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n628), .A2(new_n383), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n385), .ZN(new_n698));
  AOI22_X1  g512(.A1(new_n628), .A2(new_n386), .B1(new_n470), .B2(G472), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n696), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT105), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n684), .B1(new_n379), .B2(new_n381), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n700), .A2(new_n701), .A3(new_n702), .A4(new_n680), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n695), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G128), .ZN(G30));
  XOR2_X1   g519(.A(new_n310), .B(KEYINPUT38), .Z(new_n706));
  INV_X1    g520(.A(new_n583), .ZN(new_n707));
  INV_X1    g521(.A(new_n614), .ZN(new_n708));
  NOR4_X1   g522(.A1(new_n706), .A2(new_n707), .A3(new_n708), .A4(new_n634), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n678), .B(KEYINPUT39), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n665), .A2(new_n710), .ZN(new_n711));
  OR2_X1    g525(.A1(new_n711), .A2(KEYINPUT40), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(KEYINPUT40), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n464), .A2(new_n435), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n187), .B1(new_n455), .B2(new_n427), .ZN(new_n715));
  OAI21_X1  g529(.A(G472), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  OAI211_X1 g530(.A(new_n453), .B(new_n716), .C1(KEYINPUT32), .C2(new_n475), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n718), .A2(new_n672), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n709), .A2(new_n712), .A3(new_n713), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G143), .ZN(G45));
  NOR2_X1   g535(.A1(new_n650), .A2(new_n679), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n702), .A2(new_n476), .A3(new_n672), .A4(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G146), .ZN(G48));
  OAI21_X1  g538(.A(new_n187), .B1(new_n372), .B2(new_n373), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(G469), .ZN(new_n726));
  INV_X1    g540(.A(new_n316), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n726), .A2(new_n374), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(KEYINPUT106), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT106), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n726), .A2(new_n730), .A3(new_n374), .A4(new_n727), .ZN(new_n731));
  AND2_X1   g545(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n476), .A2(new_n530), .A3(new_n652), .A4(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT107), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n626), .B1(new_n698), .B2(new_n699), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n736), .A2(KEYINPUT107), .A3(new_n652), .A4(new_n732), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(KEYINPUT41), .B(G113), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n738), .B(new_n739), .ZN(G15));
  NAND4_X1  g554(.A1(new_n476), .A2(new_n530), .A3(new_n659), .A4(new_n732), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G116), .ZN(G18));
  AND4_X1   g556(.A1(new_n633), .A2(new_n729), .A3(new_n637), .A4(new_n731), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n476), .A2(new_n743), .A3(new_n623), .A4(new_n672), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G119), .ZN(G21));
  OAI21_X1  g559(.A(new_n434), .B1(new_n427), .B2(new_n456), .ZN(new_n746));
  AOI22_X1  g560(.A1(new_n629), .A2(G472), .B1(new_n383), .B2(new_n746), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n707), .A2(new_n708), .ZN(new_n748));
  AND3_X1   g562(.A1(new_n633), .A2(new_n637), .A3(new_n748), .ZN(new_n749));
  AND3_X1   g563(.A1(new_n729), .A2(new_n621), .A3(new_n731), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n747), .A2(new_n530), .A3(new_n749), .A4(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G122), .ZN(G24));
  NAND2_X1  g566(.A1(new_n746), .A2(new_n383), .ZN(new_n753));
  AOI21_X1  g567(.A(G902), .B1(new_n474), .B2(new_n451), .ZN(new_n754));
  INV_X1    g568(.A(G472), .ZN(new_n755));
  OAI211_X1 g569(.A(new_n672), .B(new_n753), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(new_n722), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n743), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G125), .ZN(G27));
  INV_X1    g574(.A(KEYINPUT109), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n682), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g576(.A(KEYINPUT109), .B1(new_n475), .B2(KEYINPUT32), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n762), .A2(new_n699), .A3(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n305), .A2(new_n311), .A3(new_n309), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n688), .A2(new_n370), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n727), .B1(new_n377), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT42), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n757), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n764), .A2(new_n530), .A3(new_n768), .A4(new_n770), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n476), .A2(new_n530), .A3(new_n722), .A4(new_n768), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT108), .ZN(new_n773));
  AND3_X1   g587(.A1(new_n772), .A2(new_n773), .A3(new_n769), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n773), .B1(new_n772), .B2(new_n769), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n771), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G131), .ZN(G33));
  NAND4_X1  g591(.A1(new_n476), .A2(new_n530), .A3(new_n680), .A4(new_n768), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G134), .ZN(G36));
  AND2_X1   g593(.A1(new_n707), .A2(new_n649), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT110), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n780), .B1(new_n781), .B2(KEYINPUT43), .ZN(new_n782));
  XNOR2_X1  g596(.A(KEYINPUT110), .B(KEYINPUT43), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n782), .B1(new_n780), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n697), .B1(new_n755), .B2(new_n754), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n784), .A2(new_n785), .A3(new_n672), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT44), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n765), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n788), .B1(new_n787), .B2(new_n786), .ZN(new_n789));
  AOI21_X1  g603(.A(KEYINPUT45), .B1(new_n689), .B2(new_n690), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT45), .ZN(new_n791));
  OAI21_X1  g605(.A(G469), .B1(new_n688), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n376), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT46), .ZN(new_n794));
  OR2_X1    g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n374), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n796), .B1(new_n793), .B2(new_n794), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n316), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(new_n710), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n789), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G137), .ZN(G39));
  XOR2_X1   g615(.A(KEYINPUT111), .B(KEYINPUT47), .Z(new_n802));
  OR2_X1    g616(.A1(new_n798), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(KEYINPUT111), .A2(KEYINPUT47), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n798), .A2(new_n804), .ZN(new_n805));
  NOR4_X1   g619(.A1(new_n476), .A2(new_n530), .A3(new_n757), .A4(new_n765), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n803), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  XOR2_X1   g621(.A(KEYINPUT112), .B(G140), .Z(new_n808));
  XNOR2_X1  g622(.A(new_n807), .B(new_n808), .ZN(G42));
  INV_X1    g623(.A(new_n765), .ZN(new_n810));
  AOI21_X1  g624(.A(KEYINPUT116), .B1(new_n732), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n811), .A2(new_n616), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n732), .A2(KEYINPUT116), .A3(new_n810), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n812), .A2(new_n784), .A3(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT117), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n812), .A2(KEYINPUT117), .A3(new_n784), .A4(new_n813), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n756), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n803), .A2(new_n805), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n726), .A2(new_n374), .A3(new_n317), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n747), .A2(new_n530), .ZN(new_n824));
  INV_X1    g638(.A(new_n616), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n784), .A2(new_n825), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n824), .A2(new_n826), .A3(new_n765), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n823), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n812), .A2(new_n813), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n718), .A2(new_n530), .ZN(new_n830));
  NOR4_X1   g644(.A1(new_n829), .A2(new_n830), .A3(new_n583), .A4(new_n649), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n706), .A2(new_n634), .A3(new_n732), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n824), .A2(new_n826), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT50), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n833), .A2(new_n834), .A3(KEYINPUT50), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n820), .A2(new_n828), .A3(new_n832), .A4(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT51), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n756), .B1(new_n816), .B2(new_n817), .ZN(new_n843));
  OAI21_X1  g657(.A(KEYINPUT118), .B1(new_n843), .B2(new_n831), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT119), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n823), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n821), .A2(KEYINPUT119), .A3(new_n822), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n846), .A2(new_n827), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n841), .B1(new_n837), .B2(new_n838), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n844), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n843), .A2(KEYINPUT118), .A3(new_n831), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n842), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n829), .A2(new_n830), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n853), .A2(new_n583), .A3(new_n649), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n206), .A2(G952), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n855), .B1(new_n834), .B2(new_n743), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT48), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n764), .A2(new_n530), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n857), .B1(new_n818), .B2(new_n859), .ZN(new_n860));
  AOI211_X1 g674(.A(KEYINPUT48), .B(new_n858), .C1(new_n816), .C2(new_n817), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n854), .B(new_n856), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  OR2_X1    g676(.A1(new_n862), .A2(KEYINPUT120), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(KEYINPUT120), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n852), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NOR4_X1   g679(.A1(new_n696), .A2(new_n583), .A3(new_n614), .A4(new_n679), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n866), .A2(new_n476), .A3(new_n665), .A4(new_n810), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(new_n778), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n758), .A2(new_n768), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(KEYINPUT114), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT114), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n758), .A2(new_n871), .A3(new_n768), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n868), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n776), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n303), .B1(new_n308), .B2(new_n282), .ZN(new_n875));
  OAI211_X1 g689(.A(new_n311), .B(new_n658), .C1(new_n875), .C2(new_n635), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT113), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n310), .A2(KEYINPUT113), .A3(new_n311), .A4(new_n658), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n310), .A2(new_n651), .A3(new_n311), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n627), .A2(new_n881), .A3(new_n630), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n624), .A2(new_n741), .A3(new_n882), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n744), .A2(new_n674), .A3(new_n751), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n883), .A2(new_n738), .A3(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n874), .A2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT52), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n695), .A2(new_n703), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n767), .A2(new_n679), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n717), .A2(new_n696), .A3(new_n749), .A4(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n759), .A2(new_n723), .A3(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n887), .B1(new_n888), .B2(new_n891), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n759), .A2(new_n723), .A3(new_n890), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n893), .A2(KEYINPUT52), .A3(new_n704), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n886), .A2(KEYINPUT53), .A3(new_n895), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n883), .A2(new_n738), .A3(new_n884), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n897), .A2(new_n776), .A3(new_n873), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n723), .A2(KEYINPUT52), .A3(new_n890), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n899), .A2(new_n704), .A3(new_n759), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT52), .B1(new_n893), .B2(new_n704), .ZN(new_n901));
  OAI21_X1  g715(.A(KEYINPUT115), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT115), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n899), .A2(new_n704), .A3(new_n759), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n892), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n898), .B1(new_n902), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n896), .B1(new_n906), .B2(KEYINPUT53), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n902), .A2(new_n905), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT53), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n874), .A2(new_n909), .A3(new_n885), .ZN(new_n910));
  AOI21_X1  g724(.A(KEYINPUT54), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(new_n894), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n912), .A2(new_n901), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n909), .B1(new_n913), .B2(new_n898), .ZN(new_n914));
  AOI22_X1  g728(.A1(new_n907), .A2(KEYINPUT54), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n865), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n916), .B1(G952), .B2(G953), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n780), .A2(new_n318), .A3(new_n311), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n726), .A2(new_n374), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n919), .A2(KEYINPUT49), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n919), .A2(KEYINPUT49), .ZN(new_n921));
  NOR4_X1   g735(.A1(new_n626), .A2(new_n918), .A3(new_n920), .A4(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n922), .A2(new_n718), .A3(new_n706), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n917), .A2(new_n923), .ZN(G75));
  NOR3_X1   g738(.A1(new_n900), .A2(new_n901), .A3(KEYINPUT115), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n903), .B1(new_n892), .B2(new_n904), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n910), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n914), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n928), .A2(G210), .A3(G902), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT56), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n300), .B(new_n284), .ZN(new_n931));
  XNOR2_X1  g745(.A(KEYINPUT121), .B(KEYINPUT55), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n931), .B(new_n932), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n929), .A2(new_n930), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n933), .B1(new_n929), .B2(new_n930), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n206), .A2(G952), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(G51));
  XNOR2_X1  g751(.A(new_n375), .B(KEYINPUT57), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT122), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT54), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n927), .A2(new_n939), .A3(new_n914), .A4(new_n940), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n897), .A2(KEYINPUT53), .A3(new_n776), .A4(new_n873), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n942), .B1(new_n905), .B2(new_n902), .ZN(new_n943));
  AOI21_X1  g757(.A(KEYINPUT53), .B1(new_n886), .B2(new_n895), .ZN(new_n944));
  OAI21_X1  g758(.A(KEYINPUT54), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n941), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n939), .B1(new_n911), .B2(new_n914), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n938), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  OR2_X1    g762(.A1(new_n372), .A2(new_n373), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n928), .A2(G902), .ZN(new_n951));
  OR3_X1    g765(.A1(new_n951), .A2(new_n790), .A3(new_n792), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n936), .B1(new_n950), .B2(new_n952), .ZN(G54));
  INV_X1    g767(.A(new_n576), .ZN(new_n954));
  NAND2_X1  g768(.A1(KEYINPUT58), .A2(G475), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n954), .B1(new_n951), .B2(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(new_n936), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n951), .A2(new_n954), .A3(new_n955), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n958), .A2(new_n959), .ZN(G60));
  NAND2_X1  g774(.A1(G478), .A2(G902), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT59), .Z(new_n962));
  OAI21_X1  g776(.A(new_n646), .B1(new_n915), .B2(new_n962), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n646), .A2(new_n962), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n964), .B1(new_n946), .B2(new_n947), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n963), .A2(new_n957), .A3(new_n965), .ZN(G63));
  NOR2_X1   g780(.A1(new_n943), .A2(new_n944), .ZN(new_n967));
  NAND2_X1  g781(.A1(G217), .A2(G902), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT123), .Z(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(KEYINPUT60), .Z(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n527), .B1(new_n967), .B2(new_n971), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n928), .A2(new_n669), .A3(new_n970), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n972), .A2(new_n957), .A3(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT61), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n974), .B(new_n975), .ZN(G66));
  INV_X1    g790(.A(G224), .ZN(new_n977));
  OAI21_X1  g791(.A(G953), .B1(new_n617), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n978), .B1(new_n897), .B2(G953), .ZN(new_n979));
  INV_X1    g793(.A(new_n300), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n980), .B1(G898), .B2(new_n206), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n979), .B(new_n981), .ZN(G69));
  AOI21_X1  g796(.A(new_n206), .B1(G227), .B2(G900), .ZN(new_n983));
  INV_X1    g797(.A(new_n807), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n765), .B1(new_n650), .B2(new_n657), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n736), .A2(new_n665), .A3(new_n710), .A4(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n800), .A2(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT124), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n800), .A2(KEYINPUT124), .A3(new_n986), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n984), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  AND3_X1   g805(.A1(new_n704), .A2(new_n723), .A3(new_n759), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(new_n720), .ZN(new_n993));
  OR2_X1    g807(.A1(new_n993), .A2(KEYINPUT62), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(KEYINPUT62), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n991), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n996), .A2(new_n206), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n416), .A2(new_n402), .ZN(new_n998));
  AND2_X1   g812(.A1(new_n568), .A2(new_n569), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n998), .B(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n997), .A2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g815(.A(KEYINPUT125), .B1(new_n206), .B2(G900), .ZN(new_n1002));
  INV_X1    g816(.A(new_n1002), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n859), .A2(new_n710), .A3(new_n749), .A4(new_n798), .ZN(new_n1004));
  AND3_X1   g818(.A1(new_n1004), .A2(new_n778), .A3(new_n807), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(new_n776), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n800), .A2(new_n992), .ZN(new_n1007));
  OR2_X1    g821(.A1(new_n1007), .A2(KEYINPUT126), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1007), .A2(KEYINPUT126), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1006), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n1000), .A2(G953), .ZN(new_n1011));
  INV_X1    g825(.A(new_n1011), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1003), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(new_n1013), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n983), .B1(new_n1001), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g829(.A(new_n1000), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1016), .B1(new_n996), .B2(new_n206), .ZN(new_n1017));
  INV_X1    g831(.A(new_n983), .ZN(new_n1018));
  NOR3_X1   g832(.A1(new_n1017), .A2(new_n1013), .A3(new_n1018), .ZN(new_n1019));
  NOR2_X1   g833(.A1(new_n1015), .A2(new_n1019), .ZN(G72));
  NAND2_X1  g834(.A1(G472), .A2(G902), .ZN(new_n1021));
  XOR2_X1   g835(.A(new_n1021), .B(KEYINPUT63), .Z(new_n1022));
  OAI21_X1  g836(.A(new_n1022), .B1(new_n996), .B2(new_n885), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n936), .B1(new_n1023), .B2(new_n714), .ZN(new_n1024));
  INV_X1    g838(.A(new_n430), .ZN(new_n1025));
  OAI211_X1 g839(.A(new_n907), .B(new_n1022), .C1(new_n1025), .C2(new_n466), .ZN(new_n1026));
  INV_X1    g840(.A(new_n1010), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n1022), .B1(new_n1027), .B2(new_n885), .ZN(new_n1028));
  NOR2_X1   g842(.A1(new_n460), .A2(new_n427), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  AND3_X1   g844(.A1(new_n1024), .A2(new_n1026), .A3(new_n1030), .ZN(G57));
endmodule


