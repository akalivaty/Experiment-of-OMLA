

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594;

  XNOR2_X1 U325 ( .A(n440), .B(KEYINPUT55), .ZN(n456) );
  XNOR2_X1 U326 ( .A(n319), .B(n308), .ZN(n563) );
  XOR2_X1 U327 ( .A(n334), .B(n333), .Z(n293) );
  INV_X1 U328 ( .A(KEYINPUT115), .ZN(n371) );
  XNOR2_X1 U329 ( .A(n371), .B(KEYINPUT45), .ZN(n372) );
  XNOR2_X1 U330 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U331 ( .A(n368), .B(KEYINPUT114), .ZN(n369) );
  XOR2_X1 U332 ( .A(G218GAT), .B(G162GAT), .Z(n425) );
  XNOR2_X1 U333 ( .A(n370), .B(n369), .ZN(n378) );
  XNOR2_X1 U334 ( .A(n335), .B(n293), .ZN(n336) );
  XNOR2_X1 U335 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U336 ( .A(n585), .B(KEYINPUT41), .Z(n570) );
  INV_X1 U337 ( .A(G190GAT), .ZN(n459) );
  INV_X1 U338 ( .A(G183GAT), .ZN(n462) );
  XNOR2_X1 U339 ( .A(n459), .B(KEYINPUT58), .ZN(n460) );
  XNOR2_X1 U340 ( .A(n461), .B(n460), .ZN(G1351GAT) );
  XOR2_X1 U341 ( .A(KEYINPUT7), .B(G50GAT), .Z(n295) );
  XNOR2_X1 U342 ( .A(G36GAT), .B(G29GAT), .ZN(n294) );
  XNOR2_X1 U343 ( .A(n295), .B(n294), .ZN(n296) );
  XNOR2_X1 U344 ( .A(KEYINPUT8), .B(n296), .ZN(n319) );
  XNOR2_X1 U345 ( .A(G85GAT), .B(G92GAT), .ZN(n321) );
  XNOR2_X1 U346 ( .A(n425), .B(n321), .ZN(n298) );
  NAND2_X1 U347 ( .A1(G232GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U348 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U349 ( .A(KEYINPUT9), .B(G106GAT), .Z(n300) );
  XNOR2_X1 U350 ( .A(G43GAT), .B(G99GAT), .ZN(n299) );
  XNOR2_X1 U351 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U352 ( .A(n302), .B(n301), .ZN(n307) );
  XOR2_X1 U353 ( .A(G190GAT), .B(G134GAT), .Z(n442) );
  XOR2_X1 U354 ( .A(KEYINPUT10), .B(KEYINPUT70), .Z(n304) );
  XNOR2_X1 U355 ( .A(KEYINPUT71), .B(KEYINPUT11), .ZN(n303) );
  XNOR2_X1 U356 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U357 ( .A(n442), .B(n305), .ZN(n306) );
  XNOR2_X1 U358 ( .A(n307), .B(n306), .ZN(n308) );
  INV_X1 U359 ( .A(n563), .ZN(n458) );
  XOR2_X1 U360 ( .A(G15GAT), .B(G113GAT), .Z(n310) );
  XNOR2_X1 U361 ( .A(G169GAT), .B(G43GAT), .ZN(n309) );
  XNOR2_X1 U362 ( .A(n310), .B(n309), .ZN(n451) );
  XOR2_X1 U363 ( .A(n451), .B(KEYINPUT29), .Z(n312) );
  NAND2_X1 U364 ( .A1(G229GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U365 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U366 ( .A(KEYINPUT65), .B(KEYINPUT64), .Z(n314) );
  XNOR2_X1 U367 ( .A(G197GAT), .B(KEYINPUT30), .ZN(n313) );
  XNOR2_X1 U368 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U369 ( .A(n316), .B(n315), .Z(n318) );
  XOR2_X1 U370 ( .A(G141GAT), .B(G22GAT), .Z(n426) );
  XOR2_X1 U371 ( .A(G8GAT), .B(G1GAT), .Z(n342) );
  XNOR2_X1 U372 ( .A(n426), .B(n342), .ZN(n317) );
  XNOR2_X1 U373 ( .A(n318), .B(n317), .ZN(n320) );
  XOR2_X1 U374 ( .A(n320), .B(n319), .Z(n554) );
  INV_X1 U375 ( .A(n554), .ZN(n580) );
  XNOR2_X1 U376 ( .A(G176GAT), .B(KEYINPUT31), .ZN(n322) );
  XNOR2_X1 U377 ( .A(n322), .B(n321), .ZN(n339) );
  XNOR2_X1 U378 ( .A(G99GAT), .B(G71GAT), .ZN(n323) );
  XNOR2_X1 U379 ( .A(n323), .B(G120GAT), .ZN(n441) );
  NAND2_X1 U380 ( .A1(n441), .A2(KEYINPUT32), .ZN(n327) );
  INV_X1 U381 ( .A(n441), .ZN(n325) );
  INV_X1 U382 ( .A(KEYINPUT32), .ZN(n324) );
  NAND2_X1 U383 ( .A1(n325), .A2(n324), .ZN(n326) );
  NAND2_X1 U384 ( .A1(n327), .A2(n326), .ZN(n329) );
  AND2_X1 U385 ( .A1(G230GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U386 ( .A(n329), .B(n328), .ZN(n337) );
  XOR2_X1 U387 ( .A(G78GAT), .B(G148GAT), .Z(n331) );
  XNOR2_X1 U388 ( .A(G106GAT), .B(G204GAT), .ZN(n330) );
  XNOR2_X1 U389 ( .A(n331), .B(n330), .ZN(n421) );
  XNOR2_X1 U390 ( .A(G57GAT), .B(G64GAT), .ZN(n332) );
  XNOR2_X1 U391 ( .A(n332), .B(KEYINPUT13), .ZN(n343) );
  XNOR2_X1 U392 ( .A(n421), .B(n343), .ZN(n335) );
  XOR2_X1 U393 ( .A(KEYINPUT67), .B(KEYINPUT33), .Z(n334) );
  XNOR2_X1 U394 ( .A(KEYINPUT69), .B(KEYINPUT68), .ZN(n333) );
  XOR2_X1 U395 ( .A(n339), .B(n338), .Z(n585) );
  NOR2_X1 U396 ( .A1(n580), .A2(n570), .ZN(n341) );
  XNOR2_X1 U397 ( .A(KEYINPUT46), .B(KEYINPUT113), .ZN(n340) );
  XNOR2_X1 U398 ( .A(n341), .B(n340), .ZN(n367) );
  XOR2_X1 U399 ( .A(n343), .B(n342), .Z(n345) );
  NAND2_X1 U400 ( .A1(G231GAT), .A2(G233GAT), .ZN(n344) );
  XNOR2_X1 U401 ( .A(n345), .B(n344), .ZN(n349) );
  XOR2_X1 U402 ( .A(KEYINPUT74), .B(KEYINPUT73), .Z(n347) );
  XNOR2_X1 U403 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n346) );
  XNOR2_X1 U404 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U405 ( .A(n349), .B(n348), .ZN(n353) );
  XOR2_X1 U406 ( .A(KEYINPUT77), .B(KEYINPUT75), .Z(n351) );
  XNOR2_X1 U407 ( .A(KEYINPUT72), .B(KEYINPUT76), .ZN(n350) );
  XNOR2_X1 U408 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U409 ( .A(n353), .B(n352), .ZN(n357) );
  XOR2_X1 U410 ( .A(G71GAT), .B(G127GAT), .Z(n355) );
  XNOR2_X1 U411 ( .A(G15GAT), .B(G183GAT), .ZN(n354) );
  XNOR2_X1 U412 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U413 ( .A(n357), .B(n356), .ZN(n365) );
  XOR2_X1 U414 ( .A(KEYINPUT80), .B(KEYINPUT79), .Z(n359) );
  XNOR2_X1 U415 ( .A(KEYINPUT78), .B(KEYINPUT12), .ZN(n358) );
  XNOR2_X1 U416 ( .A(n359), .B(n358), .ZN(n363) );
  XOR2_X1 U417 ( .A(G155GAT), .B(G78GAT), .Z(n361) );
  XNOR2_X1 U418 ( .A(G22GAT), .B(G211GAT), .ZN(n360) );
  XNOR2_X1 U419 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U420 ( .A(n363), .B(n362), .Z(n364) );
  XNOR2_X1 U421 ( .A(n365), .B(n364), .ZN(n588) );
  INV_X1 U422 ( .A(n588), .ZN(n561) );
  NOR2_X1 U423 ( .A1(n563), .A2(n561), .ZN(n366) );
  AND2_X1 U424 ( .A1(n367), .A2(n366), .ZN(n370) );
  INV_X1 U425 ( .A(KEYINPUT47), .ZN(n368) );
  XOR2_X1 U426 ( .A(KEYINPUT66), .B(n580), .Z(n566) );
  XOR2_X1 U427 ( .A(n563), .B(KEYINPUT36), .Z(n591) );
  NOR2_X1 U428 ( .A1(n588), .A2(n591), .ZN(n373) );
  NAND2_X1 U429 ( .A1(n374), .A2(n585), .ZN(n375) );
  NOR2_X1 U430 ( .A1(n566), .A2(n375), .ZN(n376) );
  XNOR2_X1 U431 ( .A(KEYINPUT116), .B(n376), .ZN(n377) );
  NOR2_X1 U432 ( .A1(n378), .A2(n377), .ZN(n379) );
  XNOR2_X1 U433 ( .A(KEYINPUT48), .B(n379), .ZN(n537) );
  XNOR2_X1 U434 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n380) );
  XNOR2_X1 U435 ( .A(n380), .B(G211GAT), .ZN(n422) );
  XOR2_X1 U436 ( .A(G218GAT), .B(n422), .Z(n382) );
  NAND2_X1 U437 ( .A1(G226GAT), .A2(G233GAT), .ZN(n381) );
  XNOR2_X1 U438 ( .A(n382), .B(n381), .ZN(n386) );
  XOR2_X1 U439 ( .A(KEYINPUT96), .B(G64GAT), .Z(n384) );
  XNOR2_X1 U440 ( .A(G8GAT), .B(KEYINPUT72), .ZN(n383) );
  XNOR2_X1 U441 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U442 ( .A(n386), .B(n385), .Z(n391) );
  XOR2_X1 U443 ( .A(G92GAT), .B(G204GAT), .Z(n388) );
  XNOR2_X1 U444 ( .A(G169GAT), .B(G36GAT), .ZN(n387) );
  XNOR2_X1 U445 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U446 ( .A(G190GAT), .B(n389), .ZN(n390) );
  XNOR2_X1 U447 ( .A(n391), .B(n390), .ZN(n396) );
  XOR2_X1 U448 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n393) );
  XNOR2_X1 U449 ( .A(G183GAT), .B(G176GAT), .ZN(n392) );
  XNOR2_X1 U450 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U451 ( .A(KEYINPUT18), .B(n394), .ZN(n446) );
  INV_X1 U452 ( .A(n446), .ZN(n395) );
  XOR2_X1 U453 ( .A(n396), .B(n395), .Z(n526) );
  NOR2_X1 U454 ( .A1(n537), .A2(n526), .ZN(n398) );
  INV_X1 U455 ( .A(KEYINPUT54), .ZN(n397) );
  XNOR2_X1 U456 ( .A(n398), .B(n397), .ZN(n575) );
  XOR2_X1 U457 ( .A(KEYINPUT1), .B(KEYINPUT95), .Z(n400) );
  XNOR2_X1 U458 ( .A(KEYINPUT93), .B(KEYINPUT94), .ZN(n399) );
  XNOR2_X1 U459 ( .A(n400), .B(n399), .ZN(n412) );
  XOR2_X1 U460 ( .A(G57GAT), .B(G148GAT), .Z(n402) );
  XNOR2_X1 U461 ( .A(G141GAT), .B(G1GAT), .ZN(n401) );
  XNOR2_X1 U462 ( .A(n402), .B(n401), .ZN(n406) );
  XOR2_X1 U463 ( .A(KEYINPUT6), .B(KEYINPUT92), .Z(n404) );
  XNOR2_X1 U464 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(n403) );
  XNOR2_X1 U465 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U466 ( .A(n406), .B(n405), .Z(n410) );
  XNOR2_X1 U467 ( .A(G127GAT), .B(KEYINPUT82), .ZN(n407) );
  XNOR2_X1 U468 ( .A(n407), .B(KEYINPUT0), .ZN(n450) );
  XNOR2_X1 U469 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n408) );
  XNOR2_X1 U470 ( .A(n408), .B(KEYINPUT2), .ZN(n434) );
  XNOR2_X1 U471 ( .A(n450), .B(n434), .ZN(n409) );
  XNOR2_X1 U472 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U473 ( .A(n412), .B(n411), .ZN(n420) );
  NAND2_X1 U474 ( .A1(G225GAT), .A2(G233GAT), .ZN(n418) );
  XOR2_X1 U475 ( .A(G85GAT), .B(G162GAT), .Z(n414) );
  XNOR2_X1 U476 ( .A(G113GAT), .B(G120GAT), .ZN(n413) );
  XNOR2_X1 U477 ( .A(n414), .B(n413), .ZN(n416) );
  XOR2_X1 U478 ( .A(G29GAT), .B(G134GAT), .Z(n415) );
  XNOR2_X1 U479 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U480 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U481 ( .A(n420), .B(n419), .Z(n524) );
  XNOR2_X1 U482 ( .A(n422), .B(n421), .ZN(n438) );
  XOR2_X1 U483 ( .A(KEYINPUT23), .B(KEYINPUT90), .Z(n424) );
  XNOR2_X1 U484 ( .A(KEYINPUT89), .B(KEYINPUT88), .ZN(n423) );
  XNOR2_X1 U485 ( .A(n424), .B(n423), .ZN(n430) );
  XOR2_X1 U486 ( .A(KEYINPUT22), .B(n425), .Z(n428) );
  XNOR2_X1 U487 ( .A(G50GAT), .B(n426), .ZN(n427) );
  XNOR2_X1 U488 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U489 ( .A(n430), .B(n429), .Z(n432) );
  NAND2_X1 U490 ( .A1(G228GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U491 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U492 ( .A(n433), .B(KEYINPUT24), .Z(n436) );
  XNOR2_X1 U493 ( .A(n434), .B(KEYINPUT91), .ZN(n435) );
  XNOR2_X1 U494 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U495 ( .A(n438), .B(n437), .ZN(n472) );
  NAND2_X1 U496 ( .A1(n524), .A2(n472), .ZN(n439) );
  OR2_X1 U497 ( .A1(n575), .A2(n439), .ZN(n440) );
  XOR2_X1 U498 ( .A(n441), .B(KEYINPUT85), .Z(n444) );
  XNOR2_X1 U499 ( .A(n442), .B(KEYINPUT86), .ZN(n443) );
  XNOR2_X1 U500 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U501 ( .A(n446), .B(n445), .Z(n455) );
  XOR2_X1 U502 ( .A(KEYINPUT84), .B(KEYINPUT83), .Z(n448) );
  NAND2_X1 U503 ( .A1(G227GAT), .A2(G233GAT), .ZN(n447) );
  XNOR2_X1 U504 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U505 ( .A(n449), .B(KEYINPUT20), .Z(n453) );
  XNOR2_X1 U506 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U507 ( .A(n453), .B(n452), .ZN(n454) );
  XOR2_X1 U508 ( .A(n455), .B(n454), .Z(n539) );
  INV_X1 U509 ( .A(n539), .ZN(n505) );
  NAND2_X1 U510 ( .A1(n456), .A2(n505), .ZN(n457) );
  XNOR2_X1 U511 ( .A(n457), .B(KEYINPUT122), .ZN(n571) );
  NOR2_X1 U512 ( .A1(n458), .A2(n571), .ZN(n461) );
  NOR2_X1 U513 ( .A1(n588), .A2(n571), .ZN(n464) );
  XNOR2_X1 U514 ( .A(n462), .B(KEYINPUT124), .ZN(n463) );
  XNOR2_X1 U515 ( .A(n464), .B(n463), .ZN(G1350GAT) );
  AND2_X1 U516 ( .A1(n585), .A2(n566), .ZN(n496) );
  XOR2_X1 U517 ( .A(n539), .B(KEYINPUT87), .Z(n467) );
  XNOR2_X1 U518 ( .A(n472), .B(KEYINPUT28), .ZN(n533) );
  INV_X1 U519 ( .A(n533), .ZN(n538) );
  INV_X1 U520 ( .A(n526), .ZN(n503) );
  XOR2_X1 U521 ( .A(n503), .B(KEYINPUT97), .Z(n465) );
  XNOR2_X1 U522 ( .A(n465), .B(KEYINPUT27), .ZN(n469) );
  INV_X1 U523 ( .A(n524), .ZN(n576) );
  NAND2_X1 U524 ( .A1(n469), .A2(n576), .ZN(n536) );
  NOR2_X1 U525 ( .A1(n538), .A2(n536), .ZN(n466) );
  NAND2_X1 U526 ( .A1(n467), .A2(n466), .ZN(n478) );
  NOR2_X1 U527 ( .A1(n472), .A2(n505), .ZN(n468) );
  XNOR2_X1 U528 ( .A(n468), .B(KEYINPUT26), .ZN(n577) );
  NAND2_X1 U529 ( .A1(n577), .A2(n469), .ZN(n475) );
  NOR2_X1 U530 ( .A1(n526), .A2(n539), .ZN(n470) );
  XOR2_X1 U531 ( .A(KEYINPUT98), .B(n470), .Z(n471) );
  NAND2_X1 U532 ( .A1(n472), .A2(n471), .ZN(n473) );
  XOR2_X1 U533 ( .A(KEYINPUT25), .B(n473), .Z(n474) );
  NAND2_X1 U534 ( .A1(n475), .A2(n474), .ZN(n476) );
  NAND2_X1 U535 ( .A1(n476), .A2(n524), .ZN(n477) );
  NAND2_X1 U536 ( .A1(n478), .A2(n477), .ZN(n493) );
  NOR2_X1 U537 ( .A1(n563), .A2(n588), .ZN(n479) );
  XNOR2_X1 U538 ( .A(n479), .B(KEYINPUT16), .ZN(n480) );
  XOR2_X1 U539 ( .A(KEYINPUT81), .B(n480), .Z(n481) );
  AND2_X1 U540 ( .A1(n493), .A2(n481), .ZN(n511) );
  NAND2_X1 U541 ( .A1(n496), .A2(n511), .ZN(n490) );
  NOR2_X1 U542 ( .A1(n524), .A2(n490), .ZN(n483) );
  XNOR2_X1 U543 ( .A(KEYINPUT34), .B(KEYINPUT99), .ZN(n482) );
  XNOR2_X1 U544 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U545 ( .A(G1GAT), .B(n484), .ZN(G1324GAT) );
  NOR2_X1 U546 ( .A1(n526), .A2(n490), .ZN(n485) );
  XOR2_X1 U547 ( .A(KEYINPUT100), .B(n485), .Z(n486) );
  XNOR2_X1 U548 ( .A(G8GAT), .B(n486), .ZN(G1325GAT) );
  NOR2_X1 U549 ( .A1(n539), .A2(n490), .ZN(n488) );
  XNOR2_X1 U550 ( .A(KEYINPUT101), .B(KEYINPUT35), .ZN(n487) );
  XNOR2_X1 U551 ( .A(n488), .B(n487), .ZN(n489) );
  XOR2_X1 U552 ( .A(G15GAT), .B(n489), .Z(G1326GAT) );
  NOR2_X1 U553 ( .A1(n533), .A2(n490), .ZN(n491) );
  XOR2_X1 U554 ( .A(KEYINPUT102), .B(n491), .Z(n492) );
  XNOR2_X1 U555 ( .A(G22GAT), .B(n492), .ZN(G1327GAT) );
  XOR2_X1 U556 ( .A(KEYINPUT38), .B(KEYINPUT104), .Z(n498) );
  NAND2_X1 U557 ( .A1(n588), .A2(n493), .ZN(n494) );
  NOR2_X1 U558 ( .A1(n591), .A2(n494), .ZN(n495) );
  XOR2_X1 U559 ( .A(KEYINPUT37), .B(n495), .Z(n523) );
  NAND2_X1 U560 ( .A1(n496), .A2(n523), .ZN(n497) );
  XNOR2_X1 U561 ( .A(n498), .B(n497), .ZN(n508) );
  NAND2_X1 U562 ( .A1(n576), .A2(n508), .ZN(n502) );
  XOR2_X1 U563 ( .A(KEYINPUT105), .B(KEYINPUT39), .Z(n500) );
  XNOR2_X1 U564 ( .A(G29GAT), .B(KEYINPUT103), .ZN(n499) );
  XNOR2_X1 U565 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U566 ( .A(n502), .B(n501), .ZN(G1328GAT) );
  NAND2_X1 U567 ( .A1(n508), .A2(n503), .ZN(n504) );
  XNOR2_X1 U568 ( .A(G36GAT), .B(n504), .ZN(G1329GAT) );
  NAND2_X1 U569 ( .A1(n508), .A2(n505), .ZN(n506) );
  XNOR2_X1 U570 ( .A(n506), .B(KEYINPUT40), .ZN(n507) );
  XNOR2_X1 U571 ( .A(G43GAT), .B(n507), .ZN(G1330GAT) );
  NAND2_X1 U572 ( .A1(n508), .A2(n538), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n509), .B(KEYINPUT106), .ZN(n510) );
  XNOR2_X1 U574 ( .A(G50GAT), .B(n510), .ZN(G1331GAT) );
  NOR2_X1 U575 ( .A1(n554), .A2(n570), .ZN(n522) );
  NAND2_X1 U576 ( .A1(n522), .A2(n511), .ZN(n518) );
  NOR2_X1 U577 ( .A1(n524), .A2(n518), .ZN(n512) );
  XOR2_X1 U578 ( .A(G57GAT), .B(n512), .Z(n513) );
  XNOR2_X1 U579 ( .A(KEYINPUT42), .B(n513), .ZN(G1332GAT) );
  NOR2_X1 U580 ( .A1(n526), .A2(n518), .ZN(n515) );
  XNOR2_X1 U581 ( .A(G64GAT), .B(KEYINPUT107), .ZN(n514) );
  XNOR2_X1 U582 ( .A(n515), .B(n514), .ZN(G1333GAT) );
  NOR2_X1 U583 ( .A1(n539), .A2(n518), .ZN(n516) );
  XOR2_X1 U584 ( .A(KEYINPUT108), .B(n516), .Z(n517) );
  XNOR2_X1 U585 ( .A(G71GAT), .B(n517), .ZN(G1334GAT) );
  NOR2_X1 U586 ( .A1(n533), .A2(n518), .ZN(n520) );
  XNOR2_X1 U587 ( .A(KEYINPUT109), .B(KEYINPUT43), .ZN(n519) );
  XNOR2_X1 U588 ( .A(n520), .B(n519), .ZN(n521) );
  XOR2_X1 U589 ( .A(G78GAT), .B(n521), .Z(G1335GAT) );
  NAND2_X1 U590 ( .A1(n523), .A2(n522), .ZN(n532) );
  NOR2_X1 U591 ( .A1(n524), .A2(n532), .ZN(n525) );
  XOR2_X1 U592 ( .A(G85GAT), .B(n525), .Z(G1336GAT) );
  NOR2_X1 U593 ( .A1(n526), .A2(n532), .ZN(n528) );
  XNOR2_X1 U594 ( .A(KEYINPUT110), .B(KEYINPUT111), .ZN(n527) );
  XNOR2_X1 U595 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U596 ( .A(G92GAT), .B(n529), .ZN(G1337GAT) );
  NOR2_X1 U597 ( .A1(n539), .A2(n532), .ZN(n530) );
  XOR2_X1 U598 ( .A(KEYINPUT112), .B(n530), .Z(n531) );
  XNOR2_X1 U599 ( .A(G99GAT), .B(n531), .ZN(G1338GAT) );
  NOR2_X1 U600 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U601 ( .A(G106GAT), .B(n534), .Z(n535) );
  XNOR2_X1 U602 ( .A(KEYINPUT44), .B(n535), .ZN(G1339GAT) );
  NOR2_X1 U603 ( .A1(n537), .A2(n536), .ZN(n552) );
  NOR2_X1 U604 ( .A1(n539), .A2(n538), .ZN(n540) );
  NAND2_X1 U605 ( .A1(n552), .A2(n540), .ZN(n541) );
  XNOR2_X1 U606 ( .A(KEYINPUT117), .B(n541), .ZN(n549) );
  NAND2_X1 U607 ( .A1(n549), .A2(n566), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n542), .B(KEYINPUT118), .ZN(n543) );
  XNOR2_X1 U609 ( .A(G113GAT), .B(n543), .ZN(G1340GAT) );
  XOR2_X1 U610 ( .A(G120GAT), .B(KEYINPUT49), .Z(n545) );
  INV_X1 U611 ( .A(n570), .ZN(n556) );
  NAND2_X1 U612 ( .A1(n549), .A2(n556), .ZN(n544) );
  XNOR2_X1 U613 ( .A(n545), .B(n544), .ZN(G1341GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT119), .B(KEYINPUT50), .Z(n547) );
  NAND2_X1 U615 ( .A1(n549), .A2(n561), .ZN(n546) );
  XNOR2_X1 U616 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U617 ( .A(G127GAT), .B(n548), .ZN(G1342GAT) );
  XOR2_X1 U618 ( .A(G134GAT), .B(KEYINPUT51), .Z(n551) );
  NAND2_X1 U619 ( .A1(n549), .A2(n563), .ZN(n550) );
  XNOR2_X1 U620 ( .A(n551), .B(n550), .ZN(G1343GAT) );
  NAND2_X1 U621 ( .A1(n577), .A2(n552), .ZN(n553) );
  XOR2_X1 U622 ( .A(KEYINPUT120), .B(n553), .Z(n564) );
  NAND2_X1 U623 ( .A1(n554), .A2(n564), .ZN(n555) );
  XNOR2_X1 U624 ( .A(G141GAT), .B(n555), .ZN(G1344GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT121), .B(KEYINPUT52), .Z(n558) );
  NAND2_X1 U626 ( .A1(n556), .A2(n564), .ZN(n557) );
  XNOR2_X1 U627 ( .A(n558), .B(n557), .ZN(n560) );
  XOR2_X1 U628 ( .A(G148GAT), .B(KEYINPUT53), .Z(n559) );
  XNOR2_X1 U629 ( .A(n560), .B(n559), .ZN(G1345GAT) );
  NAND2_X1 U630 ( .A1(n564), .A2(n561), .ZN(n562) );
  XNOR2_X1 U631 ( .A(n562), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U632 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n565), .B(G162GAT), .ZN(G1347GAT) );
  INV_X1 U634 ( .A(n566), .ZN(n567) );
  NOR2_X1 U635 ( .A1(n571), .A2(n567), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n568), .B(KEYINPUT123), .ZN(n569) );
  XNOR2_X1 U637 ( .A(G169GAT), .B(n569), .ZN(G1348GAT) );
  NOR2_X1 U638 ( .A1(n571), .A2(n570), .ZN(n573) );
  XNOR2_X1 U639 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n572) );
  XNOR2_X1 U640 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U641 ( .A(G176GAT), .B(n574), .ZN(G1349GAT) );
  NOR2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n578) );
  NAND2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U644 ( .A(KEYINPUT125), .B(n579), .Z(n590) );
  NOR2_X1 U645 ( .A1(n580), .A2(n590), .ZN(n584) );
  XNOR2_X1 U646 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n581), .B(KEYINPUT60), .ZN(n582) );
  XNOR2_X1 U648 ( .A(KEYINPUT126), .B(n582), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1352GAT) );
  NOR2_X1 U650 ( .A1(n585), .A2(n590), .ZN(n587) );
  XNOR2_X1 U651 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(G1353GAT) );
  NOR2_X1 U653 ( .A1(n588), .A2(n590), .ZN(n589) );
  XOR2_X1 U654 ( .A(G211GAT), .B(n589), .Z(G1354GAT) );
  NOR2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n593) );
  XNOR2_X1 U656 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n592) );
  XNOR2_X1 U657 ( .A(n593), .B(n592), .ZN(n594) );
  XNOR2_X1 U658 ( .A(G218GAT), .B(n594), .ZN(G1355GAT) );
endmodule

