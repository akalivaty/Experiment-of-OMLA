//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 1 0 1 0 1 0 1 0 0 1 0 0 0 1 0 1 1 0 1 0 1 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 0 0 0 1 0 0 1 0 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n757, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n846, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n906, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947;
  XNOR2_X1  g000(.A(G15gat), .B(G43gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G71gat), .B(G99gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT26), .ZN(new_n205));
  INV_X1    g004(.A(G169gat), .ZN(new_n206));
  INV_X1    g005(.A(G176gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G183gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT27), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT27), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G183gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT66), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI21_X1  g020(.A(G190gat), .B1(new_n216), .B2(KEYINPUT66), .ZN(new_n222));
  AOI21_X1  g021(.A(KEYINPUT28), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT28), .ZN(new_n224));
  NOR3_X1   g023(.A1(new_n219), .A2(new_n224), .A3(G190gat), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n214), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n212), .A2(KEYINPUT65), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT65), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n228), .A2(G183gat), .A3(G190gat), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT24), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n227), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(G190gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n215), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n231), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n206), .A2(new_n207), .A3(KEYINPUT23), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT23), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n237), .B1(G169gat), .B2(G176gat), .ZN(new_n238));
  AND4_X1   g037(.A1(KEYINPUT25), .A2(new_n236), .A3(new_n238), .A4(new_n210), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n235), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n212), .A2(new_n230), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n242), .A2(new_n233), .A3(new_n234), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n236), .A2(new_n238), .A3(new_n210), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n241), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n240), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n226), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT70), .ZN(new_n250));
  AND2_X1   g049(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n251));
  NOR2_X1   g050(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n252));
  INV_X1    g051(.A(G120gat), .ZN(new_n253));
  NOR3_X1   g052(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(G113gat), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n255), .A2(G120gat), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n250), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n253), .A2(G113gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(KEYINPUT69), .B(G113gat), .ZN(new_n259));
  OAI211_X1 g058(.A(KEYINPUT70), .B(new_n258), .C1(new_n259), .C2(new_n253), .ZN(new_n260));
  INV_X1    g059(.A(G127gat), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n261), .A2(G134gat), .ZN(new_n262));
  INV_X1    g061(.A(G134gat), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n263), .A2(G127gat), .ZN(new_n264));
  NOR3_X1   g063(.A1(new_n262), .A2(new_n264), .A3(KEYINPUT1), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n257), .A2(new_n260), .A3(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT1), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n255), .A2(G120gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n258), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G127gat), .B(G134gat), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT67), .ZN(new_n271));
  AOI22_X1  g070(.A1(new_n267), .A2(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(KEYINPUT67), .B1(new_n262), .B2(new_n264), .ZN(new_n273));
  AOI21_X1  g072(.A(KEYINPUT68), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n253), .A2(G113gat), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n267), .B1(new_n256), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n263), .A2(G127gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n261), .A2(G134gat), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n277), .A2(new_n278), .A3(new_n271), .ZN(new_n279));
  AND4_X1   g078(.A1(KEYINPUT68), .A2(new_n273), .A3(new_n276), .A4(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n266), .B1(new_n274), .B2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT71), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT68), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n276), .A2(new_n279), .ZN(new_n285));
  INV_X1    g084(.A(new_n273), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n272), .A2(KEYINPUT68), .A3(new_n273), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT71), .B1(new_n289), .B2(new_n266), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n249), .B1(new_n283), .B2(new_n290), .ZN(new_n291));
  AND2_X1   g090(.A1(G227gat), .A2(G233gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n281), .A2(new_n282), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n289), .A2(KEYINPUT71), .A3(new_n266), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n293), .A2(new_n294), .A3(new_n248), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n291), .A2(new_n292), .A3(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT33), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n204), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT72), .ZN(new_n299));
  AND3_X1   g098(.A1(new_n296), .A2(new_n299), .A3(KEYINPUT32), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n299), .B1(new_n296), .B2(KEYINPUT32), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n298), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT34), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n296), .A2(KEYINPUT32), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n204), .A2(new_n297), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  AND3_X1   g106(.A1(new_n302), .A2(new_n303), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n303), .B1(new_n302), .B2(new_n307), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n292), .B1(new_n291), .B2(new_n295), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NOR3_X1   g110(.A1(new_n308), .A2(new_n309), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n313));
  INV_X1    g112(.A(new_n204), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n301), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n296), .A2(new_n299), .A3(KEYINPUT32), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(KEYINPUT34), .B1(new_n318), .B2(new_n306), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n302), .A2(new_n303), .A3(new_n307), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n310), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n312), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT75), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n243), .A2(new_n210), .A3(new_n236), .A4(new_n238), .ZN(new_n324));
  AOI22_X1  g123(.A1(new_n324), .A2(new_n241), .B1(new_n235), .B2(new_n239), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT66), .B1(new_n216), .B2(new_n218), .ZN(new_n326));
  OAI21_X1  g125(.A(KEYINPUT66), .B1(new_n217), .B2(G183gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(new_n232), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n224), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n219), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n330), .A2(KEYINPUT28), .A3(new_n232), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n213), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(G226gat), .A2(G233gat), .ZN(new_n333));
  NOR3_X1   g132(.A1(new_n325), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(KEYINPUT74), .B1(new_n325), .B2(new_n332), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT74), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n226), .A2(new_n247), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n333), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n339), .A2(KEYINPUT29), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n334), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  XOR2_X1   g140(.A(G197gat), .B(G204gat), .Z(new_n342));
  AOI21_X1  g141(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  XOR2_X1   g143(.A(G211gat), .B(G218gat), .Z(new_n345));
  OR3_X1    g144(.A1(new_n344), .A2(KEYINPUT73), .A3(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n345), .B1(new_n344), .B2(KEYINPUT73), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  OR2_X1    g147(.A1(new_n341), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n335), .A2(new_n337), .A3(new_n339), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n248), .A2(new_n340), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n350), .A2(new_n348), .A3(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(G8gat), .B(G36gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n353), .B(G64gat), .ZN(new_n354));
  INV_X1    g153(.A(G92gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n354), .B(new_n355), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n349), .A2(KEYINPUT30), .A3(new_n352), .A4(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n356), .B1(new_n349), .B2(new_n352), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n323), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n359), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n361), .A2(KEYINPUT75), .A3(new_n357), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n349), .A2(new_n352), .A3(new_n356), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT30), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n360), .A2(new_n362), .A3(new_n365), .ZN(new_n366));
  XOR2_X1   g165(.A(KEYINPUT76), .B(KEYINPUT0), .Z(new_n367));
  XNOR2_X1  g166(.A(G1gat), .B(G29gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n367), .B(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(G57gat), .B(G85gat), .ZN(new_n370));
  XOR2_X1   g169(.A(new_n369), .B(new_n370), .Z(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  XNOR2_X1  g171(.A(G141gat), .B(G148gat), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(G155gat), .ZN(new_n375));
  INV_X1    g174(.A(G162gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(G155gat), .A2(G162gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(KEYINPUT2), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n374), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n378), .B(new_n377), .C1(new_n373), .C2(KEYINPUT2), .ZN(new_n382));
  AND2_X1   g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n293), .A2(KEYINPUT4), .A3(new_n294), .A4(new_n383), .ZN(new_n384));
  OAI211_X1 g183(.A(new_n383), .B(new_n266), .C1(new_n274), .C2(new_n280), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT4), .ZN(new_n386));
  NAND2_X1  g185(.A1(G225gat), .A2(G233gat), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n385), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT3), .ZN(new_n390));
  AND3_X1   g189(.A1(new_n381), .A2(new_n382), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n390), .B1(new_n381), .B2(new_n382), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(new_n281), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n384), .A2(new_n389), .A3(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT5), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n382), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n281), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(new_n385), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n396), .B1(new_n399), .B2(new_n388), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n395), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT78), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n394), .A2(new_n396), .A3(new_n387), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n385), .A2(KEYINPUT4), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT77), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n385), .A2(KEYINPUT77), .A3(KEYINPUT4), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n293), .A2(new_n386), .A3(new_n294), .A4(new_n383), .ZN(new_n409));
  AOI211_X1 g208(.A(new_n402), .B(new_n403), .C1(new_n408), .C2(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT77), .B1(new_n385), .B2(KEYINPUT4), .ZN(new_n411));
  AND3_X1   g210(.A1(new_n385), .A2(KEYINPUT77), .A3(KEYINPUT4), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n409), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n403), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT78), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n372), .B(new_n401), .C1(new_n410), .C2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT6), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(KEYINPUT79), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n401), .B1(new_n410), .B2(new_n415), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(new_n371), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT79), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n416), .A2(new_n422), .A3(new_n417), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n419), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n420), .A2(KEYINPUT6), .A3(new_n371), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n366), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT29), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n427), .B1(new_n397), .B2(KEYINPUT3), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n348), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  OR2_X1    g229(.A1(new_n344), .A2(new_n345), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n344), .A2(new_n345), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n431), .A2(new_n427), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n383), .B1(new_n433), .B2(new_n390), .ZN(new_n434));
  INV_X1    g233(.A(G228gat), .ZN(new_n435));
  INV_X1    g234(.A(G233gat), .ZN(new_n436));
  OAI22_X1  g235(.A1(new_n430), .A2(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n435), .A2(new_n436), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n429), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n346), .A2(new_n427), .A3(new_n347), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n383), .B1(new_n440), .B2(new_n390), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n442), .A2(KEYINPUT81), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT81), .ZN(new_n444));
  NOR3_X1   g243(.A1(new_n439), .A2(new_n441), .A3(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n437), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(G22gat), .ZN(new_n447));
  INV_X1    g246(.A(G22gat), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n448), .B(new_n437), .C1(new_n443), .C2(new_n445), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g249(.A(G78gat), .B(G106gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n451), .B(KEYINPUT31), .ZN(new_n452));
  INV_X1    g251(.A(G50gat), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n452), .B(new_n453), .ZN(new_n454));
  XOR2_X1   g253(.A(new_n454), .B(KEYINPUT80), .Z(new_n455));
  NAND2_X1  g254(.A1(new_n450), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n442), .B(KEYINPUT81), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT82), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n457), .A2(new_n458), .A3(new_n448), .A4(new_n437), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n449), .A2(KEYINPUT82), .ZN(new_n460));
  INV_X1    g259(.A(new_n454), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n459), .A2(new_n460), .A3(new_n447), .A4(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n456), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n322), .A2(new_n426), .A3(KEYINPUT35), .A4(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n365), .A2(new_n361), .A3(new_n357), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n421), .A2(new_n417), .A3(new_n416), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n465), .B1(new_n466), .B2(new_n425), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n311), .B1(new_n308), .B2(new_n309), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n319), .A2(new_n310), .A3(new_n320), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n467), .A2(new_n468), .A3(new_n469), .A4(new_n463), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT35), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n464), .A2(new_n472), .ZN(new_n473));
  AND2_X1   g272(.A1(new_n456), .A2(new_n462), .ZN(new_n474));
  AND3_X1   g273(.A1(new_n420), .A2(KEYINPUT6), .A3(new_n371), .ZN(new_n475));
  AOI22_X1  g274(.A1(new_n418), .A2(KEYINPUT79), .B1(new_n371), .B2(new_n420), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n475), .B1(new_n476), .B2(new_n423), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n474), .B1(new_n477), .B2(new_n366), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n466), .A2(new_n425), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT37), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n352), .B(new_n480), .C1(new_n341), .C2(new_n348), .ZN(new_n481));
  INV_X1    g280(.A(new_n348), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n350), .A2(new_n482), .A3(new_n351), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n483), .B(KEYINPUT37), .C1(new_n341), .C2(new_n482), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT38), .ZN(new_n485));
  INV_X1    g284(.A(new_n356), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n481), .A2(new_n484), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT85), .ZN(new_n488));
  AND2_X1   g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n363), .B1(new_n487), .B2(new_n488), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT86), .B1(new_n479), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT86), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n466), .A2(new_n491), .A3(new_n494), .A4(new_n425), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT87), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n480), .B1(new_n349), .B2(new_n352), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n486), .ZN(new_n498));
  OR2_X1    g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n496), .B1(new_n499), .B2(KEYINPUT38), .ZN(new_n500));
  OAI211_X1 g299(.A(new_n496), .B(KEYINPUT38), .C1(new_n497), .C2(new_n498), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n493), .A2(new_n495), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n465), .A2(new_n421), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n387), .B1(new_n413), .B2(new_n394), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n398), .A2(new_n385), .A3(new_n387), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n507), .A2(KEYINPUT84), .ZN(new_n508));
  OAI21_X1  g307(.A(KEYINPUT39), .B1(new_n507), .B2(KEYINPUT84), .ZN(new_n509));
  OR3_X1    g308(.A1(new_n506), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  XOR2_X1   g309(.A(KEYINPUT83), .B(KEYINPUT39), .Z(new_n511));
  AOI21_X1  g310(.A(new_n371), .B1(new_n506), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(KEYINPUT40), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n505), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n510), .A2(KEYINPUT40), .A3(new_n512), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n474), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT36), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n517), .B1(new_n312), .B2(new_n321), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n468), .A2(new_n469), .A3(KEYINPUT36), .ZN(new_n519));
  AOI22_X1  g318(.A1(new_n504), .A2(new_n516), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n473), .B1(new_n478), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(G29gat), .A2(G36gat), .ZN(new_n522));
  OAI21_X1  g321(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  NOR3_X1   g323(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n522), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(G43gat), .B(G50gat), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n526), .A2(KEYINPUT15), .A3(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(KEYINPUT15), .ZN(new_n529));
  XOR2_X1   g328(.A(new_n522), .B(KEYINPUT90), .Z(new_n530));
  OR2_X1    g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT89), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n523), .B1(new_n525), .B2(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n533), .B1(new_n532), .B2(new_n525), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n528), .B1(new_n531), .B2(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(G15gat), .B(G22gat), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT16), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n536), .B1(new_n537), .B2(G1gat), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n538), .B1(G1gat), .B2(new_n536), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n539), .B(G8gat), .ZN(new_n540));
  OAI21_X1  g339(.A(KEYINPUT92), .B1(new_n535), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n535), .A2(new_n540), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(G229gat), .A2(G233gat), .ZN(new_n544));
  XOR2_X1   g343(.A(new_n544), .B(KEYINPUT13), .Z(new_n545));
  NAND2_X1  g344(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n535), .B(KEYINPUT17), .ZN(new_n547));
  INV_X1    g346(.A(new_n540), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n549), .A2(KEYINPUT18), .A3(new_n544), .A4(new_n542), .ZN(new_n550));
  XNOR2_X1  g349(.A(G169gat), .B(G197gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(G113gat), .B(G141gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  XOR2_X1   g352(.A(KEYINPUT88), .B(KEYINPUT11), .Z(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT12), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n546), .A2(new_n550), .A3(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n549), .A2(new_n544), .A3(new_n542), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(KEYINPUT91), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT18), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT91), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n549), .A2(new_n561), .A3(new_n544), .A4(new_n542), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n559), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n557), .B1(new_n563), .B2(KEYINPUT93), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT93), .ZN(new_n565));
  NAND4_X1  g364(.A1(new_n559), .A2(new_n565), .A3(new_n560), .A4(new_n562), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n563), .A2(new_n546), .A3(new_n550), .ZN(new_n567));
  INV_X1    g366(.A(new_n556), .ZN(new_n568));
  AOI22_X1  g367(.A1(new_n564), .A2(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G57gat), .B(G64gat), .ZN(new_n570));
  AOI21_X1  g369(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(G71gat), .B(G78gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(KEYINPUT95), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT21), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n548), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(new_n215), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n574), .A2(new_n576), .ZN(new_n579));
  NAND2_X1  g378(.A1(G231gat), .A2(G233gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  XOR2_X1   g380(.A(G127gat), .B(G155gat), .Z(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT94), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n581), .B(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n578), .B(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(G211gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n585), .B(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G190gat), .B(G218gat), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  XOR2_X1   g389(.A(G99gat), .B(G106gat), .Z(new_n591));
  INV_X1    g390(.A(G85gat), .ZN(new_n592));
  OAI21_X1  g391(.A(KEYINPUT7), .B1(new_n592), .B2(new_n355), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT7), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n594), .A2(G85gat), .A3(G92gat), .ZN(new_n595));
  AOI22_X1  g394(.A1(new_n591), .A2(KEYINPUT97), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(G99gat), .ZN(new_n597));
  INV_X1    g396(.A(G106gat), .ZN(new_n598));
  OAI21_X1  g397(.A(KEYINPUT8), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  XOR2_X1   g398(.A(KEYINPUT96), .B(G85gat), .Z(new_n600));
  OAI211_X1 g399(.A(new_n596), .B(new_n599), .C1(G92gat), .C2(new_n600), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n591), .A2(KEYINPUT97), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n547), .A2(new_n604), .ZN(new_n605));
  AND2_X1   g404(.A1(G232gat), .A2(G233gat), .ZN(new_n606));
  AOI22_X1  g405(.A1(new_n603), .A2(new_n535), .B1(KEYINPUT41), .B2(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n590), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n605), .A2(new_n590), .A3(new_n607), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g410(.A(G134gat), .B(G162gat), .Z(new_n612));
  NOR2_X1   g411(.A1(new_n606), .A2(KEYINPUT41), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n614), .B1(new_n608), .B2(KEYINPUT98), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n609), .A2(KEYINPUT98), .A3(new_n610), .A4(new_n614), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n588), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(G230gat), .A2(G233gat), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n604), .A2(new_n574), .ZN(new_n622));
  INV_X1    g421(.A(new_n574), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n603), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n621), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT99), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n621), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT10), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n622), .A2(new_n629), .A3(new_n624), .ZN(new_n630));
  OR3_X1    g429(.A1(new_n604), .A2(new_n629), .A3(new_n575), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n628), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(G120gat), .B(G148gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(G176gat), .ZN(new_n635));
  INV_X1    g434(.A(G204gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n627), .A2(new_n633), .A3(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n637), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n639), .B1(new_n632), .B2(new_n625), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT100), .ZN(new_n641));
  AND3_X1   g440(.A1(new_n638), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n641), .B1(new_n638), .B2(new_n640), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n620), .A2(new_n644), .ZN(new_n645));
  NOR3_X1   g444(.A1(new_n521), .A2(new_n569), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(new_n477), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g447(.A1(new_n646), .A2(new_n465), .ZN(new_n649));
  XOR2_X1   g448(.A(KEYINPUT16), .B(G8gat), .Z(new_n650));
  NAND3_X1  g449(.A1(new_n649), .A2(KEYINPUT42), .A3(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(G8gat), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n649), .A2(new_n650), .ZN(new_n653));
  XOR2_X1   g452(.A(KEYINPUT101), .B(KEYINPUT42), .Z(new_n654));
  AND3_X1   g453(.A1(new_n653), .A2(KEYINPUT102), .A3(new_n654), .ZN(new_n655));
  AOI21_X1  g454(.A(KEYINPUT102), .B1(new_n653), .B2(new_n654), .ZN(new_n656));
  OAI221_X1 g455(.A(new_n651), .B1(new_n652), .B2(new_n649), .C1(new_n655), .C2(new_n656), .ZN(G1325gat));
  AOI21_X1  g456(.A(G15gat), .B1(new_n646), .B2(new_n322), .ZN(new_n658));
  XOR2_X1   g457(.A(new_n658), .B(KEYINPUT103), .Z(new_n659));
  NAND2_X1  g458(.A1(new_n518), .A2(new_n519), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  AND2_X1   g460(.A1(new_n661), .A2(G15gat), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n659), .B1(new_n646), .B2(new_n662), .ZN(G1326gat));
  NAND2_X1  g462(.A1(new_n646), .A2(new_n474), .ZN(new_n664));
  XNOR2_X1  g463(.A(KEYINPUT43), .B(G22gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(G1327gat));
  NOR2_X1   g465(.A1(new_n521), .A2(new_n569), .ZN(new_n667));
  INV_X1    g466(.A(new_n644), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n668), .A2(new_n588), .A3(new_n618), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(G29gat), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n670), .A2(new_n671), .A3(new_n477), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT45), .ZN(new_n673));
  INV_X1    g472(.A(new_n569), .ZN(new_n674));
  INV_X1    g473(.A(new_n588), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n674), .A2(new_n675), .A3(new_n644), .ZN(new_n676));
  INV_X1    g475(.A(new_n418), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n475), .B1(new_n677), .B2(new_n421), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n494), .B1(new_n678), .B2(new_n491), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n495), .A2(new_n503), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n516), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT104), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n682), .B1(new_n426), .B2(new_n463), .ZN(new_n683));
  OAI211_X1 g482(.A(KEYINPUT104), .B(new_n474), .C1(new_n477), .C2(new_n366), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n681), .A2(new_n683), .A3(new_n660), .A4(new_n684), .ZN(new_n685));
  NOR4_X1   g484(.A1(new_n312), .A2(new_n321), .A3(new_n474), .A4(new_n471), .ZN(new_n686));
  AOI22_X1  g485(.A1(new_n686), .A2(new_n426), .B1(new_n471), .B2(new_n470), .ZN(new_n687));
  AND3_X1   g486(.A1(new_n685), .A2(KEYINPUT105), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(KEYINPUT105), .B1(new_n685), .B2(new_n687), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n618), .A2(KEYINPUT44), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  OR3_X1    g490(.A1(new_n688), .A2(new_n689), .A3(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n520), .A2(new_n478), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(new_n687), .ZN(new_n695));
  INV_X1    g494(.A(new_n618), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n693), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n676), .B1(new_n692), .B2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n477), .ZN(new_n701));
  OAI21_X1  g500(.A(G29gat), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n673), .A2(new_n702), .ZN(G1328gat));
  INV_X1    g502(.A(G36gat), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n670), .A2(new_n704), .A3(new_n465), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT106), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT46), .ZN(new_n707));
  OR2_X1    g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n706), .A2(new_n707), .ZN(new_n709));
  INV_X1    g508(.A(new_n465), .ZN(new_n710));
  OAI21_X1  g509(.A(G36gat), .B1(new_n700), .B2(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n708), .A2(new_n709), .A3(new_n711), .ZN(G1329gat));
  XOR2_X1   g511(.A(KEYINPUT107), .B(KEYINPUT47), .Z(new_n713));
  INV_X1    g512(.A(G43gat), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n714), .B1(new_n699), .B2(new_n661), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT108), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n667), .A2(new_n714), .A3(new_n322), .A4(new_n669), .ZN(new_n718));
  XOR2_X1   g517(.A(new_n718), .B(KEYINPUT109), .Z(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(new_n715), .B2(new_n716), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n713), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n718), .A2(KEYINPUT47), .ZN(new_n722));
  OR2_X1    g521(.A1(new_n715), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n721), .A2(new_n723), .ZN(G1330gat));
  INV_X1    g523(.A(KEYINPUT110), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n699), .A2(new_n474), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n725), .B1(new_n726), .B2(new_n453), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n670), .A2(new_n453), .A3(new_n474), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n728), .B1(new_n726), .B2(new_n453), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT48), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n727), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  OAI221_X1 g530(.A(new_n728), .B1(new_n725), .B2(KEYINPUT48), .C1(new_n726), .C2(new_n453), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(G1331gat));
  NOR2_X1   g532(.A1(new_n688), .A2(new_n689), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n674), .A2(new_n619), .A3(new_n644), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n477), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g538(.A(new_n710), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(KEYINPUT111), .ZN(new_n742));
  NOR2_X1   g541(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n742), .B(new_n743), .ZN(G1333gat));
  INV_X1    g543(.A(G71gat), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n737), .A2(new_n745), .A3(new_n322), .ZN(new_n746));
  OAI21_X1  g545(.A(G71gat), .B1(new_n736), .B2(new_n660), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(KEYINPUT112), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT112), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n746), .A2(new_n750), .A3(new_n747), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT50), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n749), .A2(KEYINPUT50), .A3(new_n751), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(G1334gat));
  NAND2_X1  g555(.A1(new_n737), .A2(new_n474), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g557(.A1(new_n685), .A2(new_n687), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(new_n696), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT113), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n674), .A2(new_n588), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n618), .B1(new_n685), .B2(new_n687), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(KEYINPUT113), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n762), .A2(new_n763), .A3(new_n765), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n644), .B1(new_n766), .B2(KEYINPUT51), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT51), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n762), .A2(new_n768), .A3(new_n763), .A4(new_n765), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n701), .A2(new_n600), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n763), .A2(new_n668), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n688), .A2(new_n689), .A3(new_n691), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n774), .B1(new_n775), .B2(new_n697), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n600), .B1(new_n776), .B2(new_n701), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n772), .A2(new_n777), .ZN(G1336gat));
  OAI211_X1 g577(.A(new_n465), .B(new_n774), .C1(new_n775), .C2(new_n697), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(G92gat), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n764), .A2(KEYINPUT113), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n763), .B1(new_n764), .B2(KEYINPUT113), .ZN(new_n782));
  OAI21_X1  g581(.A(KEYINPUT51), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n710), .A2(G92gat), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n783), .A2(new_n769), .A3(new_n668), .A4(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n780), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT115), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n785), .A2(KEYINPUT114), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(new_n780), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n785), .A2(KEYINPUT114), .ZN(new_n792));
  OAI21_X1  g591(.A(KEYINPUT52), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n789), .A2(new_n793), .ZN(G1337gat));
  NOR3_X1   g593(.A1(new_n776), .A2(new_n597), .A3(new_n660), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n770), .A2(new_n322), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n795), .B1(new_n796), .B2(new_n597), .ZN(G1338gat));
  NOR2_X1   g596(.A1(new_n463), .A2(G106gat), .ZN(new_n798));
  AND4_X1   g597(.A1(new_n668), .A2(new_n783), .A3(new_n769), .A4(new_n798), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n474), .B(new_n774), .C1(new_n775), .C2(new_n697), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(G106gat), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(KEYINPUT118), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT117), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n799), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n767), .A2(new_n803), .A3(new_n769), .A4(new_n798), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT116), .ZN(new_n806));
  AND3_X1   g605(.A1(new_n800), .A2(new_n806), .A3(G106gat), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n806), .B1(new_n800), .B2(G106gat), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n805), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(KEYINPUT53), .B1(new_n804), .B2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(new_n799), .ZN(new_n811));
  NOR2_X1   g610(.A1(KEYINPUT118), .A2(KEYINPUT53), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n811), .A2(new_n801), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n810), .A2(new_n813), .ZN(G1339gat));
  NAND2_X1  g613(.A1(new_n322), .A2(new_n463), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n564), .A2(new_n566), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n543), .A2(new_n545), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n549), .A2(new_n542), .ZN(new_n818));
  OAI22_X1  g617(.A1(new_n817), .A2(KEYINPUT119), .B1(new_n818), .B2(new_n544), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n817), .A2(KEYINPUT119), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n555), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n816), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n630), .A2(new_n631), .A3(new_n628), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n633), .A2(KEYINPUT54), .A3(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n637), .B1(new_n632), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT55), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n824), .A2(KEYINPUT55), .A3(new_n826), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n829), .A2(new_n638), .A3(new_n830), .ZN(new_n831));
  OAI22_X1  g630(.A1(new_n644), .A2(new_n822), .B1(new_n831), .B2(new_n569), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n832), .A2(new_n618), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n696), .A2(new_n638), .A3(new_n830), .A4(new_n829), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n834), .A2(new_n822), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n675), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n620), .A2(new_n569), .A3(new_n644), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n815), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n701), .A2(new_n465), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n674), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(G113gat), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n842), .B1(new_n259), .B2(new_n841), .ZN(G1340gat));
  NAND2_X1  g642(.A1(new_n840), .A2(new_n668), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n844), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g644(.A1(new_n840), .A2(new_n588), .ZN(new_n846));
  XNOR2_X1  g645(.A(new_n846), .B(G127gat), .ZN(G1342gat));
  INV_X1    g646(.A(KEYINPUT120), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n840), .A2(new_n696), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n848), .B1(new_n849), .B2(G134gat), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n840), .A2(KEYINPUT120), .A3(new_n263), .A4(new_n696), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  OR2_X1    g651(.A1(new_n852), .A2(KEYINPUT56), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(KEYINPUT56), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n849), .A2(G134gat), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(G1343gat));
  AOI21_X1  g655(.A(new_n463), .B1(new_n836), .B2(new_n837), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n660), .ZN(new_n858));
  OR3_X1    g657(.A1(new_n858), .A2(KEYINPUT121), .A3(new_n701), .ZN(new_n859));
  OAI21_X1  g658(.A(KEYINPUT121), .B1(new_n858), .B2(new_n701), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n859), .A2(new_n710), .A3(new_n860), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n861), .A2(G141gat), .A3(new_n569), .ZN(new_n862));
  XNOR2_X1  g661(.A(new_n857), .B(KEYINPUT57), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n660), .A2(new_n839), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n863), .A2(new_n674), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(G141gat), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT58), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(new_n858), .ZN(new_n869));
  NOR4_X1   g668(.A1(new_n701), .A2(new_n569), .A3(G141gat), .A4(new_n465), .ZN(new_n870));
  AOI22_X1  g669(.A1(new_n865), .A2(G141gat), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI22_X1  g670(.A1(new_n862), .A2(new_n868), .B1(new_n867), .B2(new_n871), .ZN(G1344gat));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n863), .A2(new_n864), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n873), .B(G148gat), .C1(new_n874), .C2(new_n644), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n835), .B1(new_n832), .B2(new_n618), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n675), .B1(new_n876), .B2(KEYINPUT122), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT122), .ZN(new_n878));
  AOI211_X1 g677(.A(new_n878), .B(new_n835), .C1(new_n618), .C2(new_n832), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n837), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(KEYINPUT57), .B1(new_n880), .B2(new_n474), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT57), .ZN(new_n882));
  AOI211_X1 g681(.A(new_n882), .B(new_n463), .C1(new_n836), .C2(new_n837), .ZN(new_n883));
  OAI211_X1 g682(.A(new_n668), .B(new_n864), .C1(new_n881), .C2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(G148gat), .ZN(new_n885));
  AOI21_X1  g684(.A(KEYINPUT123), .B1(new_n885), .B2(KEYINPUT59), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT123), .ZN(new_n887));
  AOI211_X1 g686(.A(new_n887), .B(new_n873), .C1(new_n884), .C2(G148gat), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n875), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  OR2_X1    g688(.A1(new_n644), .A2(G148gat), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n889), .B1(new_n861), .B2(new_n890), .ZN(G1345gat));
  OAI21_X1  g690(.A(G155gat), .B1(new_n874), .B2(new_n675), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n588), .A2(new_n375), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n892), .B1(new_n861), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(KEYINPUT124), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT124), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n892), .B(new_n896), .C1(new_n861), .C2(new_n893), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n895), .A2(new_n897), .ZN(G1346gat));
  OAI21_X1  g697(.A(G162gat), .B1(new_n874), .B2(new_n618), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n696), .A2(new_n376), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n899), .B1(new_n861), .B2(new_n900), .ZN(G1347gat));
  NOR2_X1   g700(.A1(new_n477), .A2(new_n710), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n838), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n903), .A2(new_n569), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n904), .B(new_n206), .ZN(G1348gat));
  NOR2_X1   g704(.A1(new_n903), .A2(new_n644), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(new_n207), .ZN(G1349gat));
  INV_X1    g706(.A(KEYINPUT125), .ZN(new_n908));
  INV_X1    g707(.A(new_n903), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(new_n588), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n908), .B1(new_n910), .B2(new_n219), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n909), .A2(KEYINPUT125), .A3(new_n330), .A4(new_n588), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n910), .A2(G183gat), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT60), .ZN(G1350gat));
  NOR2_X1   g714(.A1(new_n903), .A2(new_n618), .ZN(new_n916));
  NAND2_X1  g715(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  XOR2_X1   g717(.A(KEYINPUT61), .B(G190gat), .Z(new_n919));
  OAI21_X1  g718(.A(new_n918), .B1(new_n916), .B2(new_n919), .ZN(G1351gat));
  NOR3_X1   g719(.A1(new_n858), .A2(new_n477), .A3(new_n710), .ZN(new_n921));
  AOI21_X1  g720(.A(G197gat), .B1(new_n921), .B2(new_n674), .ZN(new_n922));
  OR2_X1    g721(.A1(new_n881), .A2(new_n883), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n660), .A2(new_n902), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n674), .A2(G197gat), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n922), .B1(new_n926), .B2(new_n927), .ZN(G1352gat));
  NAND3_X1  g727(.A1(new_n921), .A2(new_n636), .A3(new_n668), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n929), .B1(KEYINPUT126), .B2(KEYINPUT62), .ZN(new_n930));
  XNOR2_X1  g729(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n930), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n923), .A2(new_n668), .A3(new_n925), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(G204gat), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n934), .ZN(G1353gat));
  OAI211_X1 g734(.A(new_n588), .B(new_n925), .C1(new_n881), .C2(new_n883), .ZN(new_n936));
  AND3_X1   g735(.A1(new_n936), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n937));
  AOI21_X1  g736(.A(KEYINPUT63), .B1(new_n936), .B2(G211gat), .ZN(new_n938));
  INV_X1    g737(.A(new_n921), .ZN(new_n939));
  OR2_X1    g738(.A1(new_n675), .A2(G211gat), .ZN(new_n940));
  OAI22_X1  g739(.A1(new_n937), .A2(new_n938), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT127), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI221_X1 g742(.A(KEYINPUT127), .B1(new_n939), .B2(new_n940), .C1(new_n937), .C2(new_n938), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(G1354gat));
  AOI21_X1  g744(.A(G218gat), .B1(new_n921), .B2(new_n696), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n696), .A2(G218gat), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n946), .B1(new_n926), .B2(new_n947), .ZN(G1355gat));
endmodule


