//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 1 0 0 0 1 0 1 0 1 1 1 0 0 0 1 1 1 0 0 1 0 1 1 0 0 0 0 1 1 1 0 1 0 1 1 1 1 1 1 0 0 0 0 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:31 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n734, new_n735, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT72), .ZN(new_n188));
  INV_X1    g002(.A(G140), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G125), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n188), .B1(new_n190), .B2(KEYINPUT16), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT16), .ZN(new_n192));
  NAND4_X1  g006(.A1(new_n192), .A2(new_n189), .A3(KEYINPUT72), .A4(G125), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G125), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G140), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n190), .A2(new_n196), .A3(KEYINPUT16), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(KEYINPUT71), .ZN(new_n198));
  XNOR2_X1  g012(.A(G125), .B(G140), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT71), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(new_n200), .A3(KEYINPUT16), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n194), .A2(new_n198), .A3(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G146), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n194), .A2(new_n198), .A3(new_n201), .A4(G146), .ZN(new_n205));
  INV_X1    g019(.A(G131), .ZN(new_n206));
  NOR2_X1   g020(.A1(G237), .A2(G953), .ZN(new_n207));
  AND2_X1   g021(.A1(KEYINPUT86), .A2(G143), .ZN(new_n208));
  NOR2_X1   g022(.A1(KEYINPUT86), .A2(G143), .ZN(new_n209));
  OAI211_X1 g023(.A(G214), .B(new_n207), .C1(new_n208), .C2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n207), .A2(G214), .ZN(new_n211));
  NAND2_X1  g025(.A1(KEYINPUT86), .A2(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n206), .B1(new_n210), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT17), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n204), .A2(new_n205), .A3(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT89), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n204), .A2(KEYINPUT89), .A3(new_n205), .A4(new_n215), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT17), .ZN(new_n220));
  AND3_X1   g034(.A1(new_n210), .A2(new_n213), .A3(new_n206), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT88), .ZN(new_n222));
  NOR3_X1   g036(.A1(new_n221), .A2(new_n214), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n210), .A2(new_n213), .ZN(new_n224));
  NOR3_X1   g038(.A1(new_n224), .A2(KEYINPUT88), .A3(G131), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n220), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n218), .A2(new_n219), .A3(new_n226), .ZN(new_n227));
  XNOR2_X1  g041(.A(G113), .B(G122), .ZN(new_n228));
  INV_X1    g042(.A(G104), .ZN(new_n229));
  XNOR2_X1  g043(.A(new_n228), .B(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n224), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT18), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n231), .B1(new_n232), .B2(new_n206), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT87), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n234), .B1(new_n199), .B2(new_n203), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n235), .B1(new_n203), .B2(new_n199), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n224), .A2(KEYINPUT18), .A3(G131), .ZN(new_n237));
  OR3_X1    g051(.A1(new_n199), .A2(KEYINPUT87), .A3(new_n203), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n233), .A2(new_n236), .A3(new_n237), .A4(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n227), .A2(new_n230), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n230), .B1(new_n227), .B2(new_n239), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n187), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(KEYINPUT91), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT91), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n245), .B(new_n187), .C1(new_n241), .C2(new_n242), .ZN(new_n246));
  XOR2_X1   g060(.A(KEYINPUT90), .B(G475), .Z(new_n247));
  NAND3_X1  g061(.A1(new_n244), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G134), .ZN(new_n249));
  INV_X1    g063(.A(G128), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n250), .A2(G143), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(G143), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n251), .B1(KEYINPUT13), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT92), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n249), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G143), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G128), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT13), .ZN(new_n258));
  OAI21_X1  g072(.A(KEYINPUT92), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n255), .B1(new_n253), .B2(new_n259), .ZN(new_n260));
  XNOR2_X1  g074(.A(G116), .B(G122), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G107), .ZN(new_n263));
  INV_X1    g077(.A(G107), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  AND2_X1   g079(.A1(new_n257), .A2(new_n252), .ZN(new_n266));
  AOI22_X1  g080(.A1(new_n263), .A2(new_n265), .B1(new_n249), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n260), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n266), .B(new_n249), .ZN(new_n269));
  INV_X1    g083(.A(G116), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n270), .A2(KEYINPUT14), .A3(G122), .ZN(new_n271));
  OAI211_X1 g085(.A(G107), .B(new_n271), .C1(new_n262), .C2(KEYINPUT14), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n269), .A2(new_n265), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n268), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g088(.A(KEYINPUT9), .B(G234), .ZN(new_n275));
  INV_X1    g089(.A(G217), .ZN(new_n276));
  NOR3_X1   g090(.A1(new_n275), .A2(new_n276), .A3(G953), .ZN(new_n277));
  XOR2_X1   g091(.A(new_n277), .B(KEYINPUT93), .Z(new_n278));
  OR2_X1    g092(.A1(new_n274), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n274), .A2(new_n278), .ZN(new_n280));
  AOI21_X1  g094(.A(G902), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G478), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n282), .A2(KEYINPUT15), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n281), .B(new_n283), .ZN(new_n284));
  OR3_X1    g098(.A1(new_n221), .A2(new_n214), .A3(new_n222), .ZN(new_n285));
  INV_X1    g099(.A(new_n225), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n199), .B(KEYINPUT19), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n203), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n285), .A2(new_n205), .A3(new_n286), .A4(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(new_n239), .ZN(new_n290));
  INV_X1    g104(.A(new_n230), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n240), .A2(new_n292), .ZN(new_n293));
  NOR2_X1   g107(.A1(G475), .A2(G902), .ZN(new_n294));
  AOI21_X1  g108(.A(KEYINPUT20), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT20), .ZN(new_n296));
  INV_X1    g110(.A(new_n294), .ZN(new_n297));
  AOI211_X1 g111(.A(new_n296), .B(new_n297), .C1(new_n240), .C2(new_n292), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n248), .A2(new_n284), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n203), .A2(G143), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n256), .A2(G146), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(KEYINPUT1), .B1(new_n256), .B2(G146), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT65), .ZN(new_n305));
  OAI21_X1  g119(.A(G128), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(KEYINPUT65), .B1(new_n301), .B2(KEYINPUT1), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n303), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n250), .A2(KEYINPUT1), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n309), .A2(new_n301), .A3(new_n302), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n308), .A2(new_n195), .A3(new_n311), .ZN(new_n312));
  AND2_X1   g126(.A1(KEYINPUT0), .A2(G128), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n301), .A2(new_n302), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT64), .ZN(new_n315));
  XNOR2_X1  g129(.A(G143), .B(G146), .ZN(new_n316));
  XNOR2_X1  g130(.A(KEYINPUT0), .B(G128), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n314), .B(new_n315), .C1(new_n316), .C2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n313), .ZN(new_n319));
  OR2_X1    g133(.A1(KEYINPUT0), .A2(G128), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n303), .A2(KEYINPUT64), .A3(new_n319), .A4(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n318), .A2(G125), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n312), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT7), .ZN(new_n324));
  INV_X1    g138(.A(G224), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n325), .A2(G953), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n323), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(KEYINPUT3), .B1(new_n229), .B2(G107), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT3), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(new_n264), .A3(G104), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n229), .A2(G107), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n328), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G101), .ZN(new_n333));
  AOI21_X1  g147(.A(G101), .B1(new_n229), .B2(G107), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n328), .A2(new_n334), .A3(new_n330), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n333), .A2(KEYINPUT4), .A3(new_n335), .ZN(new_n336));
  XOR2_X1   g150(.A(KEYINPUT75), .B(KEYINPUT4), .Z(new_n337));
  NAND3_X1  g151(.A1(new_n332), .A2(G101), .A3(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT67), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n339), .B1(new_n270), .B2(G119), .ZN(new_n340));
  INV_X1    g154(.A(G119), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n341), .A2(KEYINPUT67), .A3(G116), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n270), .A2(G119), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n340), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(KEYINPUT2), .B(G113), .ZN(new_n345));
  AND3_X1   g159(.A1(new_n344), .A2(KEYINPUT66), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n345), .B1(new_n344), .B2(KEYINPUT66), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n336), .B(new_n338), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  AND3_X1   g162(.A1(new_n340), .A2(new_n342), .A3(new_n343), .ZN(new_n349));
  INV_X1    g163(.A(new_n345), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n340), .A2(new_n342), .A3(KEYINPUT5), .A4(new_n343), .ZN(new_n351));
  NOR3_X1   g165(.A1(new_n270), .A2(KEYINPUT5), .A3(G119), .ZN(new_n352));
  INV_X1    g166(.A(G113), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AOI22_X1  g168(.A1(new_n349), .A2(new_n350), .B1(new_n351), .B2(new_n354), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n229), .A2(G107), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n264), .A2(G104), .ZN(new_n357));
  OAI21_X1  g171(.A(G101), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT76), .ZN(new_n359));
  AND3_X1   g173(.A1(new_n358), .A2(new_n335), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n359), .B1(new_n358), .B2(new_n335), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n355), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  XNOR2_X1  g176(.A(G110), .B(G122), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n348), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n326), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n312), .A2(KEYINPUT7), .A3(new_n365), .A4(new_n322), .ZN(new_n366));
  AND3_X1   g180(.A1(new_n327), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n363), .B(KEYINPUT8), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n358), .A2(new_n335), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(KEYINPUT83), .B1(new_n355), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n362), .ZN(new_n372));
  NOR3_X1   g186(.A1(new_n355), .A2(new_n370), .A3(KEYINPUT83), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n368), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(G902), .B1(new_n367), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n348), .A2(new_n362), .ZN(new_n376));
  INV_X1    g190(.A(new_n363), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n378), .A2(KEYINPUT6), .A3(new_n364), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n323), .B(new_n326), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT6), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n376), .A2(new_n381), .A3(new_n377), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n379), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n375), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(G210), .B1(G237), .B2(G902), .ZN(new_n385));
  XOR2_X1   g199(.A(new_n385), .B(KEYINPUT84), .Z(new_n386));
  NAND2_X1  g200(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n386), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n375), .A2(new_n383), .A3(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT85), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n387), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  OR2_X1    g205(.A1(new_n389), .A2(new_n390), .ZN(new_n392));
  NAND2_X1  g206(.A1(G234), .A2(G237), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(G902), .A3(G953), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(KEYINPUT21), .B(G898), .ZN(new_n396));
  INV_X1    g210(.A(G953), .ZN(new_n397));
  AND2_X1   g211(.A1(new_n397), .A2(G952), .ZN(new_n398));
  AOI22_X1  g212(.A1(new_n395), .A2(new_n396), .B1(new_n393), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(G214), .B1(G237), .B2(G902), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n391), .A2(new_n392), .A3(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n300), .A2(new_n403), .ZN(new_n404));
  XOR2_X1   g218(.A(KEYINPUT68), .B(KEYINPUT27), .Z(new_n405));
  NAND2_X1  g219(.A1(new_n207), .A2(G210), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n405), .B(new_n406), .ZN(new_n407));
  XNOR2_X1  g221(.A(KEYINPUT26), .B(G101), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n407), .B(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT28), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n346), .A2(new_n347), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT11), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n414), .B1(new_n249), .B2(G137), .ZN(new_n415));
  INV_X1    g229(.A(G137), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n416), .A2(KEYINPUT11), .A3(G134), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n249), .A2(G137), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n415), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G131), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n415), .A2(new_n417), .A3(new_n206), .A4(new_n418), .ZN(new_n421));
  AOI22_X1  g235(.A1(new_n318), .A2(new_n321), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n249), .A2(G137), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n416), .A2(G134), .ZN(new_n424));
  OAI21_X1  g238(.A(G131), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n421), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n426), .B1(new_n308), .B2(new_n311), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n413), .B1(new_n422), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT1), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n429), .B1(G143), .B2(new_n203), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n250), .B1(new_n430), .B2(KEYINPUT65), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n304), .A2(new_n305), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n316), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n421), .B(new_n425), .C1(new_n433), .C2(new_n310), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n318), .A2(new_n321), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n420), .A2(new_n421), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n434), .A2(new_n412), .A3(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n411), .B1(new_n428), .B2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n438), .A2(new_n411), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n410), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT30), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n434), .A2(new_n443), .A3(new_n437), .ZN(new_n444));
  OAI21_X1  g258(.A(KEYINPUT30), .B1(new_n427), .B2(new_n422), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n413), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n447), .A2(new_n438), .A3(new_n410), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT31), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n438), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n451), .B1(new_n446), .B2(new_n413), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n452), .A2(KEYINPUT31), .A3(new_n410), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n442), .B1(new_n450), .B2(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(G472), .A2(G902), .ZN(new_n455));
  XOR2_X1   g269(.A(new_n455), .B(KEYINPUT69), .Z(new_n456));
  OAI21_X1  g270(.A(KEYINPUT32), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n441), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n409), .B1(new_n458), .B2(new_n439), .ZN(new_n459));
  AOI21_X1  g273(.A(KEYINPUT31), .B1(new_n452), .B2(new_n410), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n412), .B1(new_n444), .B2(new_n445), .ZN(new_n461));
  NOR4_X1   g275(.A1(new_n461), .A2(new_n451), .A3(new_n449), .A4(new_n409), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n459), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT32), .ZN(new_n464));
  INV_X1    g278(.A(new_n456), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n457), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n440), .A2(new_n441), .A3(new_n410), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT29), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n468), .B(new_n469), .C1(new_n410), .C2(new_n452), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT70), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n458), .B1(new_n439), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n440), .A2(KEYINPUT70), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n472), .A2(new_n473), .A3(KEYINPUT29), .A4(new_n410), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n470), .A2(new_n187), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(G472), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n467), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n276), .B1(G234), .B2(new_n187), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT25), .ZN(new_n480));
  XNOR2_X1  g294(.A(KEYINPUT22), .B(G137), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n397), .A2(G221), .A3(G234), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n481), .B(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n204), .A2(new_n205), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n250), .A2(G119), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT23), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n341), .A2(G128), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n250), .A2(KEYINPUT23), .A3(G119), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(G110), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n489), .A2(new_n486), .ZN(new_n493));
  XNOR2_X1  g307(.A(KEYINPUT24), .B(G110), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n485), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(G110), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n488), .A2(new_n490), .A3(new_n498), .A4(new_n489), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n493), .A2(new_n494), .ZN(new_n500));
  AOI22_X1  g314(.A1(new_n499), .A2(new_n500), .B1(new_n203), .B2(new_n199), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n205), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n484), .B1(new_n497), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n497), .A2(KEYINPUT73), .A3(new_n502), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT73), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n495), .B1(new_n204), .B2(new_n205), .ZN(new_n506));
  INV_X1    g320(.A(new_n502), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n503), .B1(new_n509), .B2(new_n484), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n480), .B1(new_n510), .B2(G902), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n483), .B1(new_n504), .B2(new_n508), .ZN(new_n512));
  OAI211_X1 g326(.A(KEYINPUT25), .B(new_n187), .C1(new_n512), .C2(new_n503), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n479), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(KEYINPUT73), .B1(new_n497), .B2(new_n502), .ZN(new_n515));
  NOR3_X1   g329(.A1(new_n506), .A2(new_n507), .A3(new_n505), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n484), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n503), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n478), .A2(G902), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n514), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n404), .A2(new_n477), .A3(new_n521), .ZN(new_n522));
  XNOR2_X1  g336(.A(G110), .B(G140), .ZN(new_n523));
  INV_X1    g337(.A(G227), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n524), .A2(G953), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n523), .B(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n369), .A2(KEYINPUT76), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n358), .A2(new_n335), .A3(new_n359), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n527), .A2(new_n528), .A3(new_n311), .A4(new_n308), .ZN(new_n529));
  AOI22_X1  g343(.A1(new_n304), .A2(G128), .B1(new_n301), .B2(new_n302), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n530), .A2(new_n310), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n531), .A2(new_n369), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n436), .A2(KEYINPUT12), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(KEYINPUT77), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT77), .ZN(new_n538));
  AOI211_X1 g352(.A(new_n538), .B(new_n535), .C1(new_n529), .C2(new_n533), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n360), .A2(new_n361), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n433), .A2(new_n310), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n532), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n436), .B1(new_n543), .B2(KEYINPUT78), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT78), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n534), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n540), .B1(new_n547), .B2(KEYINPUT12), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n308), .A2(new_n311), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n549), .B(KEYINPUT10), .C1(new_n361), .C2(new_n360), .ZN(new_n550));
  INV_X1    g364(.A(new_n436), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT10), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n552), .B1(new_n531), .B2(new_n369), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n336), .A2(new_n435), .A3(new_n338), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n550), .A2(new_n551), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(KEYINPUT79), .B1(new_n548), .B2(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n551), .B1(new_n534), .B2(new_n545), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n543), .A2(KEYINPUT78), .ZN(new_n558));
  AOI21_X1  g372(.A(KEYINPUT12), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n538), .B1(new_n543), .B2(new_n535), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n534), .A2(KEYINPUT77), .A3(new_n536), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  OAI211_X1 g376(.A(KEYINPUT79), .B(new_n555), .C1(new_n559), .C2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n526), .B1(new_n556), .B2(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(KEYINPUT10), .B1(new_n433), .B2(new_n310), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n554), .B(new_n553), .C1(new_n566), .C2(new_n541), .ZN(new_n567));
  AND3_X1   g381(.A1(new_n567), .A2(KEYINPUT80), .A3(new_n436), .ZN(new_n568));
  AOI21_X1  g382(.A(KEYINPUT80), .B1(new_n567), .B2(new_n436), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n526), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n555), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n565), .A2(G469), .A3(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT82), .ZN(new_n576));
  INV_X1    g390(.A(new_n555), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n567), .A2(new_n436), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT80), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n567), .A2(KEYINPUT80), .A3(new_n436), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n577), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n576), .B1(new_n582), .B2(new_n571), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n555), .B1(new_n568), .B2(new_n569), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n584), .A2(KEYINPUT82), .A3(new_n526), .ZN(new_n585));
  AND3_X1   g399(.A1(new_n555), .A2(KEYINPUT81), .A3(new_n571), .ZN(new_n586));
  AOI21_X1  g400(.A(KEYINPUT81), .B1(new_n555), .B2(new_n571), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n548), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n583), .A2(new_n585), .A3(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(G469), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n590), .A2(new_n591), .A3(new_n187), .ZN(new_n592));
  NAND2_X1  g406(.A1(G469), .A2(G902), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n575), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(G221), .B1(new_n275), .B2(G902), .ZN(new_n595));
  XOR2_X1   g409(.A(new_n595), .B(KEYINPUT74), .Z(new_n596));
  NAND2_X1  g410(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n522), .A2(new_n597), .ZN(new_n598));
  XOR2_X1   g412(.A(new_n598), .B(G101), .Z(G3));
  OAI21_X1  g413(.A(G472), .B1(new_n454), .B2(G902), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n463), .A2(new_n465), .ZN(new_n601));
  AND2_X1   g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n594), .A2(new_n596), .A3(new_n521), .A4(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n227), .A2(new_n239), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(new_n291), .ZN(new_n606));
  AOI21_X1  g420(.A(G902), .B1(new_n606), .B2(new_n240), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n247), .B1(new_n607), .B2(new_n245), .ZN(new_n608));
  INV_X1    g422(.A(new_n246), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n299), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n401), .B1(new_n387), .B2(new_n389), .ZN(new_n612));
  INV_X1    g426(.A(new_n399), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AND4_X1   g428(.A1(KEYINPUT94), .A2(new_n279), .A3(KEYINPUT33), .A4(new_n280), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT94), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n280), .A2(new_n616), .ZN(new_n617));
  AOI22_X1  g431(.A1(new_n617), .A2(KEYINPUT33), .B1(new_n279), .B2(new_n280), .ZN(new_n618));
  OAI21_X1  g432(.A(G478), .B1(new_n615), .B2(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n282), .A2(new_n187), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n620), .B1(new_n281), .B2(new_n282), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NOR3_X1   g436(.A1(new_n611), .A2(new_n614), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n604), .A2(new_n623), .ZN(new_n624));
  XOR2_X1   g438(.A(KEYINPUT34), .B(G104), .Z(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G6));
  NOR2_X1   g440(.A1(new_n610), .A2(new_n284), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n628), .A2(new_n614), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n604), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT35), .B(G107), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G9));
  NAND3_X1  g446(.A1(new_n594), .A2(new_n596), .A3(new_n602), .ZN(new_n633));
  AOI21_X1  g447(.A(KEYINPUT25), .B1(new_n519), .B2(new_n187), .ZN(new_n634));
  INV_X1    g448(.A(new_n513), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n478), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n484), .A2(KEYINPUT36), .ZN(new_n637));
  AND2_X1   g451(.A1(new_n509), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n509), .A2(new_n637), .ZN(new_n639));
  NOR4_X1   g453(.A1(new_n638), .A2(new_n639), .A3(G902), .A4(new_n478), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n636), .A2(new_n641), .A3(KEYINPUT95), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT95), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n643), .B1(new_n514), .B2(new_n640), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n404), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n633), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT37), .B(G110), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G12));
  NAND3_X1  g463(.A1(new_n645), .A2(new_n477), .A3(new_n612), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n650), .A2(new_n597), .ZN(new_n651));
  INV_X1    g465(.A(G900), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n395), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n398), .A2(new_n393), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n628), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n651), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G128), .ZN(G30));
  INV_X1    g473(.A(new_n597), .ZN(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT97), .B(KEYINPUT39), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n655), .B(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(KEYINPUT40), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n391), .A2(new_n392), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(KEYINPUT38), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n452), .A2(new_n409), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n428), .A2(new_n438), .A3(new_n409), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n187), .ZN(new_n669));
  OAI21_X1  g483(.A(G472), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n454), .A2(KEYINPUT32), .A3(new_n456), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n464), .B1(new_n463), .B2(new_n465), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n670), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT96), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n467), .A2(KEYINPUT96), .A3(new_n670), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n284), .A2(new_n401), .ZN(new_n678));
  AND4_X1   g492(.A1(new_n610), .A2(new_n642), .A3(new_n644), .A4(new_n678), .ZN(new_n679));
  AND3_X1   g493(.A1(new_n666), .A2(new_n677), .A3(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT40), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n660), .A2(new_n681), .A3(new_n662), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n664), .A2(new_n680), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(KEYINPUT98), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(new_n256), .ZN(G45));
  AOI211_X1 g499(.A(new_n656), .B(new_n622), .C1(new_n248), .C2(new_n299), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n651), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G146), .ZN(G48));
  INV_X1    g502(.A(new_n595), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT100), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n584), .A2(new_n526), .ZN(new_n691));
  AOI22_X1  g505(.A1(new_n691), .A2(new_n576), .B1(new_n548), .B2(new_n588), .ZN(new_n692));
  AOI21_X1  g506(.A(G902), .B1(new_n692), .B2(new_n585), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n690), .B1(new_n693), .B2(new_n591), .ZN(new_n694));
  OAI21_X1  g508(.A(G469), .B1(new_n693), .B2(KEYINPUT99), .ZN(new_n695));
  AND3_X1   g509(.A1(new_n590), .A2(KEYINPUT99), .A3(new_n187), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n694), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n590), .A2(new_n187), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT99), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n590), .A2(KEYINPUT99), .A3(new_n187), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n700), .A2(new_n690), .A3(G469), .A4(new_n701), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n689), .B1(new_n697), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n477), .A2(new_n521), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  AND2_X1   g519(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n623), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT41), .B(G113), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G15));
  NAND2_X1  g523(.A1(new_n706), .A2(new_n629), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G116), .ZN(G18));
  AND4_X1   g525(.A1(new_n477), .A2(new_n645), .A3(new_n284), .A4(new_n611), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n703), .A2(new_n613), .A3(new_n612), .A4(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G119), .ZN(G21));
  NOR2_X1   g528(.A1(new_n460), .A2(new_n462), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n410), .B1(new_n472), .B2(new_n473), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n465), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AND2_X1   g531(.A1(new_n600), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n718), .A2(new_n521), .A3(new_n613), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n387), .A2(new_n389), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n610), .A2(new_n720), .A3(new_n678), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(KEYINPUT101), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT101), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n610), .A2(new_n723), .A3(new_n720), .A4(new_n678), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n719), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  AOI21_X1  g539(.A(KEYINPUT99), .B1(new_n590), .B2(new_n187), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n696), .A2(new_n726), .A3(new_n591), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n592), .A2(KEYINPUT100), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n702), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  AND4_X1   g543(.A1(KEYINPUT102), .A2(new_n725), .A3(new_n595), .A4(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(KEYINPUT102), .B1(new_n703), .B2(new_n725), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  XOR2_X1   g546(.A(new_n732), .B(G122), .Z(G24));
  AND3_X1   g547(.A1(new_n686), .A2(new_n645), .A3(new_n718), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n729), .A2(new_n734), .A3(new_n595), .A4(new_n612), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G125), .ZN(G27));
  INV_X1    g550(.A(KEYINPUT104), .ZN(new_n737));
  AOI211_X1 g551(.A(new_n689), .B(new_n401), .C1(new_n391), .C2(new_n392), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT103), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n565), .A2(new_n739), .A3(G469), .A4(new_n574), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n740), .A2(new_n592), .A3(new_n593), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n555), .B1(new_n559), .B2(new_n562), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT79), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n563), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n573), .B1(new_n745), .B2(new_n526), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n739), .B1(new_n746), .B2(G469), .ZN(new_n747));
  OAI211_X1 g561(.A(new_n737), .B(new_n738), .C1(new_n741), .C2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n592), .A2(new_n593), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n575), .A2(KEYINPUT103), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n750), .A2(new_n751), .A3(new_n740), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n737), .B1(new_n752), .B2(new_n738), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n705), .B(new_n686), .C1(new_n749), .C2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT42), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n738), .B1(new_n741), .B2(new_n747), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(KEYINPUT104), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n704), .B1(new_n758), .B2(new_n748), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n759), .A2(KEYINPUT42), .A3(new_n686), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n756), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G131), .ZN(G33));
  INV_X1    g576(.A(new_n657), .ZN(new_n763));
  AOI211_X1 g577(.A(new_n704), .B(new_n763), .C1(new_n758), .C2(new_n748), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(new_n249), .ZN(G36));
  OR2_X1    g579(.A1(new_n746), .A2(KEYINPUT45), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n746), .A2(KEYINPUT45), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n766), .A2(G469), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n593), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT46), .ZN(new_n770));
  OAI21_X1  g584(.A(KEYINPUT105), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT105), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n768), .A2(new_n772), .A3(KEYINPUT46), .A4(new_n593), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  AOI22_X1  g588(.A1(new_n769), .A2(new_n770), .B1(new_n591), .B2(new_n693), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n689), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n776), .A2(new_n662), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT43), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(KEYINPUT106), .ZN(new_n779));
  XOR2_X1   g593(.A(KEYINPUT106), .B(KEYINPUT43), .Z(new_n780));
  INV_X1    g594(.A(new_n622), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n611), .A2(new_n781), .ZN(new_n782));
  MUX2_X1   g596(.A(new_n779), .B(new_n780), .S(new_n782), .Z(new_n783));
  AOI21_X1  g597(.A(new_n602), .B1(new_n644), .B2(new_n642), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n783), .A2(KEYINPUT44), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(KEYINPUT44), .B1(new_n783), .B2(new_n784), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n665), .A2(new_n401), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n785), .A2(new_n786), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n777), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G137), .ZN(G39));
  NOR3_X1   g605(.A1(new_n788), .A2(new_n477), .A3(new_n521), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(new_n686), .ZN(new_n793));
  XOR2_X1   g607(.A(new_n793), .B(KEYINPUT107), .Z(new_n794));
  NOR2_X1   g608(.A1(new_n776), .A2(KEYINPUT47), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT47), .ZN(new_n796));
  AOI211_X1 g610(.A(new_n796), .B(new_n689), .C1(new_n774), .C2(new_n775), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n794), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G140), .ZN(G42));
  INV_X1    g613(.A(new_n654), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n729), .A2(new_n800), .A3(new_n738), .ZN(new_n801));
  AND4_X1   g615(.A1(new_n521), .A2(new_n801), .A3(new_n675), .A4(new_n676), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n622), .B1(new_n248), .B2(new_n299), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n703), .A2(new_n612), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n783), .A2(new_n521), .A3(new_n800), .A4(new_n718), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n801), .A2(new_n783), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(new_n705), .ZN(new_n809));
  OR2_X1    g623(.A1(new_n809), .A2(KEYINPUT48), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(KEYINPUT48), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n807), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n610), .A2(new_n781), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n645), .A2(new_n718), .ZN(new_n814));
  AOI22_X1  g628(.A1(new_n802), .A2(new_n813), .B1(new_n814), .B2(new_n808), .ZN(new_n815));
  INV_X1    g629(.A(new_n729), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n816), .A2(new_n596), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n795), .A2(new_n797), .A3(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n806), .A2(new_n788), .ZN(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n815), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n703), .A2(new_n401), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT111), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n806), .A2(new_n666), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n824), .A2(new_n825), .A3(KEYINPUT50), .ZN(new_n826));
  AOI21_X1  g640(.A(KEYINPUT50), .B1(new_n824), .B2(new_n825), .ZN(new_n827));
  OAI21_X1  g641(.A(KEYINPUT51), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n812), .B1(new_n821), .B2(new_n828), .ZN(new_n829));
  OR2_X1    g643(.A1(new_n818), .A2(new_n820), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT112), .ZN(new_n831));
  OR3_X1    g645(.A1(new_n826), .A2(new_n827), .A3(new_n831), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n831), .B1(new_n826), .B2(new_n827), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n830), .A2(new_n832), .A3(new_n833), .A4(new_n815), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT51), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n829), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n703), .B(new_n705), .C1(new_n623), .C2(new_n629), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n713), .B(new_n837), .C1(new_n730), .C2(new_n731), .ZN(new_n838));
  OAI22_X1  g652(.A1(new_n597), .A2(new_n522), .B1(new_n633), .B2(new_n646), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n627), .A2(new_n803), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n603), .A2(new_n403), .A3(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n712), .A2(new_n660), .A3(new_n655), .A4(new_n787), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n734), .B1(new_n749), .B2(new_n753), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n838), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n764), .B1(new_n756), .B2(new_n760), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT110), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n656), .A2(new_n689), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n636), .A2(new_n641), .A3(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n677), .A2(new_n752), .A3(new_n851), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n722), .A2(new_n724), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n848), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n850), .B1(new_n675), .B2(new_n676), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n722), .A2(new_n724), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n855), .A2(new_n856), .A3(KEYINPUT110), .A4(new_n752), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n650), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n859), .B(new_n660), .C1(new_n657), .C2(new_n686), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n735), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g675(.A(KEYINPUT52), .B1(new_n858), .B2(new_n861), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n735), .A2(new_n860), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n854), .A2(new_n857), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT52), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n846), .A2(new_n847), .A3(new_n862), .A4(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT53), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n865), .B1(new_n863), .B2(new_n864), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n872), .A2(KEYINPUT53), .A3(new_n847), .A4(new_n846), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT54), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n869), .A2(new_n873), .A3(KEYINPUT54), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n836), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g693(.A(G953), .B1(new_n879), .B2(KEYINPUT113), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT113), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n398), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n816), .A2(KEYINPUT49), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n883), .B(KEYINPUT109), .Z(new_n884));
  NAND2_X1  g698(.A1(new_n816), .A2(KEYINPUT49), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n666), .A2(new_n677), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n521), .A2(new_n596), .A3(new_n400), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n782), .A2(new_n887), .ZN(new_n888));
  XOR2_X1   g702(.A(new_n888), .B(KEYINPUT108), .Z(new_n889));
  NAND4_X1  g703(.A1(new_n884), .A2(new_n885), .A3(new_n886), .A4(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n880), .A2(new_n882), .A3(new_n890), .ZN(G75));
  NOR2_X1   g705(.A1(new_n397), .A2(G952), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n187), .B1(new_n869), .B2(new_n873), .ZN(new_n893));
  AOI21_X1  g707(.A(KEYINPUT56), .B1(new_n893), .B2(new_n386), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n379), .A2(new_n382), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(new_n380), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT55), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  OR3_X1    g712(.A1(new_n894), .A2(KEYINPUT114), .A3(new_n897), .ZN(new_n899));
  OAI21_X1  g713(.A(KEYINPUT114), .B1(new_n894), .B2(new_n897), .ZN(new_n900));
  AOI211_X1 g714(.A(new_n892), .B(new_n898), .C1(new_n899), .C2(new_n900), .ZN(G51));
  INV_X1    g715(.A(new_n768), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n874), .A2(G902), .A3(new_n902), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT117), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n590), .B(KEYINPUT115), .Z(new_n905));
  AND3_X1   g719(.A1(new_n869), .A2(KEYINPUT54), .A3(new_n873), .ZN(new_n906));
  AOI21_X1  g720(.A(KEYINPUT54), .B1(new_n869), .B2(new_n873), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n593), .B(KEYINPUT57), .Z(new_n909));
  AOI21_X1  g723(.A(new_n905), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n904), .B1(new_n910), .B2(KEYINPUT116), .ZN(new_n911));
  OR2_X1    g725(.A1(new_n910), .A2(KEYINPUT116), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n892), .B1(new_n911), .B2(new_n912), .ZN(G54));
  INV_X1    g727(.A(new_n892), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n893), .A2(KEYINPUT58), .A3(G475), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n914), .B1(new_n915), .B2(new_n293), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n916), .B1(new_n293), .B2(new_n915), .ZN(G60));
  INV_X1    g731(.A(KEYINPUT119), .ZN(new_n918));
  OR2_X1    g732(.A1(new_n615), .A2(new_n618), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  XNOR2_X1  g734(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(new_n620), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n906), .A2(new_n907), .A3(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n918), .B1(new_n924), .B2(new_n892), .ZN(new_n925));
  OAI211_X1 g739(.A(KEYINPUT119), .B(new_n914), .C1(new_n878), .C2(new_n923), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n876), .A2(new_n877), .A3(new_n922), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n919), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n925), .A2(new_n926), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(KEYINPUT120), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT120), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n925), .A2(new_n926), .A3(new_n931), .A4(new_n928), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n930), .A2(new_n932), .ZN(G63));
  NAND2_X1  g747(.A1(G217), .A2(G902), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT121), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT60), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n874), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n638), .A2(new_n639), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n874), .A2(new_n936), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n892), .B1(new_n940), .B2(new_n510), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n939), .A2(new_n941), .A3(KEYINPUT61), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT123), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n939), .A2(new_n941), .A3(KEYINPUT123), .A4(KEYINPUT61), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT122), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n939), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n937), .A2(KEYINPUT122), .A3(new_n938), .ZN(new_n949));
  AND3_X1   g763(.A1(new_n948), .A2(new_n949), .A3(new_n941), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n946), .B1(KEYINPUT61), .B2(new_n950), .ZN(G66));
  OAI21_X1  g765(.A(G953), .B1(new_n396), .B2(new_n325), .ZN(new_n952));
  INV_X1    g766(.A(new_n842), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n838), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n952), .B1(new_n954), .B2(G953), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n895), .B1(G898), .B2(new_n397), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(G69));
  XOR2_X1   g771(.A(new_n446), .B(new_n287), .Z(new_n958));
  AOI21_X1  g772(.A(new_n958), .B1(G900), .B2(G953), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n863), .B(KEYINPUT124), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n960), .B1(new_n777), .B2(new_n789), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT126), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n777), .A2(new_n705), .A3(new_n856), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n963), .A2(new_n798), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n962), .A2(new_n847), .A3(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n959), .B1(new_n965), .B2(G953), .ZN(new_n966));
  OAI21_X1  g780(.A(KEYINPUT62), .B1(new_n960), .B2(new_n684), .ZN(new_n967));
  NOR4_X1   g781(.A1(new_n663), .A2(new_n704), .A3(new_n788), .A4(new_n840), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n967), .A2(new_n790), .A3(new_n798), .A4(new_n969), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n960), .A2(new_n684), .A3(KEYINPUT62), .ZN(new_n971));
  OR3_X1    g785(.A1(new_n970), .A2(KEYINPUT125), .A3(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(KEYINPUT125), .B1(new_n970), .B2(new_n971), .ZN(new_n973));
  AOI21_X1  g787(.A(G953), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(new_n958), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n966), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OAI221_X1 g790(.A(G953), .B1(new_n524), .B2(new_n652), .C1(new_n958), .C2(KEYINPUT127), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n966), .B(new_n977), .C1(new_n974), .C2(new_n975), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n980), .ZN(G72));
  AND3_X1   g795(.A1(new_n972), .A2(new_n954), .A3(new_n973), .ZN(new_n982));
  NAND2_X1  g796(.A1(G472), .A2(G902), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(KEYINPUT63), .Z(new_n984));
  INV_X1    g798(.A(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n667), .B1(new_n982), .B2(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(new_n954), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n984), .B1(new_n965), .B2(new_n987), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n988), .A2(new_n409), .A3(new_n452), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n409), .B1(new_n461), .B2(new_n451), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n985), .B1(new_n448), .B2(new_n990), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n892), .B1(new_n874), .B2(new_n991), .ZN(new_n992));
  AND3_X1   g806(.A1(new_n986), .A2(new_n989), .A3(new_n992), .ZN(G57));
endmodule


