//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 0 0 1 1 1 0 0 1 1 1 1 1 0 1 1 1 0 1 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 0 0 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:24 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  XNOR2_X1  g0001(.A(new_n201), .B(KEYINPUT64), .ZN(new_n202));
  NOR2_X1   g0002(.A1(new_n202), .A2(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G116), .A2(G270), .ZN(new_n208));
  INV_X1    g0008(.A(G50), .ZN(new_n209));
  INV_X1    g0009(.A(G226), .ZN(new_n210));
  OAI21_X1  g0010(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  XNOR2_X1  g0011(.A(KEYINPUT66), .B(G77), .ZN(new_n212));
  AND2_X1   g0012(.A1(new_n212), .A2(G244), .ZN(new_n213));
  INV_X1    g0013(.A(G68), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(KEYINPUT65), .ZN(new_n215));
  INV_X1    g0015(.A(KEYINPUT65), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G68), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  AOI211_X1 g0018(.A(new_n211), .B(new_n213), .C1(G238), .C2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT67), .Z(new_n223));
  AOI21_X1  g0023(.A(new_n207), .B1(new_n219), .B2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(KEYINPUT1), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT68), .ZN(new_n227));
  NOR2_X1   g0027(.A1(G58), .A2(G68), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(G50), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(G1), .A2(G13), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n232), .A2(new_n206), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  INV_X1    g0034(.A(G13), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n207), .A2(new_n235), .ZN(new_n236));
  INV_X1    g0036(.A(new_n236), .ZN(new_n237));
  OAI211_X1 g0037(.A(new_n237), .B(G250), .C1(G257), .C2(G264), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT0), .ZN(new_n239));
  OAI211_X1 g0039(.A(new_n234), .B(new_n239), .C1(new_n224), .C2(new_n225), .ZN(new_n240));
  NOR2_X1   g0040(.A1(new_n227), .A2(new_n240), .ZN(G361));
  XNOR2_X1  g0041(.A(G238), .B(G244), .ZN(new_n242));
  INV_X1    g0042(.A(G232), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(KEYINPUT2), .B(G226), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G264), .B(G270), .Z(new_n247));
  XNOR2_X1  g0047(.A(G250), .B(G257), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G358));
  XNOR2_X1  g0050(.A(G87), .B(G97), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(KEYINPUT69), .ZN(new_n252));
  XOR2_X1   g0052(.A(G107), .B(G116), .Z(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XOR2_X1   g0054(.A(G68), .B(G77), .Z(new_n255));
  XOR2_X1   g0055(.A(G50), .B(G58), .Z(new_n256));
  XNOR2_X1  g0056(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n254), .B(new_n257), .ZN(G351));
  INV_X1    g0058(.A(G41), .ZN(new_n259));
  INV_X1    g0059(.A(G45), .ZN(new_n260));
  AOI21_X1  g0060(.A(G1), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(G33), .A2(G41), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n262), .A2(G1), .A3(G13), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n261), .A2(new_n263), .A3(G274), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n265), .B1(G238), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(G33), .A2(G97), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT3), .B(G33), .ZN(new_n271));
  INV_X1    g0071(.A(G1698), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n270), .B1(new_n273), .B2(new_n210), .ZN(new_n274));
  OR2_X1    g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n272), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n274), .B1(G232), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n269), .B1(new_n278), .B2(new_n263), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT13), .ZN(new_n280));
  XNOR2_X1  g0080(.A(new_n279), .B(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G169), .ZN(new_n282));
  OAI21_X1  g0082(.A(KEYINPUT14), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  XNOR2_X1  g0083(.A(new_n279), .B(KEYINPUT13), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT14), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n284), .A2(new_n285), .A3(G169), .ZN(new_n286));
  INV_X1    g0086(.A(G179), .ZN(new_n287));
  OAI211_X1 g0087(.A(new_n283), .B(new_n286), .C1(new_n287), .C2(new_n284), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT12), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n290));
  NOR3_X1   g0090(.A1(new_n218), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n290), .ZN(new_n292));
  AOI21_X1  g0092(.A(KEYINPUT12), .B1(new_n292), .B2(new_n214), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(new_n232), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n292), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n205), .A2(G20), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n297), .A2(G68), .A3(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G33), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n300), .A2(G20), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G77), .ZN(new_n303));
  NOR2_X1   g0103(.A1(G20), .A2(G33), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  OAI22_X1  g0105(.A1(new_n302), .A2(new_n303), .B1(new_n209), .B2(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n218), .A2(new_n206), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n296), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT11), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n294), .B(new_n299), .C1(new_n308), .C2(new_n309), .ZN(new_n310));
  AND2_X1   g0110(.A1(new_n308), .A2(new_n309), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n288), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n284), .A2(G200), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n281), .A2(G190), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n315), .A2(new_n316), .A3(new_n312), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n202), .A2(G20), .ZN(new_n319));
  XOR2_X1   g0119(.A(KEYINPUT8), .B(G58), .Z(new_n320));
  AOI22_X1  g0120(.A1(new_n320), .A2(new_n301), .B1(G150), .B2(new_n304), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n319), .A2(new_n321), .B1(new_n232), .B2(new_n295), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n297), .A2(G50), .A3(new_n298), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n323), .B1(G50), .B2(new_n290), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  AND2_X1   g0126(.A1(KEYINPUT3), .A2(G33), .ZN(new_n327));
  NOR2_X1   g0127(.A1(KEYINPUT3), .A2(G33), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n277), .A2(G223), .B1(new_n329), .B2(new_n212), .ZN(new_n330));
  INV_X1    g0130(.A(G222), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n330), .B1(new_n331), .B2(new_n273), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n232), .B1(G33), .B2(G41), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n265), .B1(G226), .B2(new_n268), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n326), .B1(new_n337), .B2(G169), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n336), .A2(G179), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT9), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n341), .A2(new_n326), .B1(new_n337), .B2(G190), .ZN(new_n342));
  AOI22_X1  g0142(.A1(KEYINPUT9), .A2(new_n325), .B1(new_n336), .B2(G200), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT10), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT10), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n342), .A2(new_n346), .A3(new_n343), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n340), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n277), .A2(G238), .ZN(new_n349));
  INV_X1    g0149(.A(G107), .ZN(new_n350));
  OAI221_X1 g0150(.A(new_n349), .B1(new_n350), .B2(new_n271), .C1(new_n243), .C2(new_n273), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n333), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n265), .B1(G244), .B2(new_n268), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(G200), .ZN(new_n355));
  XNOR2_X1  g0155(.A(KEYINPUT15), .B(G87), .ZN(new_n356));
  OAI21_X1  g0156(.A(KEYINPUT70), .B1(new_n356), .B2(new_n302), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n212), .A2(G20), .ZN(new_n358));
  INV_X1    g0158(.A(new_n320), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n357), .B(new_n358), .C1(new_n359), .C2(new_n305), .ZN(new_n360));
  NOR3_X1   g0160(.A1(new_n356), .A2(new_n302), .A3(KEYINPUT70), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n296), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n298), .A2(G77), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n212), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n297), .A2(new_n364), .B1(new_n365), .B2(new_n292), .ZN(new_n366));
  AND2_X1   g0166(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(G190), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n355), .B(new_n367), .C1(new_n368), .C2(new_n354), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n367), .B1(new_n282), .B2(new_n354), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n352), .A2(new_n287), .A3(new_n353), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n348), .A2(new_n369), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n210), .A2(G1698), .ZN(new_n374));
  OAI221_X1 g0174(.A(new_n374), .B1(G223), .B2(G1698), .C1(new_n327), .C2(new_n328), .ZN(new_n375));
  NAND2_X1  g0175(.A1(G33), .A2(G87), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n333), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n264), .B1(new_n243), .B2(new_n267), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n378), .A2(new_n380), .A3(G179), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n263), .B1(new_n375), .B2(new_n376), .ZN(new_n382));
  OAI21_X1  g0182(.A(G169), .B1(new_n382), .B2(new_n379), .ZN(new_n383));
  AND3_X1   g0183(.A1(new_n381), .A2(KEYINPUT73), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(KEYINPUT73), .B1(new_n381), .B2(new_n383), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT18), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT16), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT71), .ZN(new_n389));
  INV_X1    g0189(.A(G159), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n389), .B1(new_n305), .B2(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n304), .A2(KEYINPUT71), .A3(G159), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n228), .B1(new_n218), .B2(G58), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n393), .B1(new_n394), .B2(new_n206), .ZN(new_n395));
  XNOR2_X1  g0195(.A(KEYINPUT65), .B(G68), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT7), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n397), .B1(new_n271), .B2(G20), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n329), .A2(KEYINPUT7), .A3(new_n206), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n396), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n388), .B1(new_n395), .B2(new_n400), .ZN(new_n401));
  NOR3_X1   g0201(.A1(new_n271), .A2(new_n397), .A3(G20), .ZN(new_n402));
  AOI21_X1  g0202(.A(KEYINPUT7), .B1(new_n329), .B2(new_n206), .ZN(new_n403));
  OAI21_X1  g0203(.A(G68), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(G58), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n229), .B1(new_n396), .B2(new_n405), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n406), .A2(G20), .B1(new_n391), .B2(new_n392), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n404), .A2(new_n407), .A3(KEYINPUT16), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n401), .A2(new_n408), .A3(new_n296), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n320), .A2(new_n298), .ZN(new_n410));
  AOI211_X1 g0210(.A(new_n296), .B(new_n292), .C1(new_n410), .C2(KEYINPUT72), .ZN(new_n411));
  OR2_X1    g0211(.A1(new_n410), .A2(KEYINPUT72), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n411), .A2(new_n412), .B1(new_n292), .B2(new_n359), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n409), .A2(new_n413), .ZN(new_n414));
  AND3_X1   g0214(.A1(new_n386), .A2(new_n387), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n387), .B1(new_n386), .B2(new_n414), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(G200), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n418), .B1(new_n378), .B2(new_n380), .ZN(new_n419));
  NOR3_X1   g0219(.A1(new_n382), .A2(new_n379), .A3(new_n368), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n409), .A2(new_n421), .A3(new_n413), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT17), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n409), .A2(new_n421), .A3(KEYINPUT17), .A4(new_n413), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n424), .A2(KEYINPUT74), .A3(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(KEYINPUT74), .B1(new_n424), .B2(new_n425), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n417), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NOR3_X1   g0229(.A1(new_n318), .A2(new_n373), .A3(new_n429), .ZN(new_n430));
  OAI211_X1 g0230(.A(G250), .B(G1698), .C1(new_n327), .C2(new_n328), .ZN(new_n431));
  NAND2_X1  g0231(.A1(G33), .A2(G283), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OAI211_X1 g0233(.A(G244), .B(new_n272), .C1(new_n327), .C2(new_n328), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT75), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n433), .B1(KEYINPUT4), .B2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT4), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n434), .A2(new_n435), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n263), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n260), .A2(G1), .ZN(new_n441));
  AND2_X1   g0241(.A1(KEYINPUT5), .A2(G41), .ZN(new_n442));
  NOR2_X1   g0242(.A1(KEYINPUT5), .A2(G41), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n444), .A2(G257), .A3(new_n263), .ZN(new_n445));
  INV_X1    g0245(.A(G274), .ZN(new_n446));
  AND2_X1   g0246(.A1(G1), .A2(G13), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n446), .B1(new_n447), .B2(new_n262), .ZN(new_n448));
  XNOR2_X1  g0248(.A(KEYINPUT5), .B(G41), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n448), .A2(new_n441), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n445), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT76), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n445), .A2(new_n450), .A3(KEYINPUT76), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(G200), .B1(new_n440), .B2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(G97), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n292), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n205), .A2(G33), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n290), .A2(new_n459), .A3(new_n232), .A4(new_n295), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n458), .B1(new_n460), .B2(new_n457), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n350), .B1(new_n398), .B2(new_n399), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  XNOR2_X1  g0263(.A(G97), .B(G107), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT6), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NOR3_X1   g0266(.A1(new_n465), .A2(new_n457), .A3(G107), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n469), .A2(G20), .B1(G77), .B2(new_n304), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n463), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n461), .B1(new_n471), .B2(new_n296), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n436), .A2(KEYINPUT4), .ZN(new_n473));
  INV_X1    g0273(.A(new_n433), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n473), .A2(new_n439), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n333), .ZN(new_n476));
  INV_X1    g0276(.A(new_n451), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n476), .A2(G190), .A3(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n456), .A2(new_n472), .A3(new_n478), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n282), .B1(new_n440), .B2(new_n451), .ZN(new_n480));
  AND3_X1   g0280(.A1(new_n445), .A2(KEYINPUT76), .A3(new_n450), .ZN(new_n481));
  AOI21_X1  g0281(.A(KEYINPUT76), .B1(new_n445), .B2(new_n450), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n476), .A2(new_n483), .A3(new_n287), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n467), .B1(new_n465), .B2(new_n464), .ZN(new_n485));
  OAI22_X1  g0285(.A1(new_n485), .A2(new_n206), .B1(new_n303), .B2(new_n305), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n296), .B1(new_n486), .B2(new_n462), .ZN(new_n487));
  INV_X1    g0287(.A(new_n461), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n480), .A2(new_n484), .A3(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT19), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n491), .B1(new_n302), .B2(new_n457), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n271), .A2(new_n206), .A3(G68), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  XOR2_X1   g0294(.A(KEYINPUT78), .B(G87), .Z(new_n495));
  NOR2_X1   g0295(.A1(G97), .A2(G107), .ZN(new_n496));
  NAND3_X1  g0296(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n495), .A2(new_n496), .B1(new_n206), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n296), .B1(new_n494), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n356), .A2(new_n292), .ZN(new_n500));
  INV_X1    g0300(.A(G87), .ZN(new_n501));
  OR2_X1    g0301(.A1(new_n460), .A2(new_n501), .ZN(new_n502));
  AND3_X1   g0302(.A1(new_n499), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  OAI211_X1 g0303(.A(G244), .B(G1698), .C1(new_n327), .C2(new_n328), .ZN(new_n504));
  OAI211_X1 g0304(.A(G238), .B(new_n272), .C1(new_n327), .C2(new_n328), .ZN(new_n505));
  NAND2_X1  g0305(.A1(G33), .A2(G116), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(G250), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n508), .B1(new_n260), .B2(G1), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n205), .A2(new_n446), .A3(G45), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n263), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(KEYINPUT77), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT77), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n263), .A2(new_n509), .A3(new_n510), .A4(new_n513), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n333), .A2(new_n507), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(G190), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n503), .B(new_n516), .C1(new_n418), .C2(new_n515), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n479), .A2(new_n490), .A3(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT25), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n292), .A2(new_n519), .A3(new_n350), .ZN(new_n520));
  OAI21_X1  g0320(.A(KEYINPUT25), .B1(new_n290), .B2(G107), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n520), .B(new_n521), .C1(new_n350), .C2(new_n460), .ZN(new_n522));
  XNOR2_X1  g0322(.A(new_n522), .B(KEYINPUT84), .ZN(new_n523));
  AND3_X1   g0323(.A1(new_n350), .A2(KEYINPUT23), .A3(G20), .ZN(new_n524));
  AOI21_X1  g0324(.A(KEYINPUT23), .B1(new_n350), .B2(G20), .ZN(new_n525));
  OAI22_X1  g0325(.A1(new_n524), .A2(new_n525), .B1(G20), .B2(new_n506), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n206), .B(G87), .C1(new_n327), .C2(new_n328), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(KEYINPUT22), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT22), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n271), .A2(new_n529), .A3(new_n206), .A4(G87), .ZN(new_n530));
  AOI211_X1 g0330(.A(KEYINPUT24), .B(new_n526), .C1(new_n528), .C2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT24), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n528), .A2(new_n530), .ZN(new_n533));
  INV_X1    g0333(.A(new_n526), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n296), .B1(new_n531), .B2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT83), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n523), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  OAI211_X1 g0338(.A(KEYINPUT83), .B(new_n296), .C1(new_n531), .C2(new_n535), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  OAI211_X1 g0341(.A(G250), .B(new_n272), .C1(new_n327), .C2(new_n328), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT85), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n271), .A2(KEYINPUT85), .A3(G250), .A4(new_n272), .ZN(new_n545));
  NAND2_X1  g0345(.A1(G33), .A2(G294), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n271), .A2(G257), .A3(G1698), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n544), .A2(new_n545), .A3(new_n546), .A4(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n333), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n444), .A2(G264), .A3(new_n263), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT86), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n444), .A2(KEYINPUT86), .A3(G264), .A4(new_n263), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n549), .A2(new_n450), .A3(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT87), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n548), .A2(new_n333), .B1(new_n552), .B2(new_n553), .ZN(new_n558));
  AOI21_X1  g0358(.A(KEYINPUT87), .B1(new_n558), .B2(new_n450), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n368), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n555), .A2(new_n418), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n518), .B1(new_n541), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n555), .A2(new_n556), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n558), .A2(KEYINPUT87), .A3(new_n450), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n564), .A2(G169), .A3(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n558), .A2(G179), .A3(new_n450), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n566), .A2(new_n567), .B1(new_n538), .B2(new_n539), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n449), .A2(new_n441), .B1(new_n447), .B2(new_n262), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n205), .A2(G45), .ZN(new_n570));
  INV_X1    g0370(.A(new_n443), .ZN(new_n571));
  NAND2_X1  g0371(.A1(KEYINPUT5), .A2(G41), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n569), .A2(G270), .B1(new_n448), .B2(new_n573), .ZN(new_n574));
  OAI211_X1 g0374(.A(G264), .B(G1698), .C1(new_n327), .C2(new_n328), .ZN(new_n575));
  OAI211_X1 g0375(.A(G257), .B(new_n272), .C1(new_n327), .C2(new_n328), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n275), .A2(G303), .A3(new_n276), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n333), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n282), .B1(new_n574), .B2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(G116), .ZN(new_n581));
  OR3_X1    g0381(.A1(new_n460), .A2(KEYINPUT79), .A3(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(KEYINPUT79), .B1(new_n460), .B2(new_n581), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n295), .A2(new_n232), .B1(G20), .B2(new_n581), .ZN(new_n585));
  AOI21_X1  g0385(.A(G20), .B1(G33), .B2(G283), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n300), .A2(G97), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT80), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n588), .B1(new_n586), .B2(new_n587), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n585), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT81), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT20), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n292), .A2(new_n581), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n584), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  OAI211_X1 g0397(.A(KEYINPUT20), .B(new_n585), .C1(new_n590), .C2(new_n591), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(KEYINPUT81), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n432), .B(new_n206), .C1(G33), .C2(new_n457), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(KEYINPUT80), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n589), .ZN(new_n602));
  AOI21_X1  g0402(.A(KEYINPUT20), .B1(new_n602), .B2(new_n585), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n580), .B1(new_n597), .B2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT21), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OAI211_X1 g0407(.A(KEYINPUT21), .B(new_n580), .C1(new_n597), .C2(new_n604), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n574), .A2(new_n579), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  OAI211_X1 g0410(.A(G179), .B(new_n610), .C1(new_n597), .C2(new_n604), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n607), .A2(new_n608), .A3(new_n611), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n568), .A2(new_n612), .ZN(new_n613));
  OR2_X1    g0413(.A1(new_n515), .A2(G169), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n499), .B(new_n500), .C1(new_n356), .C2(new_n460), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n515), .A2(new_n287), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n584), .A2(new_n595), .A3(new_n596), .ZN(new_n619));
  OR2_X1    g0419(.A1(new_n599), .A2(new_n603), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n609), .A2(G200), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT82), .ZN(new_n623));
  OR2_X1    g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n622), .A2(new_n623), .B1(G190), .B2(new_n610), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n618), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  AND4_X1   g0426(.A1(new_n430), .A2(new_n563), .A3(new_n613), .A4(new_n626), .ZN(G372));
  NAND2_X1  g0427(.A1(new_n517), .A2(new_n617), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n490), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n629), .A2(KEYINPUT26), .A3(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT26), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n632), .B1(new_n628), .B2(new_n490), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n618), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n563), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n634), .B1(new_n635), .B2(new_n613), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n430), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g0437(.A(new_n637), .B(KEYINPUT88), .Z(new_n638));
  INV_X1    g0438(.A(new_n317), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n314), .B1(new_n639), .B2(new_n372), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n640), .B1(new_n428), .B2(new_n427), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n381), .A2(new_n383), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n414), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g0443(.A(new_n643), .B(new_n387), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n345), .A2(new_n347), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n340), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n638), .A2(new_n647), .ZN(G369));
  NAND3_X1  g0448(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n649));
  OR2_X1    g0449(.A1(new_n649), .A2(KEYINPUT27), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(KEYINPUT27), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n650), .A2(G213), .A3(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(G343), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n655), .B1(new_n619), .B2(new_n620), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n612), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n624), .A2(new_n625), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n612), .A2(new_n656), .ZN(new_n660));
  OAI21_X1  g0460(.A(G330), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n562), .A2(new_n541), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n540), .A2(new_n654), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n568), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n568), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n666), .A2(new_n654), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n662), .A2(KEYINPUT89), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT89), .ZN(new_n670));
  INV_X1    g0470(.A(new_n668), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n670), .B1(new_n671), .B2(new_n661), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n667), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n612), .A2(new_n655), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n674), .B1(new_n665), .B2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n673), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g0478(.A(new_n678), .B(KEYINPUT90), .Z(G399));
  NAND3_X1  g0479(.A1(new_n495), .A2(new_n581), .A3(new_n496), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n236), .A2(G41), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n681), .A2(new_n683), .A3(G1), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n684), .B1(new_n230), .B2(new_n683), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(KEYINPUT28), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n636), .A2(new_n655), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n687), .A2(KEYINPUT29), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(KEYINPUT29), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(G330), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n563), .A2(new_n613), .A3(new_n626), .A4(new_n655), .ZN(new_n692));
  XOR2_X1   g0492(.A(KEYINPUT93), .B(KEYINPUT30), .Z(new_n693));
  NAND3_X1  g0493(.A1(new_n574), .A2(new_n579), .A3(G179), .ZN(new_n694));
  NOR3_X1   g0494(.A1(new_n440), .A2(new_n694), .A3(new_n451), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n549), .A2(new_n554), .A3(new_n515), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT91), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n558), .A2(KEYINPUT91), .A3(new_n515), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n695), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(KEYINPUT92), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT92), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n695), .A2(new_n698), .A3(new_n702), .A4(new_n699), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n693), .B1(new_n701), .B2(new_n703), .ZN(new_n704));
  NOR3_X1   g0504(.A1(new_n610), .A2(G179), .A3(new_n515), .ZN(new_n705));
  OAI211_X1 g0505(.A(new_n705), .B(new_n555), .C1(new_n440), .C2(new_n455), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT30), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n706), .B1(new_n700), .B2(new_n707), .ZN(new_n708));
  OAI211_X1 g0508(.A(KEYINPUT31), .B(new_n654), .C1(new_n704), .C2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n692), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n654), .B1(new_n704), .B2(new_n708), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT31), .ZN(new_n712));
  AOI21_X1  g0512(.A(KEYINPUT94), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n711), .A2(KEYINPUT94), .A3(new_n712), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n691), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n690), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n686), .B1(new_n717), .B2(G1), .ZN(G364));
  NOR2_X1   g0518(.A1(new_n235), .A2(G20), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n205), .B1(new_n719), .B2(G45), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n682), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n662), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n660), .B1(new_n658), .B2(new_n657), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n723), .B1(G330), .B2(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n232), .B1(G20), .B2(new_n282), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n206), .A2(new_n287), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(G200), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(new_n368), .ZN(new_n731));
  XNOR2_X1  g0531(.A(new_n731), .B(KEYINPUT97), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n206), .A2(G179), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n734), .A2(G190), .A3(G200), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n735), .B(KEYINPUT98), .ZN(new_n736));
  AOI22_X1  g0536(.A1(new_n733), .A2(G326), .B1(G303), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(G190), .A2(G200), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n729), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(G311), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n734), .A2(new_n738), .ZN(new_n741));
  INV_X1    g0541(.A(G329), .ZN(new_n742));
  OAI22_X1  g0542(.A1(new_n739), .A2(new_n740), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n729), .A2(G190), .A3(new_n418), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  AOI211_X1 g0545(.A(new_n271), .B(new_n743), .C1(G322), .C2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n730), .A2(G190), .ZN(new_n747));
  INV_X1    g0547(.A(G317), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(KEYINPUT33), .ZN(new_n749));
  OR2_X1    g0549(.A1(new_n748), .A2(KEYINPUT33), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n747), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n368), .A2(G179), .A3(G200), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(new_n206), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n734), .A2(new_n368), .A3(G200), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI22_X1  g0556(.A1(new_n754), .A2(G294), .B1(new_n756), .B2(G283), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n737), .A2(new_n746), .A3(new_n751), .A4(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n747), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT32), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n741), .A2(new_n390), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n759), .A2(new_n214), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n760), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n763), .B1(new_n495), .B2(new_n735), .ZN(new_n764));
  OAI221_X1 g0564(.A(new_n271), .B1(new_n744), .B2(new_n405), .C1(new_n365), .C2(new_n739), .ZN(new_n765));
  NOR3_X1   g0565(.A1(new_n762), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n755), .A2(new_n350), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n767), .B1(G50), .B2(new_n731), .ZN(new_n768));
  OAI211_X1 g0568(.A(new_n766), .B(new_n768), .C1(new_n457), .C2(new_n753), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n728), .B1(new_n758), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G13), .A2(G33), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(G20), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n727), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n257), .A2(G45), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n236), .A2(new_n271), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n778), .B1(new_n260), .B2(new_n231), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n237), .A2(new_n271), .ZN(new_n780));
  INV_X1    g0580(.A(G355), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n780), .A2(new_n781), .B1(G116), .B2(new_n237), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n776), .A2(new_n779), .B1(new_n782), .B2(KEYINPUT96), .ZN(new_n783));
  OR2_X1    g0583(.A1(new_n782), .A2(KEYINPUT96), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n775), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n722), .B(KEYINPUT95), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n770), .A2(new_n785), .A3(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n773), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n788), .B1(new_n725), .B2(new_n789), .ZN(new_n790));
  AND2_X1   g0590(.A1(new_n726), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(G396));
  NOR2_X1   g0592(.A1(new_n372), .A2(new_n654), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n369), .B1(new_n367), .B2(new_n655), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n793), .B1(new_n794), .B2(new_n372), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n687), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n636), .A2(new_n655), .A3(new_n795), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n692), .A2(new_n709), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n711), .A2(new_n712), .ZN(new_n801));
  INV_X1    g0601(.A(KEYINPUT94), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n800), .A2(new_n803), .A3(new_n715), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(G330), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n722), .B1(new_n799), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n806), .B1(new_n805), .B2(new_n799), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n728), .A2(new_n772), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n786), .B1(G77), .B2(new_n808), .ZN(new_n809));
  XOR2_X1   g0609(.A(new_n809), .B(KEYINPUT99), .Z(new_n810));
  INV_X1    g0610(.A(new_n741), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n271), .B1(new_n811), .B2(G311), .ZN(new_n812));
  INV_X1    g0612(.A(G294), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n812), .B1(new_n581), .B2(new_n739), .C1(new_n813), .C2(new_n744), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n754), .A2(G97), .B1(new_n756), .B2(G87), .ZN(new_n815));
  INV_X1    g0615(.A(G283), .ZN(new_n816));
  INV_X1    g0616(.A(G303), .ZN(new_n817));
  INV_X1    g0617(.A(new_n731), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n815), .B1(new_n816), .B2(new_n759), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n814), .B(new_n819), .C1(G107), .C2(new_n736), .ZN(new_n820));
  INV_X1    g0620(.A(G132), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n271), .B1(new_n741), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(G68), .B2(new_n756), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n405), .B2(new_n753), .ZN(new_n824));
  INV_X1    g0624(.A(new_n739), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n745), .A2(G143), .B1(new_n825), .B2(G159), .ZN(new_n826));
  INV_X1    g0626(.A(G137), .ZN(new_n827));
  INV_X1    g0627(.A(G150), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n826), .B1(new_n818), .B2(new_n827), .C1(new_n828), .C2(new_n759), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT34), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n824), .B(new_n831), .C1(G50), .C2(new_n736), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n829), .A2(new_n830), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n820), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n810), .B1(new_n728), .B2(new_n834), .C1(new_n795), .C2(new_n772), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n807), .A2(new_n835), .ZN(G384));
  NOR2_X1   g0636(.A1(new_n719), .A2(new_n205), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n690), .A2(new_n430), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(new_n647), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n839), .B(KEYINPUT102), .ZN(new_n840));
  INV_X1    g0640(.A(new_n793), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n798), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n313), .A2(new_n654), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n314), .A2(new_n317), .A3(new_n843), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n313), .B(new_n654), .C1(new_n639), .C2(new_n288), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n842), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n408), .A2(new_n296), .ZN(new_n848));
  AOI21_X1  g0648(.A(KEYINPUT16), .B1(new_n404), .B2(new_n407), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n413), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n652), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n850), .A2(new_n642), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n852), .A2(new_n853), .A3(new_n422), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n652), .B1(new_n409), .B2(new_n413), .ZN(new_n855));
  INV_X1    g0655(.A(new_n414), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n855), .B1(new_n856), .B2(new_n421), .ZN(new_n857));
  AOI21_X1  g0657(.A(KEYINPUT37), .B1(new_n386), .B2(new_n414), .ZN(new_n858));
  AOI22_X1  g0658(.A1(KEYINPUT37), .A2(new_n854), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n386), .A2(new_n414), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(KEYINPUT18), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n386), .A2(new_n387), .A3(new_n414), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n428), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n864), .B1(new_n865), .B2(new_n426), .ZN(new_n866));
  OAI211_X1 g0666(.A(KEYINPUT38), .B(new_n860), .C1(new_n866), .C2(new_n852), .ZN(new_n867));
  INV_X1    g0667(.A(new_n852), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n429), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(new_n860), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT38), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n847), .B1(new_n867), .B2(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n644), .A2(new_n851), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(KEYINPUT38), .B1(new_n869), .B2(new_n860), .ZN(new_n876));
  AOI211_X1 g0676(.A(new_n871), .B(new_n859), .C1(new_n429), .C2(new_n868), .ZN(new_n877));
  OAI21_X1  g0677(.A(KEYINPUT39), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT39), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n424), .A2(new_n425), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT100), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n424), .A2(KEYINPUT100), .A3(new_n425), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n644), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n857), .A2(new_n858), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n857), .A2(new_n643), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(KEYINPUT37), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n884), .A2(new_n855), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n867), .B(new_n879), .C1(new_n888), .C2(KEYINPUT38), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n878), .A2(KEYINPUT101), .A3(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n288), .A2(new_n313), .A3(new_n655), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n884), .A2(new_n855), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n887), .A2(new_n885), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n871), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT101), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n895), .A2(new_n896), .A3(new_n879), .A4(new_n867), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n890), .A2(new_n892), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n875), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n840), .B(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n895), .A2(new_n867), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n796), .B1(new_n844), .B2(new_n845), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n711), .A2(KEYINPUT103), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT103), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n904), .B(new_n654), .C1(new_n704), .C2(new_n708), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n903), .A2(new_n712), .A3(new_n905), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n906), .A2(KEYINPUT104), .A3(new_n800), .ZN(new_n907));
  AOI21_X1  g0707(.A(KEYINPUT104), .B1(new_n906), .B2(new_n800), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n901), .B(new_n902), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(KEYINPUT40), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n906), .A2(new_n800), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT104), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n906), .A2(new_n800), .A3(KEYINPUT104), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT40), .B1(new_n872), .B2(new_n867), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n915), .A2(new_n902), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n910), .A2(new_n917), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n915), .A2(new_n430), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n691), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n919), .B2(new_n918), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n837), .B1(new_n900), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n900), .B2(new_n921), .ZN(new_n923));
  OR2_X1    g0723(.A1(new_n469), .A2(KEYINPUT35), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n469), .A2(KEYINPUT35), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n924), .A2(G116), .A3(new_n233), .A4(new_n925), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT36), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n209), .B1(new_n394), .B2(new_n212), .ZN(new_n928));
  OAI211_X1 g0728(.A(new_n235), .B(G1), .C1(G50), .C2(G68), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n923), .B(new_n927), .C1(new_n928), .C2(new_n929), .ZN(G367));
  INV_X1    g0730(.A(new_n665), .ZN(new_n931));
  INV_X1    g0731(.A(new_n675), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n931), .A2(new_n674), .A3(new_n932), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n479), .B(new_n490), .C1(new_n472), .C2(new_n655), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n630), .A2(new_n654), .ZN(new_n935));
  AND3_X1   g0735(.A1(new_n934), .A2(new_n935), .A3(KEYINPUT107), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT107), .B1(new_n934), .B2(new_n935), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(KEYINPUT42), .B1(new_n933), .B2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n938), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT42), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n940), .A2(new_n941), .A3(new_n668), .A4(new_n932), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n630), .B1(new_n940), .B2(new_n568), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n939), .B(new_n942), .C1(new_n654), .C2(new_n943), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n503), .A2(new_n655), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n945), .A2(new_n617), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n946), .A2(KEYINPUT105), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(KEYINPUT105), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n629), .A2(new_n945), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(KEYINPUT43), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n944), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(KEYINPUT108), .ZN(new_n953));
  OR2_X1    g0753(.A1(new_n950), .A2(KEYINPUT43), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n954), .B(KEYINPUT106), .Z(new_n955));
  INV_X1    g0755(.A(KEYINPUT108), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n944), .A2(new_n956), .A3(new_n951), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n953), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n955), .B1(new_n953), .B2(new_n957), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n959), .A2(new_n960), .B1(new_n673), .B2(new_n938), .ZN(new_n961));
  INV_X1    g0761(.A(new_n960), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n673), .A2(new_n938), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n962), .A2(new_n958), .A3(new_n963), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n682), .B(KEYINPUT41), .Z(new_n965));
  INV_X1    g0765(.A(KEYINPUT44), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n677), .B2(new_n940), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n676), .A2(new_n938), .A3(KEYINPUT44), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n677), .A2(new_n940), .A3(KEYINPUT45), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT45), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n676), .B2(new_n938), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  AND3_X1   g0773(.A1(new_n969), .A2(new_n673), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n673), .B1(new_n969), .B2(new_n973), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n675), .B1(new_n665), .B2(new_n667), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n933), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n978), .A2(KEYINPUT109), .A3(new_n662), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT109), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n661), .A2(new_n980), .ZN(new_n981));
  OAI211_X1 g0781(.A(KEYINPUT109), .B(G330), .C1(new_n659), .C2(new_n660), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n981), .A2(new_n982), .A3(new_n933), .A4(new_n977), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n979), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n717), .A2(KEYINPUT110), .A3(new_n984), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n984), .A2(new_n689), .A3(new_n688), .A4(new_n805), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT110), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n976), .A2(new_n985), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n965), .B1(new_n989), .B2(new_n717), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n961), .B(new_n964), .C1(new_n990), .C2(new_n721), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n774), .B1(new_n237), .B2(new_n356), .C1(new_n249), .C2(new_n778), .ZN(new_n992));
  AND2_X1   g0792(.A1(new_n786), .A2(new_n992), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n744), .A2(new_n817), .B1(new_n741), .B2(new_n748), .ZN(new_n994));
  AOI211_X1 g0794(.A(new_n271), .B(new_n994), .C1(G283), .C2(new_n825), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n747), .A2(G294), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n754), .A2(G107), .B1(new_n756), .B2(G97), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT46), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n735), .B2(new_n581), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n995), .A2(new_n996), .A3(new_n997), .A4(new_n999), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n736), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n732), .B2(new_n740), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n754), .A2(G68), .B1(new_n756), .B2(new_n212), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n735), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n747), .A2(G159), .B1(new_n1004), .B2(G58), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n329), .B1(new_n745), .B2(G150), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(G50), .A2(new_n825), .B1(new_n811), .B2(G137), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n1003), .A2(new_n1005), .A3(new_n1006), .A4(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(G143), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n732), .A2(new_n1009), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n1000), .A2(new_n1002), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT47), .Z(new_n1012));
  OAI221_X1 g0812(.A(new_n993), .B1(new_n1012), .B2(new_n728), .C1(new_n789), .C2(new_n950), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n991), .A2(new_n1013), .ZN(G387));
  NAND2_X1  g0814(.A1(new_n985), .A2(new_n988), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n682), .B(KEYINPUT113), .Z(new_n1016));
  OAI211_X1 g0816(.A(new_n1015), .B(new_n1016), .C1(new_n717), .C2(new_n984), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n681), .A2(new_n780), .B1(G107), .B2(new_n237), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n246), .A2(new_n260), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT111), .ZN(new_n1020));
  AOI211_X1 g0820(.A(G45), .B(new_n680), .C1(G68), .C2(G77), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n320), .A2(new_n209), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n1022), .B(KEYINPUT50), .Z(new_n1023));
  AOI21_X1  g0823(.A(new_n778), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1018), .B1(new_n1020), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n786), .B1(new_n1025), .B2(new_n775), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n745), .A2(G317), .B1(new_n825), .B2(G303), .ZN(new_n1027));
  INV_X1    g0827(.A(G322), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1027), .B1(new_n740), .B2(new_n759), .C1(new_n732), .C2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT48), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n754), .A2(G283), .B1(new_n1004), .B2(G294), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT49), .ZN(new_n1035));
  OR2_X1    g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n755), .A2(new_n581), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n271), .B(new_n1038), .C1(G326), .C2(new_n811), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1036), .A2(new_n1037), .A3(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n731), .A2(G159), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n1041), .B(KEYINPUT112), .Z(new_n1042));
  OAI22_X1  g0842(.A1(new_n739), .A2(new_n214), .B1(new_n741), .B2(new_n828), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n329), .B(new_n1043), .C1(G50), .C2(new_n745), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n747), .A2(new_n320), .B1(new_n756), .B2(G97), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n753), .A2(new_n356), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(new_n212), .B2(new_n1004), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1042), .A2(new_n1044), .A3(new_n1045), .A4(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n728), .B1(new_n1040), .B2(new_n1048), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n1026), .B(new_n1049), .C1(new_n671), .C2(new_n773), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(new_n721), .B2(new_n984), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1017), .A2(new_n1051), .ZN(G393));
  AND2_X1   g0852(.A1(new_n989), .A2(new_n1016), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n976), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT115), .ZN(new_n1055));
  AND3_X1   g0855(.A1(new_n1015), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1055), .B1(new_n1015), .B2(new_n1054), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1053), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  AND2_X1   g0858(.A1(new_n254), .A2(new_n777), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n774), .B1(new_n457), .B2(new_n237), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n818), .A2(new_n748), .B1(new_n740), .B2(new_n744), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT52), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n759), .A2(new_n817), .B1(new_n816), .B2(new_n735), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n329), .B1(new_n741), .B2(new_n1028), .C1(new_n813), .C2(new_n739), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n753), .A2(new_n581), .ZN(new_n1065));
  NOR4_X1   g0865(.A1(new_n1063), .A2(new_n767), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(G150), .A2(new_n731), .B1(new_n745), .B2(G159), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(KEYINPUT114), .B(KEYINPUT51), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1067), .B(new_n1068), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n759), .A2(new_n209), .B1(new_n755), .B2(new_n501), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n271), .B1(new_n741), .B2(new_n1009), .C1(new_n359), .C2(new_n739), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n753), .A2(new_n303), .B1(new_n735), .B2(new_n396), .ZN(new_n1072));
  NOR3_X1   g0872(.A1(new_n1070), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n1062), .A2(new_n1066), .B1(new_n1069), .B2(new_n1073), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n786), .B1(new_n1059), .B2(new_n1060), .C1(new_n1074), .C2(new_n728), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(new_n938), .B2(new_n773), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n976), .B2(new_n721), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1058), .A2(new_n1077), .ZN(G390));
  NAND2_X1  g0878(.A1(new_n889), .A2(KEYINPUT101), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n879), .B1(new_n872), .B2(new_n867), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n897), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n892), .B1(new_n842), .B2(new_n846), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n716), .A2(KEYINPUT116), .A3(new_n795), .A4(new_n846), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n804), .A2(G330), .A3(new_n846), .A4(new_n795), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT116), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1085), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1082), .A2(new_n901), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1084), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  OAI211_X1 g0891(.A(G330), .B(new_n902), .C1(new_n907), .C2(new_n908), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1082), .B1(new_n890), .B2(new_n897), .ZN(new_n1094));
  AND2_X1   g0894(.A1(new_n1082), .A2(new_n901), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1093), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  AND2_X1   g0896(.A1(new_n1091), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1081), .A2(new_n771), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n786), .B1(new_n320), .B2(new_n808), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(KEYINPUT54), .B(G143), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n744), .A2(new_n821), .B1(new_n739), .B2(new_n1100), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n329), .B(new_n1101), .C1(G125), .C2(new_n811), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n735), .A2(new_n828), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT53), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n731), .A2(G128), .B1(new_n756), .B2(G50), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(G159), .A2(new_n754), .B1(new_n747), .B2(G137), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n1102), .A2(new_n1104), .A3(new_n1105), .A4(new_n1106), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n747), .A2(G107), .B1(new_n825), .B2(G97), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1108), .B1(new_n816), .B2(new_n818), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1109), .B(KEYINPUT118), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n329), .B1(new_n744), .B2(new_n581), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(G294), .B2(new_n811), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n754), .A2(G77), .B1(new_n756), .B2(G68), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n736), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1112), .B(new_n1113), .C1(new_n1114), .C2(new_n501), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1107), .B1(new_n1110), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1099), .B1(new_n1116), .B2(new_n727), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n1097), .A2(new_n721), .B1(new_n1098), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n842), .B1(new_n1085), .B2(new_n1088), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n915), .A2(G330), .A3(new_n795), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n846), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1119), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT117), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n804), .A2(G330), .A3(new_n795), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n1121), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1092), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1124), .B1(new_n1127), .B2(new_n842), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n842), .ZN(new_n1129));
  AOI211_X1 g0929(.A(KEYINPUT117), .B(new_n1129), .C1(new_n1092), .C2(new_n1126), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1123), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n691), .B1(new_n913), .B2(new_n914), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n430), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1133), .A2(new_n647), .A3(new_n838), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1097), .A2(new_n1131), .A3(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n1016), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1097), .B1(new_n1135), .B2(new_n1131), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1118), .B1(new_n1137), .B2(new_n1138), .ZN(G378));
  INV_X1    g0939(.A(new_n899), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n325), .A2(new_n652), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  AND2_X1   g0944(.A1(new_n348), .A2(new_n1144), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n348), .A2(new_n1144), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1142), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  AND2_X1   g0947(.A1(new_n345), .A2(new_n347), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1143), .B1(new_n1148), .B2(new_n340), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n348), .A2(new_n1144), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1149), .A2(new_n1150), .A3(new_n1141), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1147), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1152), .B1(new_n918), .B2(G330), .ZN(new_n1153));
  AND3_X1   g0953(.A1(new_n1147), .A2(KEYINPUT120), .A3(new_n1151), .ZN(new_n1154));
  AOI21_X1  g0954(.A(KEYINPUT120), .B1(new_n1147), .B2(new_n1151), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  AOI211_X1 g0956(.A(new_n691), .B(new_n1156), .C1(new_n910), .C2(new_n917), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1140), .B1(new_n1153), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1152), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n846), .A2(new_n795), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(new_n913), .B2(new_n914), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(KEYINPUT40), .A2(new_n909), .B1(new_n1161), .B2(new_n916), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1159), .B1(new_n1162), .B2(new_n691), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1156), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n918), .A2(G330), .A3(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1163), .A2(new_n1165), .A3(new_n899), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1158), .A2(new_n721), .A3(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n722), .B1(G50), .B2(new_n808), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n731), .A2(G125), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1169), .B1(new_n759), .B2(new_n821), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n745), .A2(G128), .B1(new_n825), .B2(G137), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n735), .B2(new_n1100), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1170), .B(new_n1172), .C1(G150), .C2(new_n754), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  OR2_X1    g0974(.A1(new_n1174), .A2(KEYINPUT59), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(KEYINPUT59), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n756), .A2(G159), .ZN(new_n1177));
  AOI211_X1 g0977(.A(G33), .B(G41), .C1(new_n811), .C2(G124), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .A4(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n329), .A2(new_n259), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n744), .A2(new_n350), .B1(new_n739), .B2(new_n356), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1180), .B(new_n1181), .C1(G283), .C2(new_n811), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n731), .A2(G116), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n747), .A2(G97), .B1(new_n756), .B2(G58), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n754), .A2(G68), .B1(new_n1004), .B2(new_n212), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .A4(new_n1185), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1186), .B(KEYINPUT119), .ZN(new_n1187));
  OR2_X1    g0987(.A1(new_n1187), .A2(KEYINPUT58), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1180), .B(new_n209), .C1(G33), .C2(G41), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1187), .A2(KEYINPUT58), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1179), .A2(new_n1188), .A3(new_n1189), .A4(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1168), .B1(new_n1191), .B2(new_n727), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n1164), .B2(new_n772), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1167), .A2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  AND3_X1   g0995(.A1(new_n1163), .A2(new_n899), .A3(new_n1165), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n899), .B1(new_n1163), .B2(new_n1165), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1131), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1091), .A2(new_n1096), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1135), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(KEYINPUT57), .B1(new_n1198), .B2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1158), .A2(KEYINPUT57), .A3(new_n1166), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1134), .B1(new_n1097), .B2(new_n1131), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1016), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1195), .B1(new_n1202), .B2(new_n1205), .ZN(G375));
  NAND2_X1  g1006(.A1(new_n1131), .A2(new_n1135), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n965), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1123), .B(new_n1134), .C1(new_n1128), .C2(new_n1130), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n786), .B1(G68), .B2(new_n808), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n846), .A2(new_n772), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n744), .A2(new_n827), .B1(new_n739), .B2(new_n828), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n329), .B(new_n1213), .C1(G128), .C2(new_n811), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n736), .A2(G159), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n754), .A2(G50), .B1(new_n756), .B2(G58), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1100), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(G132), .A2(new_n731), .B1(new_n747), .B2(new_n1217), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .A4(new_n1218), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n747), .A2(G116), .B1(new_n825), .B2(G107), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n813), .B2(new_n818), .ZN(new_n1221));
  XOR2_X1   g1021(.A(new_n1221), .B(KEYINPUT121), .Z(new_n1222));
  OAI21_X1  g1022(.A(new_n329), .B1(new_n744), .B2(new_n816), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n1046), .B(new_n1223), .C1(G77), .C2(new_n756), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1222), .A2(new_n1224), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n736), .A2(G97), .B1(G303), .B2(new_n811), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(new_n1226), .B(KEYINPUT122), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1219), .B1(new_n1225), .B2(new_n1227), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n1211), .B(new_n1212), .C1(new_n727), .C2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(new_n1131), .B2(new_n721), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1210), .A2(new_n1230), .ZN(G381));
  INV_X1    g1031(.A(KEYINPUT123), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(G375), .B(new_n1232), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n991), .A2(new_n1058), .A3(new_n1013), .A4(new_n1077), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1017), .A2(new_n1051), .A3(new_n791), .ZN(new_n1235));
  OR2_X1    g1035(.A1(new_n1235), .A2(G384), .ZN(new_n1236));
  NOR4_X1   g1036(.A1(G378), .A2(new_n1234), .A3(G381), .A4(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1233), .A2(new_n1237), .ZN(G407));
  INV_X1    g1038(.A(G378), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n653), .A2(G213), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1239), .A2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1233), .A2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(G407), .A2(new_n1244), .A3(G213), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT124), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(G407), .A2(new_n1244), .A3(KEYINPUT124), .A4(G213), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(G409));
  NAND2_X1  g1049(.A1(new_n1241), .A2(G2897), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1016), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(new_n1131), .B2(new_n1135), .ZN(new_n1252));
  AND2_X1   g1052(.A1(new_n1209), .A2(KEYINPUT60), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1209), .A2(KEYINPUT60), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1252), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n807), .A2(KEYINPUT125), .A3(new_n835), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1230), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT125), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(G384), .A2(new_n1259), .ZN(new_n1260));
  AND3_X1   g1060(.A1(new_n1255), .A2(new_n1258), .A3(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1260), .B1(new_n1255), .B2(new_n1258), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1250), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1260), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1207), .A2(new_n1016), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1254), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1209), .A2(KEYINPUT60), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1265), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1264), .B1(new_n1268), .B2(new_n1257), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1255), .A2(new_n1258), .A3(new_n1260), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1250), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1269), .A2(new_n1270), .A3(new_n1271), .ZN(new_n1272));
  AND2_X1   g1072(.A1(new_n1263), .A2(new_n1272), .ZN(new_n1273));
  OAI211_X1 g1073(.A(G378), .B(new_n1195), .C1(new_n1202), .C2(new_n1205), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1207), .A2(new_n1200), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1275), .A2(new_n1016), .A3(new_n1136), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1158), .A2(new_n1166), .ZN(new_n1277));
  NOR3_X1   g1077(.A1(new_n1277), .A2(new_n1204), .A3(new_n965), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n1276), .B(new_n1118), .C1(new_n1278), .C2(new_n1194), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1241), .B1(new_n1274), .B2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(KEYINPUT61), .B1(new_n1273), .B2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(G393), .A2(G396), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n1235), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT126), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1234), .A2(new_n1286), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(new_n991), .A2(new_n1013), .B1(new_n1058), .B2(new_n1077), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1285), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1288), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1290), .A2(new_n1284), .A3(new_n1286), .A4(new_n1234), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1289), .A2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1280), .A2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT63), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1292), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1280), .A2(KEYINPUT63), .A3(new_n1293), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1282), .A2(new_n1296), .A3(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT61), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1263), .A2(new_n1272), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1299), .B1(new_n1300), .B2(new_n1280), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT62), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1274), .A2(new_n1279), .ZN(new_n1303));
  AND4_X1   g1103(.A1(new_n1302), .A2(new_n1303), .A3(new_n1240), .A4(new_n1293), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1302), .B1(new_n1280), .B2(new_n1293), .ZN(new_n1305));
  NOR3_X1   g1105(.A1(new_n1301), .A2(new_n1304), .A3(new_n1305), .ZN(new_n1306));
  AND2_X1   g1106(.A1(new_n1289), .A2(new_n1291), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1298), .B1(new_n1306), .B2(new_n1307), .ZN(G405));
  NAND2_X1  g1108(.A1(G375), .A2(new_n1239), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT127), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1309), .A2(new_n1310), .A3(new_n1274), .ZN(new_n1311));
  AND2_X1   g1111(.A1(new_n1311), .A2(new_n1293), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1274), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1198), .A2(new_n1201), .A3(KEYINPUT57), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT57), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1315), .B1(new_n1277), .B2(new_n1204), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1314), .A2(new_n1316), .A3(new_n1016), .ZN(new_n1317));
  AOI21_X1  g1117(.A(G378), .B1(new_n1317), .B2(new_n1195), .ZN(new_n1318));
  OAI21_X1  g1118(.A(KEYINPUT127), .B1(new_n1313), .B2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1319), .A2(new_n1307), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1309), .A2(new_n1274), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1292), .A2(new_n1321), .A3(KEYINPUT127), .ZN(new_n1322));
  AND3_X1   g1122(.A1(new_n1312), .A2(new_n1320), .A3(new_n1322), .ZN(new_n1323));
  AOI22_X1  g1123(.A1(new_n1320), .A2(new_n1322), .B1(new_n1293), .B2(new_n1311), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1323), .A2(new_n1324), .ZN(G402));
endmodule


