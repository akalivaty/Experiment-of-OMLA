//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 1 1 1 0 0 0 0 0 0 0 0 0 1 1 1 0 1 1 0 1 0 1 0 1 0 0 0 0 0 0 1 0 1 1 1 1 0 0 1 0 1 0 0 0 0 1 1 0 1 1 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:53 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1212,
    new_n1213, new_n1214, new_n1216, new_n1217, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  INV_X1    g0006(.A(G226), .ZN(new_n207));
  INV_X1    g0007(.A(G116), .ZN(new_n208));
  INV_X1    g0008(.A(G270), .ZN(new_n209));
  OAI22_X1  g0009(.A1(new_n202), .A2(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  AOI21_X1  g0010(.A(new_n210), .B1(G58), .B2(G232), .ZN(new_n211));
  XNOR2_X1  g0011(.A(KEYINPUT64), .B(G244), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n212), .A2(G77), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G87), .A2(G250), .ZN(new_n215));
  NAND4_X1  g0015(.A1(new_n211), .A2(new_n213), .A3(new_n214), .A4(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G68), .ZN(new_n217));
  INV_X1    g0017(.A(G238), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n206), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT1), .Z(new_n221));
  NOR2_X1   g0021(.A1(new_n206), .A2(G13), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n222), .B(G250), .C1(G257), .C2(G264), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT0), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(G50), .B1(G58), .B2(G68), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n221), .B(new_n224), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT2), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(new_n207), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT65), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G264), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(new_n209), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n236), .B(new_n240), .ZN(G358));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G107), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(new_n208), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  XNOR2_X1  g0048(.A(KEYINPUT3), .B(G33), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n249), .A2(G223), .A3(G1698), .ZN(new_n250));
  INV_X1    g0050(.A(G77), .ZN(new_n251));
  INV_X1    g0051(.A(G222), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT3), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G33), .ZN(new_n256));
  AND2_X1   g0056(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n257));
  NOR2_X1   g0057(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n258));
  OAI211_X1 g0058(.A(new_n254), .B(new_n256), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  OAI221_X1 g0059(.A(new_n250), .B1(new_n251), .B2(new_n249), .C1(new_n252), .C2(new_n259), .ZN(new_n260));
  AND2_X1   g0060(.A1(G33), .A2(G41), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT69), .ZN(new_n262));
  NOR3_X1   g0062(.A1(new_n261), .A2(new_n262), .A3(new_n225), .ZN(new_n263));
  AND2_X1   g0063(.A1(G1), .A2(G13), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G33), .A2(G41), .ZN(new_n265));
  AOI21_X1  g0065(.A(KEYINPUT69), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  OR2_X1    g0066(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n260), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G1), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n269), .B(G274), .C1(G41), .C2(G45), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n269), .B1(G41), .B2(G45), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n271), .B1(new_n225), .B2(new_n261), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(KEYINPUT67), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n264), .A2(new_n265), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT67), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n274), .A2(new_n275), .A3(new_n271), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT66), .B(G226), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n273), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n268), .A2(new_n270), .A3(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G190), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n279), .A2(G200), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n203), .A2(G20), .ZN(new_n283));
  INV_X1    g0083(.A(G150), .ZN(new_n284));
  NOR2_X1   g0084(.A1(G20), .A2(G33), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n226), .A2(G33), .ZN(new_n287));
  OR2_X1    g0087(.A1(KEYINPUT8), .A2(G58), .ZN(new_n288));
  NAND2_X1  g0088(.A1(KEYINPUT8), .A2(G58), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OAI221_X1 g0090(.A(new_n283), .B1(new_n284), .B2(new_n286), .C1(new_n287), .C2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n225), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  AND2_X1   g0094(.A1(new_n292), .A2(new_n225), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n295), .B1(G1), .B2(new_n226), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G50), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT70), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n269), .A2(G13), .A3(G20), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(new_n202), .ZN(new_n300));
  AND3_X1   g0100(.A1(new_n297), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n298), .B1(new_n297), .B2(new_n300), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n294), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(KEYINPUT74), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT74), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n305), .B(new_n294), .C1(new_n301), .C2(new_n302), .ZN(new_n306));
  AND3_X1   g0106(.A1(new_n304), .A2(KEYINPUT9), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(KEYINPUT9), .B1(new_n304), .B2(new_n306), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n281), .B(new_n282), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(KEYINPUT10), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n304), .A2(new_n306), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT9), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n304), .A2(KEYINPUT9), .A3(new_n306), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT10), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n315), .A2(new_n316), .A3(new_n281), .A4(new_n282), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n310), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G179), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n280), .A2(new_n320), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n321), .B(new_n303), .C1(G169), .C2(new_n280), .ZN(new_n322));
  XNOR2_X1  g0122(.A(new_n322), .B(KEYINPUT71), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT18), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n290), .A2(new_n299), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n293), .B1(new_n269), .B2(G20), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n325), .B1(new_n326), .B2(new_n290), .ZN(new_n327));
  XNOR2_X1  g0127(.A(new_n327), .B(KEYINPUT81), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT7), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n329), .B1(new_n249), .B2(G20), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n254), .A2(new_n256), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n329), .A2(G20), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n217), .B1(new_n330), .B2(new_n333), .ZN(new_n334));
  AND2_X1   g0134(.A1(G58), .A2(G68), .ZN(new_n335));
  OAI21_X1  g0135(.A(G20), .B1(new_n335), .B2(new_n201), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(KEYINPUT78), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n285), .A2(G159), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT78), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n339), .B(G20), .C1(new_n335), .C2(new_n201), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n337), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(KEYINPUT79), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT79), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n337), .A2(new_n343), .A3(new_n338), .A4(new_n340), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n334), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n295), .B1(new_n345), .B2(KEYINPUT16), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT16), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n331), .A2(new_n226), .ZN(new_n348));
  OAI21_X1  g0148(.A(KEYINPUT80), .B1(new_n253), .B2(KEYINPUT3), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT80), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n350), .A2(new_n255), .A3(G33), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n349), .A2(new_n351), .A3(new_n254), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n348), .A2(new_n329), .B1(new_n352), .B2(new_n332), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n353), .A2(new_n217), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n347), .B1(new_n354), .B2(new_n341), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n328), .B1(new_n346), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(G169), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n254), .A2(new_n256), .A3(G226), .A4(G1698), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT82), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n249), .A2(KEYINPUT82), .A3(G226), .A4(G1698), .ZN(new_n361));
  OR2_X1    g0161(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n362));
  NAND2_X1  g0162(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n364), .A2(new_n249), .A3(G223), .ZN(new_n365));
  NAND2_X1  g0165(.A1(G33), .A2(G87), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n360), .A2(new_n361), .A3(new_n365), .A4(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n267), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n270), .B1(new_n272), .B2(new_n233), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT83), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OAI211_X1 g0171(.A(KEYINPUT83), .B(new_n270), .C1(new_n272), .C2(new_n233), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n357), .B1(new_n368), .B2(new_n373), .ZN(new_n374));
  AOI22_X1  g0174(.A1(new_n267), .A2(new_n367), .B1(new_n371), .B2(new_n372), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n374), .B1(G179), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n324), .B1(new_n356), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n342), .A2(new_n344), .ZN(new_n378));
  INV_X1    g0178(.A(new_n334), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n378), .A2(KEYINPUT16), .A3(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n380), .A2(new_n293), .A3(new_n355), .ZN(new_n381));
  INV_X1    g0181(.A(new_n328), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n375), .A2(G179), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n384), .B1(new_n357), .B2(new_n375), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n383), .A2(KEYINPUT18), .A3(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(G190), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n368), .A2(new_n373), .A3(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(new_n375), .B2(G200), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n381), .A2(new_n382), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(KEYINPUT17), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT17), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n356), .A2(new_n392), .A3(new_n389), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n377), .A2(new_n386), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  OR2_X1    g0194(.A1(KEYINPUT15), .A2(G87), .ZN(new_n395));
  NAND2_X1  g0195(.A1(KEYINPUT15), .A2(G87), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n395), .A2(new_n226), .A3(G33), .A4(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n288), .A2(new_n285), .A3(new_n289), .ZN(new_n398));
  NAND2_X1  g0198(.A1(G20), .A2(G77), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n397), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n293), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n299), .A2(G77), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n326), .A2(G77), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n401), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT72), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n402), .B1(new_n400), .B2(new_n293), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT72), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n407), .A2(new_n408), .A3(new_n404), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n406), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n249), .A2(G238), .A3(G1698), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n331), .A2(G107), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n411), .B(new_n412), .C1(new_n233), .C2(new_n259), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n267), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n273), .A2(new_n212), .A3(new_n276), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n414), .A2(new_n270), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n410), .B1(G200), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n417), .B1(new_n387), .B2(new_n416), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT73), .ZN(new_n419));
  AND4_X1   g0219(.A1(new_n408), .A2(new_n401), .A3(new_n403), .A4(new_n404), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n408), .B1(new_n407), .B2(new_n404), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n270), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n423), .B1(new_n413), .B2(new_n267), .ZN(new_n424));
  AOI21_X1  g0224(.A(G169), .B1(new_n424), .B2(new_n415), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n419), .B1(new_n422), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n424), .A2(new_n320), .A3(new_n415), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n416), .A2(new_n357), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n428), .A2(new_n410), .A3(KEYINPUT73), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n426), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n323), .A2(new_n394), .A3(new_n418), .A4(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n273), .A2(G238), .A3(new_n276), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n270), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n263), .A2(new_n266), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n207), .B1(new_n362), .B2(new_n363), .ZN(new_n435));
  NAND2_X1  g0235(.A1(G232), .A2(G1698), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n249), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(G33), .A2(G97), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n434), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT13), .B1(new_n433), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(G226), .B1(new_n257), .B2(new_n258), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n331), .B1(new_n442), .B2(new_n436), .ZN(new_n443));
  INV_X1    g0243(.A(new_n439), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n267), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT13), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n445), .A2(new_n446), .A3(new_n270), .A4(new_n432), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n441), .A2(G190), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT76), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n441), .A2(KEYINPUT76), .A3(new_n447), .A4(G190), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n217), .A2(G20), .ZN(new_n453));
  INV_X1    g0253(.A(G13), .ZN(new_n454));
  NOR3_X1   g0254(.A1(new_n453), .A2(G1), .A3(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n455), .A2(KEYINPUT77), .ZN(new_n456));
  XOR2_X1   g0256(.A(new_n456), .B(KEYINPUT12), .Z(new_n457));
  OAI221_X1 g0257(.A(new_n453), .B1(new_n287), .B2(new_n251), .C1(new_n286), .C2(new_n202), .ZN(new_n458));
  AOI21_X1  g0258(.A(KEYINPUT11), .B1(new_n458), .B2(new_n293), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n458), .A2(KEYINPUT11), .A3(new_n293), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n460), .B1(new_n217), .B2(new_n296), .ZN(new_n461));
  NOR3_X1   g0261(.A1(new_n457), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT75), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n441), .A2(new_n463), .A3(new_n447), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n433), .A2(new_n440), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n465), .A2(KEYINPUT75), .A3(new_n446), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n464), .A2(G200), .A3(new_n466), .ZN(new_n467));
  AND3_X1   g0267(.A1(new_n452), .A2(new_n462), .A3(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n462), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n464), .A2(G169), .A3(new_n466), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(KEYINPUT14), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n441), .A2(G179), .A3(new_n447), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT14), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n464), .A2(new_n466), .A3(new_n473), .A4(G169), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n471), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n468), .B1(new_n469), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NOR3_X1   g0277(.A1(new_n319), .A2(new_n431), .A3(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  XNOR2_X1  g0279(.A(KEYINPUT88), .B(KEYINPUT24), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n254), .A2(new_n256), .A3(new_n226), .A4(G87), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT22), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT22), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n249), .A2(new_n483), .A3(new_n226), .A4(G87), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n253), .A2(new_n208), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n226), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n226), .A2(G107), .ZN(new_n488));
  XNOR2_X1  g0288(.A(new_n488), .B(KEYINPUT23), .ZN(new_n489));
  AND4_X1   g0289(.A1(new_n480), .A2(new_n485), .A3(new_n487), .A4(new_n489), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n482), .A2(new_n484), .B1(new_n226), .B2(new_n486), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n480), .B1(new_n491), .B2(new_n489), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n293), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n269), .A2(G33), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n299), .A2(new_n494), .A3(new_n225), .A4(new_n292), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G107), .ZN(new_n497));
  INV_X1    g0297(.A(new_n299), .ZN(new_n498));
  INV_X1    g0298(.A(G107), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n498), .B(new_n499), .C1(KEYINPUT89), .C2(KEYINPUT25), .ZN(new_n500));
  NAND2_X1  g0300(.A1(KEYINPUT89), .A2(KEYINPUT25), .ZN(new_n501));
  XNOR2_X1  g0301(.A(new_n500), .B(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n493), .A2(new_n497), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(G33), .A2(G294), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n254), .A2(new_n256), .A3(G257), .A4(G1698), .ZN(new_n505));
  INV_X1    g0305(.A(G250), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n504), .B(new_n505), .C1(new_n259), .C2(new_n506), .ZN(new_n507));
  XNOR2_X1  g0307(.A(KEYINPUT5), .B(G41), .ZN(new_n508));
  INV_X1    g0308(.A(G45), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n509), .A2(G1), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n508), .A2(new_n510), .B1(new_n264), .B2(new_n265), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n507), .A2(new_n267), .B1(G264), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n508), .A2(G274), .A3(new_n510), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n357), .ZN(new_n515));
  INV_X1    g0315(.A(new_n514), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n320), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n503), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n495), .A2(new_n208), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n269), .A2(new_n208), .A3(G13), .A4(G20), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n292), .A2(new_n225), .B1(G20), .B2(new_n208), .ZN(new_n522));
  NAND2_X1  g0322(.A1(G33), .A2(G283), .ZN(new_n523));
  INV_X1    g0323(.A(G97), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n523), .B(new_n226), .C1(G33), .C2(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(KEYINPUT20), .B1(new_n522), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n522), .A2(KEYINPUT20), .A3(new_n525), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n520), .B(new_n521), .C1(new_n526), .C2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  XNOR2_X1  g0330(.A(KEYINPUT87), .B(G303), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n331), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n254), .A2(new_n256), .A3(G264), .A4(G1698), .ZN(new_n533));
  INV_X1    g0333(.A(G257), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n532), .B(new_n533), .C1(new_n534), .C2(new_n259), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n267), .ZN(new_n536));
  AND2_X1   g0336(.A1(KEYINPUT5), .A2(G41), .ZN(new_n537));
  NOR2_X1   g0337(.A1(KEYINPUT5), .A2(G41), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n510), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n539), .A2(G270), .A3(new_n274), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n536), .A2(new_n513), .A3(new_n541), .ZN(new_n542));
  NOR3_X1   g0342(.A1(new_n530), .A2(new_n542), .A3(new_n320), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n522), .A2(new_n525), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT20), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n519), .B1(new_n546), .B2(new_n527), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n357), .B1(new_n547), .B2(new_n521), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n542), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(KEYINPUT21), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT21), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n548), .A2(new_n551), .A3(new_n542), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n543), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n536), .A2(G190), .A3(new_n513), .A4(new_n541), .ZN(new_n554));
  INV_X1    g0354(.A(new_n513), .ZN(new_n555));
  AOI211_X1 g0355(.A(new_n555), .B(new_n540), .C1(new_n535), .C2(new_n267), .ZN(new_n556));
  INV_X1    g0356(.A(G200), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n530), .B(new_n554), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n518), .A2(new_n553), .A3(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(new_n486), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n254), .A2(new_n256), .A3(G244), .A4(G1698), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n560), .B(new_n561), .C1(new_n259), .C2(new_n218), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n267), .ZN(new_n563));
  OAI221_X1 g0363(.A(G250), .B1(G1), .B2(new_n509), .C1(new_n261), .C2(new_n225), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n510), .A2(G274), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n557), .B1(new_n563), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n226), .ZN(new_n570));
  INV_X1    g0370(.A(G87), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n571), .A2(new_n524), .A3(new_n499), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n226), .A2(G33), .A3(G97), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT19), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n570), .A2(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n254), .A2(new_n256), .A3(new_n226), .A4(G68), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n293), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n395), .A2(new_n396), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n498), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n495), .A2(new_n571), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n578), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  OAI21_X1  g0383(.A(KEYINPUT86), .B1(new_n568), .B2(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n566), .B1(new_n562), .B2(new_n267), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(G190), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n295), .B1(new_n575), .B2(new_n576), .ZN(new_n587));
  INV_X1    g0387(.A(new_n580), .ZN(new_n588));
  NOR3_X1   g0388(.A1(new_n587), .A2(new_n588), .A3(new_n581), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT86), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n589), .B(new_n590), .C1(new_n557), .C2(new_n585), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n584), .A2(new_n586), .A3(new_n591), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n578), .B(new_n580), .C1(new_n579), .C2(new_n495), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n585), .A2(G179), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n585), .A2(new_n357), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n593), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  AND2_X1   g0397(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n512), .A2(new_n387), .A3(new_n513), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(KEYINPUT90), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n514), .A2(new_n557), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT90), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n512), .A2(new_n602), .A3(new_n387), .A4(new_n513), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n600), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n485), .A2(new_n487), .A3(new_n489), .ZN(new_n605));
  INV_X1    g0405(.A(new_n480), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n491), .A2(new_n480), .A3(new_n489), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n609), .A2(new_n293), .B1(G107), .B2(new_n496), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n604), .A2(new_n610), .A3(new_n502), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT4), .ZN(new_n612));
  INV_X1    g0412(.A(G244), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n612), .B1(new_n259), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n249), .A2(G250), .A3(G1698), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n364), .A2(new_n249), .A3(KEYINPUT4), .A4(G244), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n614), .A2(new_n523), .A3(new_n615), .A4(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n267), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT85), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n539), .A2(new_n274), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n619), .B1(new_n620), .B2(new_n534), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n511), .A2(KEYINPUT85), .A3(G257), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n555), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n618), .A2(new_n623), .A3(new_n320), .ZN(new_n624));
  AOI21_X1  g0424(.A(G169), .B1(new_n618), .B2(new_n623), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT84), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n627), .B1(new_n353), .B2(new_n499), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n499), .A2(KEYINPUT6), .A3(G97), .ZN(new_n629));
  XOR2_X1   g0429(.A(G97), .B(G107), .Z(new_n630));
  OAI21_X1  g0430(.A(new_n629), .B1(new_n630), .B2(KEYINPUT6), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n631), .A2(G20), .B1(G77), .B2(new_n285), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n352), .A2(new_n332), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n330), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n634), .A2(KEYINPUT84), .A3(G107), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n628), .A2(new_n632), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n293), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n299), .A2(G97), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n638), .B1(new_n496), .B2(G97), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n626), .A2(new_n640), .ZN(new_n641));
  AND3_X1   g0441(.A1(new_n618), .A2(new_n623), .A3(new_n387), .ZN(new_n642));
  AOI21_X1  g0442(.A(G200), .B1(new_n618), .B2(new_n623), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n637), .B(new_n639), .C1(new_n642), .C2(new_n643), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n598), .A2(new_n611), .A3(new_n641), .A4(new_n644), .ZN(new_n645));
  NOR3_X1   g0445(.A1(new_n479), .A2(new_n559), .A3(new_n645), .ZN(G372));
  NAND2_X1  g0446(.A1(new_n391), .A2(new_n393), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n452), .A2(new_n462), .A3(new_n467), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT93), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n430), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n426), .A2(new_n429), .A3(KEYINPUT93), .A4(new_n427), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n475), .A2(new_n469), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n649), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n377), .A2(new_n386), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n318), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n659), .A2(new_n323), .ZN(new_n660));
  OAI21_X1  g0460(.A(KEYINPUT91), .B1(new_n595), .B2(new_n596), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT91), .ZN(new_n662));
  OAI211_X1 g0462(.A(new_n594), .B(new_n662), .C1(new_n357), .C2(new_n585), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n593), .ZN(new_n665));
  OAI211_X1 g0465(.A(new_n586), .B(new_n589), .C1(new_n557), .C2(new_n585), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n611), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n518), .A2(new_n553), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n669), .A2(new_n641), .A3(new_n644), .A4(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n598), .A2(new_n640), .A3(new_n626), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(KEYINPUT26), .ZN(new_n673));
  INV_X1    g0473(.A(new_n667), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT26), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n641), .A2(KEYINPUT92), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n641), .A2(KEYINPUT92), .ZN(new_n677));
  OAI211_X1 g0477(.A(new_n674), .B(new_n675), .C1(new_n676), .C2(new_n677), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n671), .A2(new_n673), .A3(new_n678), .A4(new_n665), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n478), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n660), .A2(new_n680), .ZN(G369));
  NOR2_X1   g0481(.A1(new_n454), .A2(G20), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(new_n269), .ZN(new_n683));
  XOR2_X1   g0483(.A(new_n683), .B(KEYINPUT94), .Z(new_n684));
  OR2_X1    g0484(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(new_n686), .A3(G213), .ZN(new_n687));
  INV_X1    g0487(.A(G343), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n503), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n518), .B1(new_n668), .B2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n515), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n692), .B1(new_n610), .B2(new_n502), .ZN(new_n693));
  INV_X1    g0493(.A(new_n689), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n693), .A2(new_n517), .A3(new_n694), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n553), .A2(new_n689), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(new_n695), .ZN(new_n699));
  INV_X1    g0499(.A(new_n696), .ZN(new_n700));
  INV_X1    g0500(.A(new_n553), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n694), .A2(new_n530), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n556), .A2(G179), .A3(new_n529), .ZN(new_n704));
  AND3_X1   g0504(.A1(new_n548), .A2(new_n551), .A3(new_n542), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n551), .B1(new_n548), .B2(new_n542), .ZN(new_n706));
  OAI211_X1 g0506(.A(new_n558), .B(new_n704), .C1(new_n705), .C2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n703), .B1(new_n707), .B2(new_n702), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(G330), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n700), .A2(new_n709), .ZN(new_n710));
  OR2_X1    g0510(.A1(new_n699), .A2(new_n710), .ZN(G399));
  NOR2_X1   g0511(.A1(new_n572), .A2(G116), .ZN(new_n712));
  INV_X1    g0512(.A(G41), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n222), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n712), .A2(new_n714), .A3(G1), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n715), .B1(new_n229), .B2(new_n714), .ZN(new_n716));
  XOR2_X1   g0516(.A(KEYINPUT95), .B(KEYINPUT28), .Z(new_n717));
  XNOR2_X1  g0517(.A(new_n716), .B(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n641), .A2(new_n644), .ZN(new_n719));
  XNOR2_X1  g0519(.A(new_n719), .B(KEYINPUT97), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n669), .A2(new_n670), .ZN(new_n722));
  OAI21_X1  g0522(.A(KEYINPUT98), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  OR2_X1    g0523(.A1(new_n672), .A2(KEYINPUT26), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT98), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n720), .A2(new_n725), .A3(new_n670), .A4(new_n669), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n674), .B1(new_n676), .B2(new_n677), .ZN(new_n727));
  AOI22_X1  g0527(.A1(new_n727), .A2(KEYINPUT26), .B1(new_n593), .B2(new_n664), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n723), .A2(new_n724), .A3(new_n726), .A4(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n729), .A2(KEYINPUT29), .A3(new_n694), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n679), .A2(new_n694), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT29), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  AOI22_X1  g0534(.A1(new_n618), .A2(new_n623), .B1(new_n512), .B2(new_n513), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n563), .A2(new_n567), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n735), .A2(new_n320), .A3(new_n542), .A4(new_n736), .ZN(new_n737));
  AND2_X1   g0537(.A1(new_n618), .A2(new_n623), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n540), .B1(new_n535), .B2(new_n267), .ZN(new_n739));
  AND3_X1   g0539(.A1(new_n739), .A2(G179), .A3(new_n585), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n738), .A2(new_n740), .A3(KEYINPUT30), .A4(new_n516), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT30), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n618), .A2(new_n623), .A3(new_n512), .A4(new_n513), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n739), .A2(G179), .A3(new_n585), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n742), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n737), .A2(new_n741), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(new_n689), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n645), .A2(new_n559), .A3(new_n689), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT31), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n746), .A2(KEYINPUT31), .A3(new_n689), .ZN(new_n751));
  XOR2_X1   g0551(.A(new_n751), .B(KEYINPUT96), .Z(new_n752));
  NAND2_X1  g0552(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G330), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n734), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n755), .B(KEYINPUT99), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n718), .B1(new_n756), .B2(G1), .ZN(G364));
  NOR3_X1   g0557(.A1(new_n387), .A2(G179), .A3(G200), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n226), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(G97), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n226), .A2(G179), .ZN(new_n762));
  NOR2_X1   g0562(.A1(G190), .A2(G200), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G159), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n226), .A2(new_n320), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR3_X1   g0568(.A1(new_n768), .A2(new_n557), .A3(G190), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  OAI221_X1 g0570(.A(new_n761), .B1(new_n766), .B2(KEYINPUT32), .C1(new_n770), .C2(new_n217), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n771), .B1(KEYINPUT32), .B2(new_n766), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n767), .A2(new_n763), .ZN(new_n773));
  NOR3_X1   g0573(.A1(new_n768), .A2(new_n387), .A3(G200), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(G58), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n249), .B1(new_n251), .B2(new_n773), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n762), .A2(new_n387), .A3(G200), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT102), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n777), .B1(G107), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n387), .A2(new_n557), .ZN(new_n782));
  INV_X1    g0582(.A(KEYINPUT101), .ZN(new_n783));
  AND3_X1   g0583(.A1(new_n767), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n783), .B1(new_n767), .B2(new_n782), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G50), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n782), .A2(new_n762), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G87), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n772), .A2(new_n781), .A3(new_n788), .A4(new_n791), .ZN(new_n792));
  XOR2_X1   g0592(.A(KEYINPUT33), .B(G317), .Z(new_n793));
  INV_X1    g0593(.A(G322), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n770), .A2(new_n793), .B1(new_n775), .B2(new_n794), .ZN(new_n795));
  XOR2_X1   g0595(.A(new_n795), .B(KEYINPUT103), .Z(new_n796));
  NAND2_X1  g0596(.A1(new_n787), .A2(G326), .ZN(new_n797));
  INV_X1    g0597(.A(G294), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n759), .A2(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n249), .B1(new_n790), .B2(G303), .ZN(new_n800));
  INV_X1    g0600(.A(G329), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n800), .B1(new_n801), .B2(new_n764), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n799), .B(new_n802), .C1(G283), .C2(new_n780), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n796), .A2(new_n797), .A3(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(G311), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n773), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n792), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n225), .B1(G20), .B2(new_n357), .ZN(new_n808));
  NOR2_X1   g0608(.A1(G13), .A2(G33), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n810), .A2(G20), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(new_n808), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n331), .A2(new_n222), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n813), .B(KEYINPUT100), .Z(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n815), .B1(new_n244), .B2(G45), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n816), .B1(G45), .B2(new_n229), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n249), .A2(G355), .A3(new_n222), .ZN(new_n818));
  OAI211_X1 g0618(.A(new_n817), .B(new_n818), .C1(G116), .C2(new_n222), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n807), .A2(new_n808), .B1(new_n812), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n269), .B1(new_n682), .B2(G45), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n714), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n811), .ZN(new_n825));
  OAI211_X1 g0625(.A(new_n820), .B(new_n824), .C1(new_n708), .C2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n824), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n709), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n708), .A2(G330), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n826), .B1(new_n828), .B2(new_n829), .ZN(G396));
  NOR2_X1   g0630(.A1(new_n694), .A2(new_n422), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n653), .A2(new_n831), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n418), .B(new_n430), .C1(new_n422), .C2(new_n694), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n731), .B(new_n834), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(new_n754), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(new_n827), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n779), .A2(new_n217), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n249), .B1(new_n789), .B2(new_n202), .C1(new_n759), .C2(new_n776), .ZN(new_n839));
  INV_X1    g0639(.A(new_n773), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n769), .A2(G150), .B1(G159), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(G143), .ZN(new_n842));
  INV_X1    g0642(.A(G137), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n841), .B1(new_n842), .B2(new_n775), .C1(new_n786), .C2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT34), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n838), .B(new_n839), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(G132), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n846), .B1(new_n845), .B2(new_n844), .C1(new_n847), .C2(new_n764), .ZN(new_n848));
  INV_X1    g0648(.A(G283), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n761), .B1(new_n770), .B2(new_n849), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n775), .A2(new_n798), .B1(new_n773), .B2(new_n208), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n850), .B(new_n851), .C1(G87), .C2(new_n780), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n787), .A2(G303), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n852), .B(new_n853), .C1(new_n805), .C2(new_n764), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n331), .B1(new_n789), .B2(new_n499), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT105), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n848), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n808), .A2(new_n809), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n858), .B(KEYINPUT104), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n857), .A2(new_n808), .B1(new_n251), .B2(new_n859), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n860), .B(new_n824), .C1(new_n834), .C2(new_n810), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n837), .A2(new_n861), .ZN(G384));
  NOR2_X1   g0662(.A1(new_n655), .A2(new_n689), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n657), .A2(new_n647), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n346), .B1(KEYINPUT16), .B2(new_n345), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n687), .B1(new_n865), .B2(new_n382), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  AOI22_X1  g0667(.A1(new_n865), .A2(new_n382), .B1(new_n376), .B2(new_n687), .ZN(new_n868));
  AND3_X1   g0668(.A1(new_n381), .A2(new_n382), .A3(new_n389), .ZN(new_n869));
  OAI21_X1  g0669(.A(KEYINPUT37), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n687), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n383), .B1(new_n385), .B2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT37), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n872), .A2(new_n873), .A3(new_n390), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n870), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n867), .A2(KEYINPUT107), .A3(KEYINPUT38), .A4(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n867), .A2(KEYINPUT38), .A3(new_n875), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n383), .A2(new_n871), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n376), .A2(new_n687), .B1(new_n381), .B2(new_n382), .ZN(new_n880));
  NOR3_X1   g0680(.A1(new_n880), .A2(new_n869), .A3(KEYINPUT37), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n873), .B1(new_n872), .B2(new_n390), .ZN(new_n882));
  OAI22_X1  g0682(.A1(new_n394), .A2(new_n879), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT38), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT107), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n877), .B1(new_n878), .B2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n886), .A2(KEYINPUT39), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n380), .A2(new_n293), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n345), .A2(KEYINPUT16), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OAI22_X1  g0690(.A1(new_n890), .A2(new_n328), .B1(new_n385), .B2(new_n871), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n873), .B1(new_n891), .B2(new_n390), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n892), .A2(new_n881), .ZN(new_n893));
  INV_X1    g0693(.A(new_n866), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n894), .B1(new_n657), .B2(new_n647), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n884), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n878), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n897), .A2(KEYINPUT39), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n863), .B1(new_n887), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n689), .A2(new_n469), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n655), .A2(new_n648), .A3(new_n900), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n469), .B(new_n689), .C1(new_n468), .C2(new_n475), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n679), .A2(new_n694), .A3(new_n834), .ZN(new_n904));
  OR2_X1    g0704(.A1(new_n430), .A2(new_n689), .ZN(new_n905));
  AND3_X1   g0705(.A1(new_n904), .A2(KEYINPUT106), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT106), .B1(new_n904), .B2(new_n905), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n897), .B(new_n903), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n658), .A2(new_n687), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n899), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n730), .A2(new_n478), .A3(new_n733), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n660), .ZN(new_n912));
  XOR2_X1   g0712(.A(new_n910), .B(new_n912), .Z(new_n913));
  INV_X1    g0713(.A(KEYINPUT109), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n751), .A2(new_n914), .ZN(new_n915));
  NAND4_X1  g0715(.A1(new_n746), .A2(KEYINPUT109), .A3(KEYINPUT31), .A4(new_n689), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AND4_X1   g0717(.A1(new_n641), .A2(new_n644), .A3(new_n597), .A4(new_n592), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n707), .B1(new_n693), .B2(new_n517), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n918), .A2(new_n919), .A3(new_n611), .A4(new_n694), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(KEYINPUT31), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n917), .B1(new_n921), .B2(new_n747), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n903), .A2(new_n834), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT40), .ZN(new_n924));
  NOR3_X1   g0724(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n915), .A2(new_n916), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n750), .A2(new_n926), .ZN(new_n927));
  AOI22_X1  g0727(.A1(new_n901), .A2(new_n902), .B1(new_n832), .B2(new_n833), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n897), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  XOR2_X1   g0729(.A(KEYINPUT108), .B(KEYINPUT40), .Z(new_n930));
  AOI22_X1  g0730(.A1(new_n886), .A2(new_n925), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n478), .A2(new_n927), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n931), .B(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(G330), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n913), .B(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n269), .B2(new_n682), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n208), .B1(new_n631), .B2(KEYINPUT35), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n937), .B(new_n227), .C1(KEYINPUT35), .C2(new_n631), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(KEYINPUT36), .ZN(new_n939));
  OAI21_X1  g0739(.A(G77), .B1(new_n776), .B2(new_n217), .ZN(new_n940));
  OAI22_X1  g0740(.A1(new_n940), .A2(new_n229), .B1(G50), .B2(new_n217), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n941), .A2(G1), .A3(new_n454), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n936), .A2(new_n939), .A3(new_n942), .ZN(G367));
  NOR2_X1   g0743(.A1(new_n759), .A2(new_n217), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n944), .B1(G159), .B2(new_n769), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n945), .B(new_n249), .C1(new_n202), .C2(new_n773), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n780), .A2(G77), .ZN(new_n947));
  OAI221_X1 g0747(.A(new_n947), .B1(new_n843), .B2(new_n764), .C1(new_n284), .C2(new_n775), .ZN(new_n948));
  AOI211_X1 g0748(.A(new_n946), .B(new_n948), .C1(G143), .C2(new_n787), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n790), .A2(G58), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n765), .A2(G317), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n780), .A2(G97), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n249), .B1(new_n840), .B2(G283), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n774), .A2(new_n531), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n789), .A2(new_n208), .ZN(new_n956));
  AOI22_X1  g0756(.A1(G107), .A2(new_n760), .B1(new_n956), .B2(KEYINPUT46), .ZN(new_n957));
  OAI221_X1 g0757(.A(new_n957), .B1(KEYINPUT46), .B2(new_n956), .C1(new_n798), .C2(new_n770), .ZN(new_n958));
  AOI211_X1 g0758(.A(new_n955), .B(new_n958), .C1(G311), .C2(new_n787), .ZN(new_n959));
  AOI22_X1  g0759(.A1(new_n949), .A2(new_n950), .B1(new_n951), .B2(new_n959), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n960), .B(KEYINPUT47), .Z(new_n961));
  AOI21_X1  g0761(.A(new_n827), .B1(new_n961), .B2(new_n808), .ZN(new_n962));
  OAI221_X1 g0762(.A(new_n812), .B1(new_n222), .B2(new_n579), .C1(new_n240), .C2(new_n815), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n689), .A2(new_n583), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n665), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n965), .B1(new_n674), .B2(new_n964), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n962), .B(new_n963), .C1(new_n825), .C2(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n641), .A2(new_n694), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n689), .A2(new_n640), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n969), .B1(new_n720), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n699), .A2(new_n971), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT112), .Z(new_n973));
  OR2_X1    g0773(.A1(new_n973), .A2(KEYINPUT44), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(KEYINPUT44), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n699), .A2(new_n971), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT45), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n974), .A2(new_n975), .A3(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(new_n710), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n696), .B(new_n697), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(new_n709), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n756), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n756), .B1(new_n979), .B2(new_n983), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n714), .B(KEYINPUT41), .Z(new_n985));
  AOI21_X1  g0785(.A(new_n822), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n971), .B(KEYINPUT110), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n641), .B1(new_n987), .B2(new_n518), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(new_n694), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n971), .A2(new_n698), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT42), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n967), .A2(KEYINPUT43), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n989), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n993), .B(KEYINPUT111), .Z(new_n994));
  AOI21_X1  g0794(.A(new_n992), .B1(new_n989), .B2(new_n991), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT43), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n995), .B1(new_n996), .B2(new_n966), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n994), .A2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n710), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n987), .A2(new_n999), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n998), .B(new_n1000), .Z(new_n1001));
  OAI21_X1  g0801(.A(new_n968), .B1(new_n986), .B2(new_n1001), .ZN(G387));
  OR2_X1    g0802(.A1(new_n756), .A2(new_n982), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1003), .A2(new_n823), .A3(new_n983), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n769), .A2(G311), .B1(new_n531), .B2(new_n840), .ZN(new_n1005));
  INV_X1    g0805(.A(G317), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n1005), .B1(new_n1006), .B2(new_n775), .C1(new_n786), .C2(new_n794), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT48), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n1008), .B1(new_n849), .B2(new_n759), .C1(new_n798), .C2(new_n789), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT49), .ZN(new_n1010));
  OR2_X1    g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n765), .A2(G326), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n249), .B1(new_n780), .B2(G116), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .A4(new_n1014), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n952), .B1(new_n202), .B2(new_n775), .C1(new_n284), .C2(new_n764), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n770), .A2(new_n290), .B1(new_n579), .B2(new_n759), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n331), .B(new_n1017), .C1(G68), .C2(new_n840), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n790), .A2(G77), .ZN(new_n1019));
  INV_X1    g0819(.A(G159), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1018), .B(new_n1019), .C1(new_n1020), .C2(new_n786), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1015), .B1(new_n1016), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1022), .A2(new_n808), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n290), .A2(G50), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT50), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n712), .B1(new_n217), .B2(new_n251), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1026));
  AOI211_X1 g0826(.A(G45), .B(new_n1026), .C1(new_n1025), .C2(new_n1024), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n814), .B1(new_n236), .B2(new_n509), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n249), .B(new_n222), .C1(G116), .C2(new_n572), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1027), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n222), .A2(G107), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n812), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1023), .B(new_n1032), .C1(new_n696), .C2(new_n825), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1004), .B1(new_n821), .B2(new_n981), .C1(new_n827), .C2(new_n1033), .ZN(G393));
  AOI21_X1  g0834(.A(new_n714), .B1(new_n979), .B2(new_n983), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n979), .B2(new_n983), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n979), .A2(new_n821), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n987), .A2(new_n811), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n812), .B1(new_n524), .B2(new_n222), .C1(new_n247), .C2(new_n815), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n770), .A2(new_n202), .B1(new_n251), .B2(new_n759), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n249), .B1(new_n764), .B2(new_n842), .C1(new_n290), .C2(new_n773), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n571), .B2(new_n779), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT51), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n1020), .A2(new_n775), .B1(new_n786), .B2(new_n284), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1043), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n1044), .B2(new_n1045), .C1(new_n217), .C2(new_n789), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n331), .B1(new_n773), .B2(new_n798), .C1(new_n849), .C2(new_n789), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n769), .A2(new_n531), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n208), .B2(new_n759), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1048), .B(new_n1050), .C1(G107), .C2(new_n780), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n805), .A2(new_n775), .B1(new_n786), .B2(new_n1006), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT52), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1051), .B(new_n1053), .C1(new_n794), .C2(new_n764), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1047), .A2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n827), .B1(new_n1055), .B2(new_n808), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1038), .A2(new_n1039), .A3(new_n1056), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1036), .A2(new_n1037), .A3(new_n1057), .ZN(G390));
  AND2_X1   g0858(.A1(new_n834), .A2(G330), .ZN(new_n1059));
  AND2_X1   g0859(.A1(new_n753), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(new_n903), .ZN(new_n1061));
  AND2_X1   g0861(.A1(new_n927), .A2(new_n1059), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1061), .B1(new_n903), .B2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n729), .A2(new_n694), .A3(new_n834), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n905), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n927), .A2(new_n903), .A3(new_n1059), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(new_n1060), .B2(new_n903), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n907), .B2(new_n906), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT114), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1068), .B(KEYINPUT114), .C1(new_n907), .C2(new_n906), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1066), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n478), .A2(G330), .A3(new_n927), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n911), .A2(new_n660), .A3(new_n1074), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT115), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1076), .B(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT113), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1067), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n903), .B1(new_n906), .B2(new_n907), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n863), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n887), .A2(new_n898), .ZN(new_n1084));
  AND2_X1   g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n863), .B1(new_n1065), .B2(new_n903), .ZN(new_n1086));
  AND2_X1   g0886(.A1(new_n1086), .A2(new_n886), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1079), .B(new_n1080), .C1(new_n1085), .C2(new_n1087), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n1083), .A2(new_n1084), .B1(new_n1086), .B2(new_n886), .ZN(new_n1089));
  OAI21_X1  g0889(.A(KEYINPUT113), .B1(new_n1089), .B2(new_n1067), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1089), .A2(new_n1061), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1088), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1078), .A2(new_n1092), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n1088), .A2(new_n1090), .A3(new_n1091), .A4(new_n1076), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1093), .A2(new_n823), .A3(new_n1094), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n1092), .A2(new_n821), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1084), .A2(new_n809), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(KEYINPUT54), .B(G143), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n249), .B1(new_n773), .B2(new_n1098), .C1(new_n775), .C2(new_n847), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n790), .A2(G150), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT53), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(G159), .B2(new_n760), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1102), .B1(new_n843), .B2(new_n770), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n1099), .B(new_n1103), .C1(G50), .C2(new_n780), .ZN(new_n1104));
  INV_X1    g0904(.A(G125), .ZN(new_n1105));
  INV_X1    g0905(.A(G128), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n1104), .B1(new_n1105), .B2(new_n764), .C1(new_n1106), .C2(new_n786), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n331), .B1(new_n770), .B2(new_n499), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n791), .B1(new_n251), .B2(new_n759), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n773), .A2(new_n524), .B1(new_n764), .B2(new_n798), .ZN(new_n1110));
  NOR4_X1   g0910(.A1(new_n838), .A2(new_n1108), .A3(new_n1109), .A4(new_n1110), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n1111), .B1(new_n208), .B2(new_n775), .C1(new_n849), .C2(new_n786), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1107), .A2(new_n1112), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n1113), .A2(new_n808), .B1(new_n290), .B2(new_n859), .ZN(new_n1114));
  AND2_X1   g0914(.A1(new_n1097), .A2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1096), .B1(new_n824), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1095), .A2(new_n1116), .ZN(G378));
  NOR2_X1   g0917(.A1(new_n922), .A2(new_n923), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n885), .A2(new_n878), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n1118), .A2(KEYINPUT40), .A3(new_n1119), .A4(new_n876), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n897), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n920), .A2(KEYINPUT31), .B1(new_n689), .B2(new_n746), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n928), .B1(new_n1122), .B2(new_n917), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n930), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1120), .A2(G330), .A3(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(KEYINPUT116), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT116), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n1120), .A2(new_n1124), .A3(new_n1127), .A4(G330), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n318), .A2(new_n322), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n311), .A2(new_n687), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT55), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1130), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n318), .A2(new_n322), .A3(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1131), .A2(new_n1132), .A3(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1133), .B1(new_n318), .B2(new_n322), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n322), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n1137), .B(new_n1130), .C1(new_n310), .C2(new_n317), .ZN(new_n1138));
  OAI21_X1  g0938(.A(KEYINPUT55), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  AND3_X1   g0939(.A1(new_n1135), .A2(new_n1139), .A3(KEYINPUT56), .ZN(new_n1140));
  AOI21_X1  g0940(.A(KEYINPUT56), .B1(new_n1135), .B2(new_n1139), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1126), .A2(new_n1128), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1135), .A2(new_n1139), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT56), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1135), .A2(new_n1139), .A3(KEYINPUT56), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1148), .A2(new_n1125), .A3(KEYINPUT116), .ZN(new_n1149));
  AND3_X1   g0949(.A1(new_n1143), .A2(new_n910), .A3(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n910), .B1(new_n1143), .B2(new_n1149), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n822), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n858), .A2(new_n202), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n780), .A2(G58), .ZN(new_n1154));
  OAI221_X1 g0954(.A(new_n1154), .B1(new_n849), .B2(new_n764), .C1(new_n579), .C2(new_n773), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n713), .B(new_n1019), .C1(new_n770), .C2(new_n524), .ZN(new_n1156));
  NOR4_X1   g0956(.A1(new_n1155), .A2(new_n249), .A3(new_n944), .A4(new_n1156), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n1157), .B1(new_n499), .B2(new_n775), .C1(new_n208), .C2(new_n786), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1158), .B(KEYINPUT58), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n759), .A2(new_n284), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n843), .A2(new_n773), .B1(new_n789), .B2(new_n1098), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n1160), .B(new_n1161), .C1(G132), .C2(new_n769), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n1162), .B1(new_n1105), .B2(new_n786), .C1(new_n1106), .C2(new_n775), .ZN(new_n1163));
  XOR2_X1   g0963(.A(new_n1163), .B(KEYINPUT59), .Z(new_n1164));
  AOI21_X1  g0964(.A(G41), .B1(new_n780), .B2(G159), .ZN(new_n1165));
  AOI21_X1  g0965(.A(G33), .B1(new_n765), .B2(G124), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(G41), .B1(KEYINPUT3), .B2(G33), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n1159), .B(new_n1167), .C1(G50), .C2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n827), .B1(new_n1169), .B2(new_n808), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1153), .B(new_n1170), .C1(new_n1148), .C2(new_n810), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n1152), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1075), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1143), .A2(new_n910), .A3(new_n1149), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n910), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1128), .A2(new_n1142), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1127), .B1(new_n931), .B2(G330), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1149), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1175), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n1094), .A2(new_n1173), .B1(new_n1174), .B2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n823), .B1(new_n1181), .B2(KEYINPUT57), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1094), .A2(new_n1173), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT117), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1180), .A2(KEYINPUT117), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  AND3_X1   g0987(.A1(new_n1183), .A2(KEYINPUT57), .A3(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1172), .B1(new_n1182), .B2(new_n1188), .ZN(G375));
  NAND2_X1  g0989(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1078), .A2(new_n985), .A3(new_n1190), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n249), .B1(new_n773), .B2(new_n284), .C1(new_n1020), .C2(new_n789), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(G50), .B2(new_n760), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1193), .B(new_n1154), .C1(new_n1106), .C2(new_n764), .ZN(new_n1194));
  XOR2_X1   g0994(.A(new_n1194), .B(KEYINPUT119), .Z(new_n1195));
  NOR2_X1   g0995(.A1(new_n786), .A2(new_n847), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n1196), .A2(KEYINPUT118), .B1(new_n770), .B2(new_n1098), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(KEYINPUT118), .B2(new_n1196), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1195), .B(new_n1198), .C1(new_n843), .C2(new_n775), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n770), .A2(new_n208), .B1(new_n579), .B2(new_n759), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n249), .B(new_n1200), .C1(G283), .C2(new_n774), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(G107), .A2(new_n840), .B1(new_n765), .B2(G303), .ZN(new_n1202));
  AND3_X1   g1002(.A1(new_n1201), .A2(new_n947), .A3(new_n1202), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n1203), .B1(new_n524), .B2(new_n789), .C1(new_n798), .C2(new_n786), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1199), .A2(new_n1204), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n1205), .A2(new_n808), .B1(new_n217), .B2(new_n859), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n901), .A2(new_n902), .A3(new_n809), .ZN(new_n1207));
  AND3_X1   g1007(.A1(new_n1206), .A2(new_n824), .A3(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1073), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1208), .B1(new_n1209), .B2(new_n822), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1191), .A2(new_n1210), .ZN(G381));
  NOR3_X1   g1011(.A1(G387), .A2(G390), .A3(G384), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(G375), .A2(G378), .ZN(new_n1213));
  NOR3_X1   g1013(.A1(G381), .A2(G393), .A3(G396), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .ZN(G407));
  INV_X1    g1015(.A(G213), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(new_n1213), .B2(new_n688), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(G407), .ZN(G409));
  XOR2_X1   g1018(.A(G393), .B(G396), .Z(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(G390), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(G387), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1221), .A2(G387), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1220), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  OR2_X1    g1025(.A1(new_n1221), .A2(G387), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1226), .A2(new_n1219), .A3(new_n1222), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1225), .A2(new_n1227), .ZN(new_n1228));
  OAI211_X1 g1028(.A(G378), .B(new_n1172), .C1(new_n1182), .C2(new_n1188), .ZN(new_n1229));
  AOI21_X1  g1029(.A(KEYINPUT117), .B1(new_n1180), .B2(new_n1174), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1151), .A2(new_n1184), .ZN(new_n1231));
  OAI21_X1  g1031(.A(KEYINPUT120), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT120), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1185), .A2(new_n1233), .A3(new_n1186), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1232), .A2(new_n1234), .A3(new_n822), .ZN(new_n1235));
  AND3_X1   g1035(.A1(new_n1235), .A2(KEYINPUT121), .A3(new_n1171), .ZN(new_n1236));
  AOI21_X1  g1036(.A(KEYINPUT121), .B1(new_n1235), .B2(new_n1171), .ZN(new_n1237));
  AND2_X1   g1037(.A1(new_n1181), .A2(new_n985), .ZN(new_n1238));
  NOR3_X1   g1038(.A1(new_n1236), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1229), .B1(new_n1239), .B2(G378), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1216), .A2(G343), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT60), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n714), .B1(new_n1190), .B2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1076), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1244), .B(new_n1245), .C1(new_n1243), .C2(new_n1190), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n1210), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1247), .A2(new_n837), .A3(new_n861), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1246), .A2(G384), .A3(new_n1210), .ZN(new_n1249));
  AND2_X1   g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1240), .A2(KEYINPUT63), .A3(new_n1242), .A4(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT123), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1235), .A2(new_n1171), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT121), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1238), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1235), .A2(KEYINPUT121), .A3(new_n1171), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1256), .A2(new_n1257), .A3(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(G378), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1241), .B1(new_n1261), .B2(new_n1229), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1262), .A2(KEYINPUT123), .A3(KEYINPUT63), .A4(new_n1250), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1228), .B1(new_n1253), .B2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT61), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT63), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT122), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1240), .A2(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1261), .A2(KEYINPUT122), .A3(new_n1229), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1268), .A2(new_n1242), .A3(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1241), .A2(G2897), .ZN(new_n1271));
  XOR2_X1   g1071(.A(new_n1250), .B(new_n1271), .Z(new_n1272));
  AOI21_X1  g1072(.A(new_n1266), .B1(new_n1270), .B2(new_n1272), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1268), .A2(new_n1242), .A3(new_n1250), .A4(new_n1269), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  OAI211_X1 g1075(.A(new_n1264), .B(new_n1265), .C1(new_n1273), .C2(new_n1275), .ZN(new_n1276));
  AND4_X1   g1076(.A1(KEYINPUT62), .A2(new_n1240), .A3(new_n1242), .A4(new_n1250), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT62), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1277), .B1(new_n1274), .B2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1240), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1272), .B1(new_n1280), .B2(new_n1241), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n1265), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1228), .B1(new_n1279), .B2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1276), .A2(new_n1283), .ZN(G405));
  NAND2_X1  g1084(.A1(G375), .A2(new_n1260), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT124), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(G375), .A2(new_n1260), .A3(KEYINPUT124), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1287), .A2(new_n1229), .A3(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT125), .ZN(new_n1290));
  AND3_X1   g1090(.A1(new_n1248), .A2(new_n1290), .A3(new_n1249), .ZN(new_n1291));
  OR2_X1    g1091(.A1(new_n1291), .A2(KEYINPUT126), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1289), .A2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1250), .A2(KEYINPUT126), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1294), .B1(new_n1291), .B2(KEYINPUT126), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1295), .A2(new_n1229), .A3(new_n1287), .A4(new_n1288), .ZN(new_n1296));
  AOI211_X1 g1096(.A(KEYINPUT127), .B(new_n1228), .C1(new_n1293), .C2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT127), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1293), .A2(new_n1296), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1228), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1298), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1302));
  NOR3_X1   g1102(.A1(new_n1297), .A2(new_n1301), .A3(new_n1302), .ZN(G402));
endmodule


