//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 1 1 0 1 1 1 0 0 0 0 1 1 0 1 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 0 1 1 1 0 0 0 0 1 1 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n645,
    new_n646, new_n647, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n800, new_n801, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n809, new_n810, new_n811, new_n812, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n887, new_n888, new_n890, new_n891, new_n892,
    new_n894, new_n895, new_n896, new_n897, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933;
  INV_X1    g000(.A(KEYINPUT102), .ZN(new_n202));
  NOR3_X1   g001(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n203));
  OAI21_X1  g002(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n204));
  AOI21_X1  g003(.A(new_n203), .B1(KEYINPUT91), .B2(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(KEYINPUT91), .B2(new_n204), .ZN(new_n206));
  XOR2_X1   g005(.A(KEYINPUT92), .B(G29gat), .Z(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G36gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT15), .ZN(new_n210));
  NOR2_X1   g009(.A1(G43gat), .A2(G50gat), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(G43gat), .A2(G50gat), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n210), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n209), .A2(new_n214), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n214), .B1(G36gat), .B2(new_n207), .ZN(new_n216));
  XNOR2_X1  g015(.A(KEYINPUT93), .B(G50gat), .ZN(new_n217));
  OAI211_X1 g016(.A(new_n210), .B(new_n213), .C1(new_n217), .C2(G43gat), .ZN(new_n218));
  INV_X1    g017(.A(new_n203), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n219), .A2(KEYINPUT94), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT94), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n204), .B1(new_n203), .B2(new_n221), .ZN(new_n222));
  OAI211_X1 g021(.A(new_n216), .B(new_n218), .C1(new_n220), .C2(new_n222), .ZN(new_n223));
  AND2_X1   g022(.A1(new_n215), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n202), .B1(new_n224), .B2(KEYINPUT17), .ZN(new_n225));
  NAND2_X1  g024(.A1(G85gat), .A2(G92gat), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n226), .B(KEYINPUT7), .ZN(new_n227));
  NAND2_X1  g026(.A1(G99gat), .A2(G106gat), .ZN(new_n228));
  INV_X1    g027(.A(G85gat), .ZN(new_n229));
  INV_X1    g028(.A(G92gat), .ZN(new_n230));
  AOI22_X1  g029(.A1(KEYINPUT8), .A2(new_n228), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n227), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(G99gat), .B(G106gat), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n232), .B(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT17), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n236), .B1(new_n235), .B2(KEYINPUT102), .ZN(new_n237));
  AOI22_X1  g036(.A1(new_n225), .A2(new_n235), .B1(new_n224), .B2(new_n237), .ZN(new_n238));
  AND2_X1   g037(.A1(G232gat), .A2(G233gat), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n238), .B1(KEYINPUT41), .B2(new_n239), .ZN(new_n240));
  XOR2_X1   g039(.A(G190gat), .B(G218gat), .Z(new_n241));
  XNOR2_X1  g040(.A(new_n241), .B(KEYINPUT103), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT104), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n240), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(G134gat), .B(G162gat), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n242), .A2(new_n243), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n239), .A2(KEYINPUT41), .ZN(new_n250));
  XOR2_X1   g049(.A(new_n249), .B(new_n250), .Z(new_n251));
  OAI21_X1  g050(.A(new_n246), .B1(new_n240), .B2(new_n244), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n248), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n251), .B1(new_n248), .B2(new_n252), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NOR2_X1   g056(.A1(G71gat), .A2(G78gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(G71gat), .A2(G78gat), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n258), .B1(KEYINPUT96), .B2(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n260), .B1(KEYINPUT96), .B2(new_n259), .ZN(new_n261));
  NOR2_X1   g060(.A1(KEYINPUT96), .A2(KEYINPUT9), .ZN(new_n262));
  INV_X1    g061(.A(G64gat), .ZN(new_n263));
  OR2_X1    g062(.A1(new_n263), .A2(G57gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(G57gat), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n262), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n261), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(KEYINPUT97), .B(G57gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(G64gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n258), .A2(KEYINPUT9), .ZN(new_n270));
  AOI22_X1  g069(.A1(new_n269), .A2(new_n265), .B1(new_n259), .B2(new_n270), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n272), .A2(KEYINPUT21), .ZN(new_n273));
  NAND2_X1  g072(.A1(G231gat), .A2(G233gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(G127gat), .B(G155gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n276), .B(KEYINPUT20), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n275), .B(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G15gat), .B(G22gat), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT16), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n279), .B1(new_n280), .B2(G1gat), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n281), .B1(G1gat), .B2(new_n279), .ZN(new_n282));
  OR2_X1    g081(.A1(new_n282), .A2(G8gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(G8gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n285), .B1(KEYINPUT21), .B2(new_n272), .ZN(new_n286));
  XOR2_X1   g085(.A(new_n286), .B(KEYINPUT101), .Z(new_n287));
  XNOR2_X1  g086(.A(new_n278), .B(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(KEYINPUT100), .B(KEYINPUT19), .ZN(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT98), .B(KEYINPUT99), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n289), .B(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(G183gat), .B(G211gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n291), .B(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n288), .B(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n257), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G8gat), .B(G36gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(G64gat), .B(G92gat), .ZN(new_n297));
  XOR2_X1   g096(.A(new_n296), .B(new_n297), .Z(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n300));
  XOR2_X1   g099(.A(new_n300), .B(KEYINPUT64), .Z(new_n301));
  OAI21_X1  g100(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n302));
  INV_X1    g101(.A(G183gat), .ZN(new_n303));
  INV_X1    g102(.A(G190gat), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  NOR2_X1   g105(.A1(G169gat), .A2(G176gat), .ZN(new_n307));
  OR2_X1    g106(.A1(new_n307), .A2(KEYINPUT23), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(KEYINPUT23), .ZN(new_n309));
  NAND2_X1  g108(.A1(G169gat), .A2(G176gat), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n311), .A2(KEYINPUT25), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n306), .A2(new_n308), .A3(new_n309), .A4(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n305), .A2(new_n300), .ZN(new_n314));
  AOI22_X1  g113(.A1(new_n307), .A2(KEYINPUT23), .B1(new_n310), .B2(KEYINPUT65), .ZN(new_n315));
  OR2_X1    g114(.A1(new_n310), .A2(KEYINPUT65), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n314), .A2(new_n308), .A3(new_n315), .A4(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(KEYINPUT25), .ZN(new_n318));
  XNOR2_X1  g117(.A(KEYINPUT27), .B(G183gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(new_n304), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n320), .B(KEYINPUT28), .ZN(new_n321));
  INV_X1    g120(.A(new_n307), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n311), .B1(new_n322), .B2(KEYINPUT26), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n323), .B1(KEYINPUT26), .B2(new_n322), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n324), .B1(new_n303), .B2(new_n304), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n313), .B(new_n318), .C1(new_n321), .C2(new_n325), .ZN(new_n326));
  AND2_X1   g125(.A1(G226gat), .A2(G233gat), .ZN(new_n327));
  AND2_X1   g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT29), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n327), .B1(new_n326), .B2(new_n329), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(G211gat), .B(G218gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n332), .B(KEYINPUT72), .ZN(new_n333));
  OR2_X1    g132(.A1(G197gat), .A2(G204gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(G197gat), .A2(G204gat), .ZN(new_n335));
  AND2_X1   g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n337));
  OR2_X1    g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n333), .B(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n331), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n337), .B1(new_n334), .B2(new_n335), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n333), .B(new_n341), .ZN(new_n342));
  XOR2_X1   g141(.A(KEYINPUT73), .B(KEYINPUT29), .Z(new_n343));
  AOI21_X1  g142(.A(new_n327), .B1(new_n326), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n342), .B1(new_n328), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n340), .A2(KEYINPUT74), .A3(new_n345), .ZN(new_n346));
  OR2_X1    g145(.A1(new_n345), .A2(KEYINPUT74), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n299), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT75), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT30), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(KEYINPUT75), .B1(new_n348), .B2(KEYINPUT30), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n346), .A2(new_n347), .A3(new_n299), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n348), .A2(KEYINPUT30), .ZN(new_n356));
  AND3_X1   g155(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(G134gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(G127gat), .ZN(new_n359));
  INV_X1    g158(.A(G127gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(G134gat), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT1), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n359), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(G113gat), .B(G120gat), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n363), .B1(KEYINPUT67), .B2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(G120gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(G113gat), .ZN(new_n367));
  INV_X1    g166(.A(G113gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(G120gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT67), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n370), .A2(new_n362), .ZN(new_n373));
  AND3_X1   g172(.A1(new_n358), .A2(KEYINPUT66), .A3(G127gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(G127gat), .B(G134gat), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT66), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n374), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  AOI22_X1  g176(.A1(new_n365), .A2(new_n372), .B1(new_n373), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(G155gat), .A2(G162gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT2), .ZN(new_n380));
  INV_X1    g179(.A(G141gat), .ZN(new_n381));
  INV_X1    g180(.A(G148gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(G141gat), .A2(G148gat), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n380), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(G155gat), .B(G162gat), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n383), .A2(KEYINPUT76), .A3(new_n384), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  AND2_X1   g187(.A1(G141gat), .A2(G148gat), .ZN(new_n389));
  NOR2_X1   g188(.A1(G141gat), .A2(G148gat), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  AND2_X1   g190(.A1(G155gat), .A2(G162gat), .ZN(new_n392));
  NOR2_X1   g191(.A1(G155gat), .A2(G162gat), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  OAI211_X1 g193(.A(new_n380), .B(new_n391), .C1(new_n394), .C2(KEYINPUT76), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n388), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT4), .B1(new_n378), .B2(new_n396), .ZN(new_n397));
  AND2_X1   g196(.A1(new_n388), .A2(new_n395), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n367), .A2(new_n369), .A3(KEYINPUT67), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n399), .A2(new_n362), .A3(new_n375), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n364), .A2(KEYINPUT67), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n359), .A2(new_n361), .A3(new_n376), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n358), .A2(KEYINPUT66), .A3(G127gat), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n364), .A2(KEYINPUT1), .ZN(new_n405));
  OAI22_X1  g204(.A1(new_n400), .A2(new_n401), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g205(.A(KEYINPUT78), .B1(new_n398), .B2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT78), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n378), .A2(new_n408), .A3(new_n396), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n397), .B1(new_n410), .B2(KEYINPUT4), .ZN(new_n411));
  XOR2_X1   g210(.A(KEYINPUT80), .B(KEYINPUT5), .Z(new_n412));
  NAND2_X1  g211(.A1(G225gat), .A2(G233gat), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n378), .B1(KEYINPUT3), .B2(new_n398), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT3), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n396), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n414), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n411), .A2(new_n412), .A3(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(KEYINPUT4), .B1(new_n398), .B2(new_n406), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(KEYINPUT77), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT77), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n423), .B(KEYINPUT4), .C1(new_n398), .C2(new_n406), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT4), .B1(new_n407), .B2(new_n409), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n418), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n398), .A2(new_n406), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n407), .A2(new_n409), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(new_n414), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(KEYINPUT79), .ZN(new_n431));
  INV_X1    g230(.A(new_n412), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT79), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n429), .A2(new_n433), .A3(new_n414), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n427), .A2(new_n431), .A3(new_n432), .A4(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT81), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT4), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n408), .B1(new_n378), .B2(new_n396), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n377), .A2(new_n373), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n372), .A2(new_n362), .A3(new_n375), .A4(new_n399), .ZN(new_n440));
  AND4_X1   g239(.A1(new_n408), .A2(new_n396), .A3(new_n439), .A4(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n437), .B1(new_n438), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n442), .A2(new_n422), .A3(new_n424), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n412), .B1(new_n443), .B2(new_n418), .ZN(new_n444));
  AND3_X1   g243(.A1(new_n429), .A2(new_n433), .A3(new_n414), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n433), .B1(new_n429), .B2(new_n414), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT81), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n444), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n420), .B1(new_n436), .B2(new_n449), .ZN(new_n450));
  XOR2_X1   g249(.A(G1gat), .B(G29gat), .Z(new_n451));
  XNOR2_X1  g250(.A(G57gat), .B(G85gat), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n451), .B(new_n452), .ZN(new_n453));
  XNOR2_X1  g252(.A(KEYINPUT82), .B(KEYINPUT0), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n453), .B(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n450), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT6), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n435), .A2(KEYINPUT81), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n448), .B1(new_n444), .B2(new_n447), .ZN(new_n460));
  OAI211_X1 g259(.A(new_n456), .B(new_n419), .C1(new_n459), .C2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT6), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT83), .B1(new_n450), .B2(new_n456), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n419), .B1(new_n459), .B2(new_n460), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT83), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n465), .A2(new_n466), .A3(new_n455), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n463), .B1(new_n464), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT84), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n458), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT6), .B1(new_n450), .B2(new_n456), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n466), .B1(new_n465), .B2(new_n455), .ZN(new_n472));
  NOR3_X1   g271(.A1(new_n450), .A2(KEYINPUT83), .A3(new_n456), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n469), .B(new_n471), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n357), .B1(new_n470), .B2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT85), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n458), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n479), .B1(new_n480), .B2(KEYINPUT84), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(new_n474), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n482), .A2(KEYINPUT85), .A3(new_n357), .ZN(new_n483));
  INV_X1    g282(.A(G227gat), .ZN(new_n484));
  INV_X1    g283(.A(G233gat), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT68), .ZN(new_n487));
  OR3_X1    g286(.A1(new_n326), .A2(new_n487), .A3(new_n378), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n378), .A2(new_n487), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n406), .A2(KEYINPUT68), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n326), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n486), .B1(new_n488), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT34), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI211_X1 g293(.A(KEYINPUT34), .B(new_n486), .C1(new_n488), .C2(new_n491), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n488), .A2(new_n486), .A3(new_n491), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(KEYINPUT32), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT33), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  XOR2_X1   g300(.A(G15gat), .B(G43gat), .Z(new_n502));
  XNOR2_X1  g301(.A(G71gat), .B(G99gat), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n502), .B(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n499), .A2(new_n501), .A3(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n504), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n498), .B(KEYINPUT32), .C1(new_n500), .C2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT69), .ZN(new_n509));
  AND3_X1   g308(.A1(new_n497), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n509), .B1(new_n497), .B2(new_n508), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n496), .A2(new_n505), .A3(new_n507), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT70), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT70), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n496), .A2(new_n505), .A3(new_n515), .A4(new_n507), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n512), .A2(new_n517), .ZN(new_n518));
  AND2_X1   g317(.A1(G228gat), .A2(G233gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n417), .A2(new_n343), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n342), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(KEYINPUT3), .B1(new_n339), .B2(new_n329), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n519), .B(new_n521), .C1(new_n522), .C2(new_n396), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT87), .ZN(new_n524));
  INV_X1    g323(.A(new_n343), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n524), .B1(new_n342), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n339), .A2(KEYINPUT87), .A3(new_n343), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n526), .A2(new_n527), .A3(new_n416), .ZN(new_n528));
  AOI22_X1  g327(.A1(new_n528), .A2(new_n398), .B1(new_n342), .B2(new_n520), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n523), .B1(new_n529), .B2(new_n519), .ZN(new_n530));
  OR2_X1    g329(.A1(new_n530), .A2(G22gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT88), .ZN(new_n532));
  OR3_X1    g331(.A1(new_n530), .A2(KEYINPUT88), .A3(G22gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n530), .A2(G22gat), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(G78gat), .B(G106gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(KEYINPUT31), .B(G50gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n536), .B(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(KEYINPUT86), .ZN(new_n539));
  AND2_X1   g338(.A1(new_n534), .A2(new_n538), .ZN(new_n540));
  AOI22_X1  g339(.A1(new_n535), .A2(new_n539), .B1(new_n531), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n518), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n478), .A2(new_n483), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT35), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n545));
  NOR3_X1   g344(.A1(new_n545), .A2(new_n541), .A3(KEYINPUT35), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n458), .B1(new_n463), .B2(new_n457), .ZN(new_n547));
  AND3_X1   g346(.A1(new_n514), .A2(KEYINPUT71), .A3(new_n516), .ZN(new_n548));
  AOI21_X1  g347(.A(KEYINPUT71), .B1(new_n514), .B2(new_n516), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n496), .B1(new_n505), .B2(new_n507), .ZN(new_n550));
  NOR3_X1   g349(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n546), .A2(new_n547), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n544), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n478), .A2(new_n483), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(new_n541), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n415), .A2(new_n417), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n411), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(new_n414), .ZN(new_n558));
  OAI211_X1 g357(.A(new_n558), .B(KEYINPUT39), .C1(new_n414), .C2(new_n429), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n559), .B(new_n456), .C1(KEYINPUT39), .C2(new_n558), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT40), .ZN(new_n561));
  AND2_X1   g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n560), .A2(new_n561), .ZN(new_n563));
  NOR3_X1   g362(.A1(new_n562), .A2(new_n563), .A3(new_n457), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n541), .B1(new_n545), .B2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT37), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n355), .B1(new_n566), .B2(new_n298), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n342), .B1(new_n328), .B2(new_n330), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT89), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n566), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  OR2_X1    g370(.A1(new_n328), .A2(new_n344), .ZN(new_n572));
  OAI211_X1 g371(.A(KEYINPUT89), .B(new_n568), .C1(new_n572), .C2(new_n342), .ZN(new_n573));
  AOI21_X1  g372(.A(KEYINPUT38), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n567), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(new_n349), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT38), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n346), .A2(new_n347), .A3(KEYINPUT37), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n577), .B1(new_n567), .B2(new_n578), .ZN(new_n579));
  OR3_X1    g378(.A1(new_n547), .A2(new_n576), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT36), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n582), .B1(new_n512), .B2(new_n517), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n583), .B1(new_n551), .B2(new_n582), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n555), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n295), .B1(new_n553), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n283), .A2(new_n236), .A3(new_n284), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n224), .B(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(G229gat), .A2(G233gat), .ZN(new_n591));
  AND2_X1   g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  XOR2_X1   g391(.A(new_n591), .B(KEYINPUT13), .Z(new_n593));
  XOR2_X1   g392(.A(new_n224), .B(new_n285), .Z(new_n594));
  AOI22_X1  g393(.A1(new_n592), .A2(KEYINPUT18), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n595), .B1(KEYINPUT18), .B2(new_n592), .ZN(new_n596));
  XNOR2_X1  g395(.A(G113gat), .B(G141gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(G197gat), .ZN(new_n598));
  XOR2_X1   g397(.A(KEYINPUT11), .B(G169gat), .Z(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(KEYINPUT90), .B(KEYINPUT12), .ZN(new_n601));
  XOR2_X1   g400(.A(new_n600), .B(new_n601), .Z(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n596), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT95), .ZN(new_n605));
  OR3_X1    g404(.A1(new_n592), .A2(new_n605), .A3(KEYINPUT18), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n605), .B1(new_n592), .B2(KEYINPUT18), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n606), .A2(new_n595), .A3(new_n602), .A4(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(G230gat), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n611), .A2(new_n485), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n234), .A2(new_n272), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT105), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  OR2_X1    g415(.A1(new_n234), .A2(new_n272), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n618), .A2(KEYINPUT10), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT10), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n614), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n613), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n618), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n622), .B1(new_n613), .B2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(G120gat), .B(G148gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(G176gat), .B(G204gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  OR2_X1    g426(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n624), .A2(new_n627), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n610), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n588), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n632), .A2(new_n482), .ZN(new_n633));
  XOR2_X1   g432(.A(new_n633), .B(G1gat), .Z(G1324gat));
  XOR2_X1   g433(.A(KEYINPUT106), .B(KEYINPUT16), .Z(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(G8gat), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n588), .A2(new_n631), .A3(new_n545), .A4(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(G8gat), .B1(new_n632), .B2(new_n357), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(new_n637), .ZN(new_n639));
  MUX2_X1   g438(.A(new_n637), .B(new_n639), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g439(.A(G15gat), .B1(new_n632), .B2(new_n584), .ZN(new_n641));
  INV_X1    g440(.A(new_n551), .ZN(new_n642));
  OR2_X1    g441(.A1(new_n642), .A2(G15gat), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n641), .B1(new_n632), .B2(new_n643), .ZN(G1326gat));
  INV_X1    g443(.A(new_n541), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n632), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g445(.A(KEYINPUT43), .B(G22gat), .Z(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(G1327gat));
  INV_X1    g447(.A(new_n294), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n631), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n552), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n652), .B1(new_n543), .B2(KEYINPUT35), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n585), .B1(new_n554), .B2(new_n541), .ZN(new_n654));
  OAI211_X1 g453(.A(new_n256), .B(new_n651), .C1(new_n653), .C2(new_n654), .ZN(new_n655));
  NOR3_X1   g454(.A1(new_n655), .A2(new_n482), .A3(new_n207), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n656), .B(KEYINPUT45), .Z(new_n657));
  OAI21_X1  g456(.A(new_n256), .B1(new_n653), .B2(new_n654), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(KEYINPUT44), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT107), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n660), .B1(new_n254), .B2(new_n255), .ZN(new_n661));
  INV_X1    g460(.A(new_n255), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n662), .A2(KEYINPUT107), .A3(new_n253), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n665), .A2(KEYINPUT44), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n666), .B1(new_n653), .B2(new_n654), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n650), .B1(new_n659), .B2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n207), .B1(new_n669), .B2(new_n482), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n657), .A2(new_n670), .ZN(G1328gat));
  OAI21_X1  g470(.A(G36gat), .B1(new_n669), .B2(new_n357), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n655), .A2(G36gat), .A3(new_n357), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(KEYINPUT46), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n672), .A2(new_n674), .ZN(G1329gat));
  INV_X1    g474(.A(KEYINPUT47), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n257), .B1(new_n553), .B2(new_n587), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT109), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n642), .A2(G43gat), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n677), .A2(new_n678), .A3(new_n651), .A4(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n679), .ZN(new_n681));
  OAI21_X1  g480(.A(KEYINPUT109), .B1(new_n655), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(KEYINPUT108), .ZN(new_n684));
  INV_X1    g483(.A(G43gat), .ZN(new_n685));
  INV_X1    g484(.A(new_n584), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n685), .B1(new_n668), .B2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n683), .ZN(new_n688));
  OAI211_X1 g487(.A(new_n676), .B(new_n684), .C1(new_n687), .C2(new_n688), .ZN(new_n689));
  AOI211_X1 g488(.A(new_n584), .B(new_n650), .C1(new_n659), .C2(new_n667), .ZN(new_n690));
  OAI221_X1 g489(.A(new_n683), .B1(KEYINPUT108), .B2(KEYINPUT47), .C1(new_n690), .C2(new_n685), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n689), .A2(new_n691), .ZN(G1330gat));
  AND2_X1   g491(.A1(new_n541), .A2(new_n217), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n668), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  OR2_X1    g494(.A1(new_n655), .A2(KEYINPUT110), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n645), .B1(new_n655), .B2(KEYINPUT110), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n217), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(KEYINPUT48), .B1(new_n695), .B2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT48), .ZN(new_n700));
  AND2_X1   g499(.A1(new_n696), .A2(new_n697), .ZN(new_n701));
  OAI211_X1 g500(.A(new_n700), .B(new_n694), .C1(new_n701), .C2(new_n217), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n699), .A2(new_n702), .ZN(G1331gat));
  INV_X1    g502(.A(new_n630), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n704), .A2(new_n609), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n588), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n706), .A2(new_n482), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(new_n268), .ZN(G1332gat));
  INV_X1    g507(.A(new_n706), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT49), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n263), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n357), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n709), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  OAI211_X1 g512(.A(new_n710), .B(new_n263), .C1(new_n706), .C2(new_n357), .ZN(new_n714));
  XNOR2_X1  g513(.A(KEYINPUT111), .B(KEYINPUT112), .ZN(new_n715));
  AND3_X1   g514(.A1(new_n713), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n715), .B1(new_n713), .B2(new_n714), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n716), .A2(new_n717), .ZN(G1333gat));
  OR3_X1    g517(.A1(new_n706), .A2(G71gat), .A3(new_n642), .ZN(new_n719));
  OAI21_X1  g518(.A(G71gat), .B1(new_n706), .B2(new_n584), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT50), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n719), .A2(KEYINPUT50), .A3(new_n720), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(G1334gat));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n541), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g526(.A1(new_n294), .A2(new_n609), .ZN(new_n728));
  OAI211_X1 g527(.A(new_n256), .B(new_n728), .C1(new_n653), .C2(new_n654), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT51), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n729), .B(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n482), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n731), .A2(new_n229), .A3(new_n732), .A4(new_n630), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n728), .A2(new_n630), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n734), .B1(new_n659), .B2(new_n667), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n735), .A2(new_n732), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n733), .B1(new_n736), .B2(new_n229), .ZN(G1336gat));
  NOR3_X1   g536(.A1(new_n357), .A2(G92gat), .A3(new_n704), .ZN(new_n738));
  AOI21_X1  g537(.A(KEYINPUT52), .B1(new_n731), .B2(new_n738), .ZN(new_n739));
  AOI211_X1 g538(.A(new_n357), .B(new_n734), .C1(new_n659), .C2(new_n667), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n739), .B1(new_n230), .B2(new_n740), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n230), .B1(new_n735), .B2(new_n545), .ZN(new_n742));
  AND3_X1   g541(.A1(new_n729), .A2(KEYINPUT113), .A3(KEYINPUT51), .ZN(new_n743));
  AOI21_X1  g542(.A(KEYINPUT51), .B1(new_n729), .B2(KEYINPUT113), .ZN(new_n744));
  INV_X1    g543(.A(new_n738), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n743), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(KEYINPUT52), .B1(new_n742), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n741), .A2(new_n747), .ZN(G1337gat));
  INV_X1    g547(.A(G99gat), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n731), .A2(new_n749), .A3(new_n630), .A4(new_n551), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n735), .A2(new_n686), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n750), .B1(new_n751), .B2(new_n749), .ZN(G1338gat));
  NOR3_X1   g551(.A1(new_n645), .A2(G106gat), .A3(new_n704), .ZN(new_n753));
  AOI21_X1  g552(.A(KEYINPUT53), .B1(new_n731), .B2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(G106gat), .ZN(new_n755));
  AOI211_X1 g554(.A(new_n645), .B(new_n734), .C1(new_n659), .C2(new_n667), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n754), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n755), .B1(new_n735), .B2(new_n541), .ZN(new_n758));
  INV_X1    g557(.A(new_n753), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n743), .A2(new_n744), .A3(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(KEYINPUT53), .B1(new_n758), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n757), .A2(new_n761), .ZN(G1339gat));
  OR3_X1    g561(.A1(new_n619), .A2(new_n613), .A3(new_n621), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n763), .A2(KEYINPUT54), .A3(new_n622), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT54), .ZN(new_n765));
  OAI211_X1 g564(.A(new_n765), .B(new_n613), .C1(new_n619), .C2(new_n621), .ZN(new_n766));
  AND3_X1   g565(.A1(new_n766), .A2(KEYINPUT114), .A3(new_n627), .ZN(new_n767));
  AOI21_X1  g566(.A(KEYINPUT114), .B1(new_n766), .B2(new_n627), .ZN(new_n768));
  OAI211_X1 g567(.A(KEYINPUT55), .B(new_n764), .C1(new_n767), .C2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n628), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT115), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n769), .A2(KEYINPUT115), .A3(new_n628), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n764), .B1(new_n767), .B2(new_n768), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT55), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n772), .A2(new_n609), .A3(new_n773), .A4(new_n776), .ZN(new_n777));
  OR2_X1    g576(.A1(new_n590), .A2(new_n591), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(KEYINPUT116), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n779), .B1(new_n593), .B2(new_n594), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n778), .A2(KEYINPUT116), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n600), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  AND2_X1   g581(.A1(new_n782), .A2(new_n608), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n630), .A2(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n664), .B1(new_n777), .B2(new_n784), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n772), .A2(new_n783), .A3(new_n773), .A4(new_n776), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n786), .A2(new_n665), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n649), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n630), .A2(new_n609), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n295), .A2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n482), .B1(new_n788), .B2(new_n792), .ZN(new_n793));
  AND3_X1   g592(.A1(new_n793), .A2(new_n357), .A3(new_n542), .ZN(new_n794));
  AOI21_X1  g593(.A(G113gat), .B1(new_n794), .B2(new_n609), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n541), .B1(new_n788), .B2(new_n792), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n796), .A2(new_n732), .A3(new_n357), .A4(new_n551), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n797), .A2(new_n368), .A3(new_n610), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n795), .A2(new_n798), .ZN(G1340gat));
  AOI21_X1  g598(.A(G120gat), .B1(new_n794), .B2(new_n630), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n797), .A2(new_n366), .A3(new_n704), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n800), .A2(new_n801), .ZN(G1341gat));
  NOR3_X1   g601(.A1(new_n797), .A2(new_n360), .A3(new_n649), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n794), .A2(new_n294), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT117), .ZN(new_n805));
  OR2_X1    g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(G127gat), .B1(new_n804), .B2(new_n805), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n803), .B1(new_n806), .B2(new_n807), .ZN(G1342gat));
  NAND3_X1  g607(.A1(new_n794), .A2(new_n358), .A3(new_n256), .ZN(new_n809));
  OR2_X1    g608(.A1(new_n809), .A2(KEYINPUT56), .ZN(new_n810));
  OAI21_X1  g609(.A(G134gat), .B1(new_n797), .B2(new_n257), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(KEYINPUT56), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n810), .A2(new_n811), .A3(new_n812), .ZN(G1343gat));
  NAND2_X1  g612(.A1(new_n584), .A2(new_n541), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n357), .B1(new_n814), .B2(KEYINPUT119), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n815), .B1(KEYINPUT119), .B2(new_n814), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n793), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n609), .A2(new_n381), .ZN(new_n818));
  XNOR2_X1  g617(.A(new_n818), .B(KEYINPUT120), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT58), .ZN(new_n820));
  OAI22_X1  g619(.A1(new_n817), .A2(new_n819), .B1(KEYINPUT121), .B2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT57), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n645), .A2(new_n822), .ZN(new_n823));
  OR2_X1    g622(.A1(new_n786), .A2(new_n665), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n766), .A2(new_n627), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT114), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n766), .A2(KEYINPUT114), .A3(new_n627), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n622), .A2(KEYINPUT54), .ZN(new_n829));
  AOI22_X1  g628(.A1(new_n827), .A2(new_n828), .B1(new_n763), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n609), .B1(new_n830), .B2(KEYINPUT55), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n784), .B1(new_n831), .B2(new_n770), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(new_n257), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n294), .B1(new_n824), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n823), .B1(new_n834), .B2(new_n791), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n645), .B1(new_n788), .B2(new_n792), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n835), .B1(new_n836), .B2(KEYINPUT57), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n584), .A2(new_n732), .A3(new_n357), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n838), .B(KEYINPUT118), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n837), .A2(new_n609), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n821), .B1(new_n840), .B2(G141gat), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n820), .A2(KEYINPUT121), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n841), .B(new_n842), .ZN(G1344gat));
  AND2_X1   g642(.A1(new_n837), .A2(new_n839), .ZN(new_n844));
  AOI211_X1 g643(.A(KEYINPUT59), .B(new_n382), .C1(new_n844), .C2(new_n630), .ZN(new_n845));
  AOI22_X1  g644(.A1(new_n770), .A2(new_n771), .B1(new_n775), .B2(new_n774), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n846), .A2(new_n256), .A3(new_n783), .A4(new_n773), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n833), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n649), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT123), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n850), .B1(new_n295), .B2(new_n790), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n257), .A2(new_n789), .A3(KEYINPUT123), .A4(new_n294), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n849), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(KEYINPUT57), .B1(new_n855), .B2(new_n541), .ZN(new_n856));
  INV_X1    g655(.A(new_n823), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n857), .B1(new_n788), .B2(new_n792), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n839), .A2(new_n630), .ZN(new_n860));
  OAI21_X1  g659(.A(G148gat), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  XNOR2_X1  g660(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n630), .A2(new_n382), .ZN(new_n864));
  OAI22_X1  g663(.A1(new_n845), .A2(new_n863), .B1(new_n817), .B2(new_n864), .ZN(G1345gat));
  INV_X1    g664(.A(G155gat), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n866), .B1(new_n844), .B2(new_n294), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n817), .A2(G155gat), .A3(new_n649), .ZN(new_n868));
  OR2_X1    g667(.A1(new_n867), .A2(new_n868), .ZN(G1346gat));
  NAND4_X1  g668(.A1(new_n837), .A2(G162gat), .A3(new_n664), .A4(new_n839), .ZN(new_n870));
  INV_X1    g669(.A(G162gat), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n871), .B1(new_n817), .B2(new_n257), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  XOR2_X1   g672(.A(new_n873), .B(KEYINPUT124), .Z(G1347gat));
  NAND4_X1  g673(.A1(new_n796), .A2(new_n482), .A3(new_n545), .A4(new_n551), .ZN(new_n875));
  INV_X1    g674(.A(G169gat), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n875), .A2(new_n876), .A3(new_n610), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n788), .A2(new_n792), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n482), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT125), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n357), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n878), .A2(KEYINPUT125), .A3(new_n482), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n881), .A2(new_n542), .A3(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(new_n609), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n877), .B1(new_n885), .B2(new_n876), .ZN(G1348gat));
  OAI21_X1  g685(.A(G176gat), .B1(new_n875), .B2(new_n704), .ZN(new_n887));
  OR2_X1    g686(.A1(new_n704), .A2(G176gat), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n887), .B1(new_n883), .B2(new_n888), .ZN(G1349gat));
  OAI21_X1  g688(.A(G183gat), .B1(new_n875), .B2(new_n649), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n294), .A2(new_n319), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n890), .B1(new_n883), .B2(new_n891), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n892), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g692(.A1(new_n884), .A2(new_n304), .A3(new_n664), .ZN(new_n894));
  OAI21_X1  g693(.A(G190gat), .B1(new_n875), .B2(new_n257), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n895), .A2(KEYINPUT61), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n895), .A2(KEYINPUT61), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n894), .B1(new_n896), .B2(new_n897), .ZN(G1351gat));
  INV_X1    g697(.A(new_n814), .ZN(new_n899));
  AND3_X1   g698(.A1(new_n881), .A2(new_n899), .A3(new_n882), .ZN(new_n900));
  AOI21_X1  g699(.A(G197gat), .B1(new_n900), .B2(new_n609), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT126), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n902), .B1(new_n856), .B2(new_n858), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n878), .A2(new_n823), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n853), .B1(new_n848), .B2(new_n649), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n822), .B1(new_n905), .B2(new_n645), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n904), .A2(new_n906), .A3(KEYINPUT126), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n903), .A2(new_n907), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n686), .A2(new_n732), .A3(new_n357), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n609), .A2(G197gat), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n901), .B1(new_n910), .B2(new_n911), .ZN(G1352gat));
  AND3_X1   g711(.A1(new_n904), .A2(new_n906), .A3(KEYINPUT126), .ZN(new_n913));
  AOI21_X1  g712(.A(KEYINPUT126), .B1(new_n904), .B2(new_n906), .ZN(new_n914));
  OAI211_X1 g713(.A(new_n630), .B(new_n909), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT127), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n908), .A2(KEYINPUT127), .A3(new_n630), .A4(new_n909), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n917), .A2(G204gat), .A3(new_n918), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n704), .A2(G204gat), .ZN(new_n920));
  NAND4_X1  g719(.A1(new_n881), .A2(new_n899), .A3(new_n882), .A4(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT62), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n921), .B(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n919), .A2(new_n923), .ZN(G1353gat));
  NAND2_X1  g723(.A1(new_n909), .A2(new_n294), .ZN(new_n925));
  OAI21_X1  g724(.A(G211gat), .B1(new_n859), .B2(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT63), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n926), .B(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(G211gat), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n900), .A2(new_n929), .A3(new_n294), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(new_n930), .ZN(G1354gat));
  AOI21_X1  g730(.A(G218gat), .B1(new_n900), .B2(new_n664), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n256), .A2(G218gat), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n932), .B1(new_n910), .B2(new_n933), .ZN(G1355gat));
endmodule


