//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 1 0 1 1 0 0 0 1 0 0 1 0 1 0 1 1 1 0 0 0 1 0 0 1 1 1 1 1 0 1 0 0 1 1 1 1 0 1 0 0 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n755, new_n757, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n851, new_n852, new_n853, new_n854, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n958, new_n959, new_n960,
    new_n961, new_n962;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G64gat), .B(G92gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G197gat), .B(G204gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT22), .ZN(new_n207));
  XOR2_X1   g006(.A(G211gat), .B(G218gat), .Z(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G211gat), .ZN(new_n210));
  INV_X1    g009(.A(G218gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n210), .A2(new_n211), .A3(KEYINPUT22), .ZN(new_n212));
  NAND2_X1  g011(.A1(G211gat), .A2(G218gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AND3_X1   g013(.A1(new_n214), .A2(KEYINPUT74), .A3(new_n206), .ZN(new_n215));
  AOI21_X1  g014(.A(KEYINPUT74), .B1(new_n214), .B2(new_n206), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n209), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G226gat), .ZN(new_n218));
  INV_X1    g017(.A(G233gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT68), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT27), .ZN(new_n222));
  INV_X1    g021(.A(G183gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n225));
  AOI21_X1  g024(.A(G190gat), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n221), .B1(new_n226), .B2(KEYINPUT28), .ZN(new_n227));
  INV_X1    g026(.A(G190gat), .ZN(new_n228));
  AND2_X1   g027(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n228), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT28), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n231), .A2(KEYINPUT68), .A3(new_n232), .ZN(new_n233));
  OAI211_X1 g032(.A(KEYINPUT28), .B(new_n228), .C1(new_n229), .C2(new_n230), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT69), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(KEYINPUT27), .B(G183gat), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n237), .A2(KEYINPUT69), .A3(KEYINPUT28), .A4(new_n228), .ZN(new_n238));
  AOI22_X1  g037(.A1(new_n227), .A2(new_n233), .B1(new_n236), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(G183gat), .A2(G190gat), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(G169gat), .A2(G176gat), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT66), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n242), .B(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(G169gat), .ZN(new_n245));
  INV_X1    g044(.A(G176gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  OR2_X1    g046(.A1(new_n247), .A2(KEYINPUT26), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(KEYINPUT26), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n244), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  NOR3_X1   g050(.A1(new_n239), .A2(new_n241), .A3(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT25), .ZN(new_n253));
  AND2_X1   g052(.A1(new_n244), .A2(new_n253), .ZN(new_n254));
  AND2_X1   g053(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n255));
  NOR2_X1   g054(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n247), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NOR2_X1   g056(.A1(G169gat), .A2(G176gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(KEYINPUT23), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT64), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n259), .A2(KEYINPUT64), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT24), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n240), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g064(.A1(G183gat), .A2(G190gat), .ZN(new_n266));
  AOI21_X1  g065(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n267));
  NOR3_X1   g066(.A1(new_n265), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n254), .A2(new_n262), .A3(new_n263), .A4(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT67), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n240), .A2(new_n271), .A3(new_n264), .ZN(new_n272));
  INV_X1    g071(.A(new_n266), .ZN(new_n273));
  AOI21_X1  g072(.A(KEYINPUT67), .B1(G183gat), .B2(G190gat), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n272), .B(new_n273), .C1(new_n264), .C2(new_n274), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n275), .A2(new_n244), .A3(new_n257), .A4(new_n259), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT25), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n270), .A2(new_n277), .ZN(new_n278));
  NOR3_X1   g077(.A1(new_n252), .A2(new_n278), .A3(KEYINPUT76), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT76), .ZN(new_n280));
  AND2_X1   g079(.A1(new_n227), .A2(new_n233), .ZN(new_n281));
  AND2_X1   g080(.A1(new_n236), .A2(new_n238), .ZN(new_n282));
  OAI211_X1 g081(.A(new_n240), .B(new_n250), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(KEYINPUT64), .B1(new_n257), .B2(new_n259), .ZN(new_n284));
  INV_X1    g083(.A(new_n263), .ZN(new_n285));
  NOR3_X1   g084(.A1(new_n284), .A2(new_n285), .A3(new_n268), .ZN(new_n286));
  AOI22_X1  g085(.A1(new_n286), .A2(new_n254), .B1(KEYINPUT25), .B2(new_n276), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n280), .B1(new_n283), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n220), .B1(new_n279), .B2(new_n288), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n220), .A2(KEYINPUT29), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT75), .ZN(new_n291));
  NOR3_X1   g090(.A1(new_n252), .A2(new_n278), .A3(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(KEYINPUT75), .B1(new_n283), .B2(new_n287), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n290), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n217), .B1(new_n289), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n291), .B1(new_n252), .B2(new_n278), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n283), .A2(new_n287), .A3(KEYINPUT75), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n296), .A2(new_n220), .A3(new_n297), .ZN(new_n298));
  OAI21_X1  g097(.A(KEYINPUT76), .B1(new_n252), .B2(new_n278), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n283), .A2(new_n287), .A3(new_n280), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n299), .A2(new_n300), .A3(new_n290), .ZN(new_n301));
  AND3_X1   g100(.A1(new_n298), .A2(new_n301), .A3(new_n217), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n205), .B1(new_n295), .B2(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n298), .A2(new_n301), .A3(new_n217), .ZN(new_n304));
  INV_X1    g103(.A(new_n220), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n305), .B1(new_n299), .B2(new_n300), .ZN(new_n306));
  INV_X1    g105(.A(new_n290), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n307), .B1(new_n296), .B2(new_n297), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  OAI211_X1 g108(.A(new_n304), .B(new_n204), .C1(new_n309), .C2(new_n217), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n303), .A2(KEYINPUT30), .A3(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT30), .ZN(new_n312));
  OAI211_X1 g111(.A(new_n312), .B(new_n205), .C1(new_n295), .C2(new_n302), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(G1gat), .B(G29gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n316), .B(G85gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(KEYINPUT0), .B(G57gat), .ZN(new_n318));
  XOR2_X1   g117(.A(new_n317), .B(new_n318), .Z(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(G127gat), .B(G134gat), .ZN(new_n321));
  INV_X1    g120(.A(G120gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(G113gat), .ZN(new_n323));
  INV_X1    g122(.A(G113gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(G120gat), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT1), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT70), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  AOI211_X1 g127(.A(KEYINPUT70), .B(KEYINPUT1), .C1(new_n323), .C2(new_n325), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n321), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n326), .A2(new_n327), .ZN(new_n331));
  INV_X1    g130(.A(new_n321), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  AND2_X1   g133(.A1(KEYINPUT78), .A2(G141gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(KEYINPUT78), .A2(G141gat), .ZN(new_n336));
  OAI21_X1  g135(.A(G148gat), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  AND2_X1   g136(.A1(KEYINPUT79), .A2(G148gat), .ZN(new_n338));
  NOR2_X1   g137(.A1(KEYINPUT79), .A2(G148gat), .ZN(new_n339));
  OAI21_X1  g138(.A(G141gat), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(G155gat), .A2(G162gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT2), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT80), .ZN(new_n344));
  AND2_X1   g143(.A1(G155gat), .A2(G162gat), .ZN(new_n345));
  NOR2_X1   g144(.A1(G155gat), .A2(G162gat), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n344), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(G155gat), .ZN(new_n348));
  INV_X1    g147(.A(G162gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n350), .A2(KEYINPUT80), .A3(new_n342), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n341), .A2(new_n343), .A3(new_n347), .A4(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n346), .B(KEYINPUT77), .ZN(new_n353));
  INV_X1    g152(.A(G141gat), .ZN(new_n354));
  INV_X1    g153(.A(G148gat), .ZN(new_n355));
  AOI21_X1  g154(.A(KEYINPUT2), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(G141gat), .A2(G148gat), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n345), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n353), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(KEYINPUT81), .B(KEYINPUT3), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n352), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT3), .ZN(new_n362));
  AOI22_X1  g161(.A1(new_n337), .A2(new_n340), .B1(KEYINPUT2), .B2(new_n342), .ZN(new_n363));
  AND2_X1   g162(.A1(new_n347), .A2(new_n351), .ZN(new_n364));
  AOI22_X1  g163(.A1(new_n363), .A2(new_n364), .B1(new_n358), .B2(new_n353), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n334), .B(new_n361), .C1(new_n362), .C2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT4), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n352), .A2(new_n359), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n367), .B1(new_n334), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(G225gat), .A2(G233gat), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n371), .B1(new_n334), .B2(new_n368), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n329), .A2(new_n321), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT1), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n324), .A2(G120gat), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n322), .A2(G113gat), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n374), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(KEYINPUT70), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(new_n331), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n373), .B1(new_n379), .B2(new_n321), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n380), .A2(KEYINPUT4), .A3(new_n365), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n366), .A2(new_n369), .A3(new_n372), .A4(new_n381), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n334), .A2(new_n368), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n365), .B1(new_n330), .B2(new_n333), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n371), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n382), .A2(KEYINPUT5), .A3(new_n385), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n371), .A2(KEYINPUT5), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n366), .A2(new_n369), .A3(new_n381), .A4(new_n387), .ZN(new_n388));
  AND3_X1   g187(.A1(new_n386), .A2(KEYINPUT86), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT86), .B1(new_n386), .B2(new_n388), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n320), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n366), .A2(new_n369), .A3(new_n381), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(new_n371), .ZN(new_n393));
  OR3_X1    g192(.A1(new_n383), .A2(new_n384), .A3(new_n371), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n393), .A2(new_n394), .A3(KEYINPUT39), .ZN(new_n395));
  OAI211_X1 g194(.A(new_n395), .B(new_n319), .C1(KEYINPUT39), .C2(new_n393), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n396), .B(KEYINPUT40), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n315), .A2(new_n391), .A3(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT85), .ZN(new_n399));
  AOI21_X1  g198(.A(KEYINPUT29), .B1(new_n365), .B2(new_n360), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n400), .A2(new_n217), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n368), .A2(KEYINPUT3), .ZN(new_n403));
  NAND2_X1  g202(.A1(G228gat), .A2(G233gat), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT29), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n368), .A2(new_n406), .A3(new_n217), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n402), .A2(new_n403), .A3(new_n405), .A4(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n360), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n368), .A2(new_n409), .ZN(new_n410));
  AND3_X1   g209(.A1(new_n407), .A2(KEYINPUT84), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT84), .B1(new_n407), .B2(new_n410), .ZN(new_n412));
  NOR3_X1   g211(.A1(new_n411), .A2(new_n412), .A3(new_n401), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n408), .B1(new_n413), .B2(new_n405), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n399), .B1(new_n414), .B2(G22gat), .ZN(new_n415));
  XOR2_X1   g214(.A(G78gat), .B(G106gat), .Z(new_n416));
  XNOR2_X1  g215(.A(new_n416), .B(KEYINPUT31), .ZN(new_n417));
  INV_X1    g216(.A(G50gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n417), .B(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n414), .A2(G22gat), .ZN(new_n421));
  INV_X1    g220(.A(G22gat), .ZN(new_n422));
  INV_X1    g221(.A(new_n412), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n407), .A2(KEYINPUT84), .A3(new_n410), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n423), .A2(new_n402), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(new_n404), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n422), .B1(new_n426), .B2(new_n408), .ZN(new_n427));
  OAI22_X1  g226(.A1(new_n415), .A2(new_n420), .B1(new_n421), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n414), .A2(G22gat), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n426), .A2(new_n422), .A3(new_n408), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n429), .A2(new_n430), .A3(new_n399), .A4(new_n419), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  XOR2_X1   g231(.A(KEYINPUT87), .B(KEYINPUT37), .Z(new_n433));
  OAI21_X1  g232(.A(new_n433), .B1(new_n295), .B2(new_n302), .ZN(new_n434));
  OAI211_X1 g233(.A(KEYINPUT37), .B(new_n304), .C1(new_n309), .C2(new_n217), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n434), .A2(new_n204), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT38), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n309), .A2(new_n217), .ZN(new_n438));
  AND2_X1   g237(.A1(new_n298), .A2(new_n301), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n438), .B(KEYINPUT37), .C1(new_n217), .C2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT38), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n440), .A2(new_n441), .A3(new_n204), .A4(new_n434), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n386), .A2(new_n388), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(new_n320), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT6), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n386), .A2(new_n319), .A3(new_n388), .ZN(new_n447));
  AND2_X1   g246(.A1(new_n447), .A2(new_n445), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n446), .B1(new_n391), .B2(new_n448), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n437), .A2(new_n442), .A3(new_n449), .A4(new_n303), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n398), .A2(new_n432), .A3(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT88), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n398), .A2(KEYINPUT88), .A3(new_n450), .A4(new_n432), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n444), .A2(KEYINPUT82), .A3(new_n445), .A4(new_n447), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT82), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n443), .B(new_n320), .C1(new_n457), .C2(KEYINPUT6), .ZN(new_n458));
  AOI221_X4 g257(.A(KEYINPUT83), .B1(new_n456), .B2(new_n458), .C1(new_n311), .C2(new_n313), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT83), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n456), .A2(new_n458), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n460), .B1(new_n314), .B2(new_n461), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n432), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n380), .B1(new_n252), .B2(new_n278), .ZN(new_n467));
  AND2_X1   g266(.A1(G227gat), .A2(G233gat), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n283), .A2(new_n287), .A3(new_n334), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT71), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT71), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n467), .A2(new_n469), .A3(new_n472), .A4(new_n468), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT32), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT33), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(G15gat), .B(G43gat), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n478), .B(G99gat), .ZN(new_n479));
  XNOR2_X1  g278(.A(KEYINPUT72), .B(G71gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n479), .B(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n477), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n475), .B1(new_n481), .B2(KEYINPUT33), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n474), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT73), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT73), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n474), .A2(new_n486), .A3(new_n483), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n482), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  AND2_X1   g287(.A1(new_n467), .A2(new_n469), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n489), .A2(new_n468), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT34), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NOR3_X1   g291(.A1(new_n489), .A2(KEYINPUT34), .A3(new_n468), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n488), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n494), .A2(new_n482), .A3(new_n485), .A4(new_n487), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT36), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n496), .A2(KEYINPUT36), .A3(new_n497), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n455), .A2(new_n466), .A3(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n496), .A2(new_n432), .A3(new_n497), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(KEYINPUT90), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT90), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n496), .A2(new_n432), .A3(new_n506), .A4(new_n497), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n463), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT35), .ZN(new_n509));
  AND3_X1   g308(.A1(new_n496), .A2(KEYINPUT89), .A3(new_n497), .ZN(new_n510));
  AOI21_X1  g309(.A(KEYINPUT89), .B1(new_n496), .B2(new_n497), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT35), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n314), .A2(new_n513), .ZN(new_n514));
  NOR3_X1   g313(.A1(new_n465), .A2(new_n514), .A3(new_n449), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n509), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n503), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(KEYINPUT99), .B(G92gat), .ZN(new_n519));
  INV_X1    g318(.A(G85gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(G99gat), .A2(G106gat), .ZN(new_n521));
  AOI22_X1  g320(.A1(new_n519), .A2(new_n520), .B1(KEYINPUT8), .B2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT98), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n523), .A2(G85gat), .A3(G92gat), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT7), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OR2_X1    g325(.A1(new_n524), .A2(new_n525), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n522), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(G99gat), .B(G106gat), .ZN(new_n529));
  OR2_X1    g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n528), .A2(new_n529), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT100), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n532), .B(new_n533), .ZN(new_n534));
  XOR2_X1   g333(.A(G43gat), .B(G50gat), .Z(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT15), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT15), .ZN(new_n538));
  AOI22_X1  g337(.A1(new_n535), .A2(new_n538), .B1(G29gat), .B2(G36gat), .ZN(new_n539));
  NOR3_X1   g338(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(KEYINPUT92), .ZN(new_n541));
  OAI21_X1  g340(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  OAI211_X1 g342(.A(new_n537), .B(new_n539), .C1(new_n541), .C2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(G29gat), .A2(G36gat), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n545), .B1(new_n543), .B2(new_n540), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n536), .A2(new_n546), .A3(KEYINPUT15), .ZN(new_n547));
  AOI21_X1  g346(.A(KEYINPUT93), .B1(new_n544), .B2(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT17), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n534), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n544), .A2(new_n547), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n532), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n550), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(G134gat), .B(G162gat), .ZN(new_n555));
  XOR2_X1   g354(.A(new_n555), .B(KEYINPUT101), .Z(new_n556));
  NAND2_X1  g355(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  XOR2_X1   g356(.A(G190gat), .B(G218gat), .Z(new_n558));
  AOI21_X1  g357(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n556), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n550), .A2(new_n561), .A3(new_n551), .A4(new_n553), .ZN(new_n562));
  AND3_X1   g361(.A1(new_n557), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n560), .B1(new_n557), .B2(new_n562), .ZN(new_n564));
  OR2_X1    g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G127gat), .B(G155gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(G211gat), .ZN(new_n567));
  XOR2_X1   g366(.A(G15gat), .B(G22gat), .Z(new_n568));
  INV_X1    g367(.A(G1gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G15gat), .B(G22gat), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT16), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n571), .B1(new_n572), .B2(G1gat), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n570), .A2(new_n573), .A3(KEYINPUT94), .ZN(new_n574));
  INV_X1    g373(.A(G8gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT21), .ZN(new_n577));
  XNOR2_X1  g376(.A(G57gat), .B(G64gat), .ZN(new_n578));
  OR2_X1    g377(.A1(new_n578), .A2(KEYINPUT96), .ZN(new_n579));
  NAND2_X1  g378(.A1(G71gat), .A2(G78gat), .ZN(new_n580));
  OR2_X1    g379(.A1(G71gat), .A2(G78gat), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT9), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n578), .A2(KEYINPUT96), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n579), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  OAI211_X1 g384(.A(new_n580), .B(new_n581), .C1(new_n578), .C2(new_n582), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  OAI211_X1 g386(.A(new_n576), .B(new_n223), .C1(new_n577), .C2(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n574), .B(G8gat), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n587), .A2(new_n577), .ZN(new_n590));
  OAI21_X1  g389(.A(G183gat), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(G231gat), .A2(G233gat), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n592), .A2(new_n593), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n567), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n596), .ZN(new_n598));
  INV_X1    g397(.A(new_n567), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n598), .A2(new_n594), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n587), .A2(new_n577), .ZN(new_n601));
  XNOR2_X1  g400(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT97), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n601), .B(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n597), .A2(new_n600), .A3(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n604), .B1(new_n597), .B2(new_n600), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n565), .A2(new_n608), .A3(KEYINPUT102), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT102), .ZN(new_n610));
  INV_X1    g409(.A(new_n607), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(new_n605), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n563), .A2(new_n564), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n610), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  AND2_X1   g413(.A1(new_n609), .A2(new_n614), .ZN(new_n615));
  AND2_X1   g414(.A1(new_n518), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n587), .ZN(new_n617));
  OAI21_X1  g416(.A(KEYINPUT103), .B1(new_n532), .B2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT103), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n530), .A2(new_n619), .A3(new_n587), .A4(new_n531), .ZN(new_n620));
  INV_X1    g419(.A(new_n529), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(KEYINPUT104), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n528), .B(new_n622), .ZN(new_n623));
  AOI22_X1  g422(.A1(new_n618), .A2(new_n620), .B1(new_n617), .B2(new_n623), .ZN(new_n624));
  XOR2_X1   g423(.A(KEYINPUT105), .B(KEYINPUT10), .Z(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n532), .A2(KEYINPUT10), .A3(new_n617), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT106), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(G230gat), .A2(G233gat), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n626), .A2(KEYINPUT106), .A3(new_n627), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT107), .ZN(new_n634));
  OR3_X1    g433(.A1(new_n624), .A2(new_n634), .A3(new_n631), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n634), .B1(new_n624), .B2(new_n631), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(G120gat), .B(G148gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(G176gat), .B(G204gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n633), .A2(new_n638), .A3(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n631), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n644), .B1(new_n626), .B2(new_n627), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n641), .B1(new_n637), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(KEYINPUT108), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT108), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n643), .A2(new_n649), .A3(new_n646), .ZN(new_n650));
  AND2_X1   g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n549), .A2(new_n576), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n589), .A2(new_n552), .ZN(new_n653));
  AND2_X1   g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(G229gat), .A2(G233gat), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n654), .A2(KEYINPUT18), .A3(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n589), .A2(new_n552), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n657), .B(KEYINPUT95), .Z(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(new_n653), .ZN(new_n659));
  XOR2_X1   g458(.A(new_n655), .B(KEYINPUT13), .Z(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n652), .A2(new_n655), .A3(new_n653), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT18), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n656), .A2(new_n661), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(G169gat), .B(G197gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT91), .B(KEYINPUT11), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(G113gat), .B(G141gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT12), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n665), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n656), .A2(new_n661), .A3(new_n671), .A4(new_n664), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n651), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n616), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n678), .A2(new_n461), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(new_n569), .ZN(G1324gat));
  INV_X1    g479(.A(new_n678), .ZN(new_n681));
  NAND2_X1  g480(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n572), .A2(new_n575), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n681), .A2(new_n315), .A3(new_n682), .A4(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT42), .ZN(new_n685));
  OR2_X1    g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(G8gat), .B1(new_n678), .B2(new_n314), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n684), .A2(new_n685), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(G1325gat));
  INV_X1    g488(.A(new_n502), .ZN(new_n690));
  AND3_X1   g489(.A1(new_n681), .A2(G15gat), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(G15gat), .B1(new_n681), .B2(new_n512), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n691), .A2(new_n692), .ZN(G1326gat));
  NOR2_X1   g492(.A1(new_n678), .A2(new_n432), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(new_n422), .ZN(new_n695));
  XNOR2_X1  g494(.A(KEYINPUT109), .B(KEYINPUT43), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(G1327gat));
  NAND2_X1  g496(.A1(new_n518), .A2(new_n613), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n677), .A2(new_n612), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n701), .A2(G29gat), .A3(new_n461), .ZN(new_n702));
  XOR2_X1   g501(.A(new_n702), .B(KEYINPUT45), .Z(new_n703));
  INV_X1    g502(.A(KEYINPUT112), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT110), .ZN(new_n705));
  AOI221_X4 g504(.A(new_n705), .B1(new_n512), .B2(new_n515), .C1(new_n508), .C2(KEYINPUT35), .ZN(new_n706));
  AOI21_X1  g505(.A(KEYINPUT110), .B1(new_n509), .B2(new_n516), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n503), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(KEYINPUT111), .B(KEYINPUT44), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n708), .A2(new_n613), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n698), .A2(KEYINPUT44), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n699), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n704), .B1(new_n714), .B2(new_n461), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n699), .B1(new_n710), .B2(new_n711), .ZN(new_n716));
  INV_X1    g515(.A(new_n461), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n716), .A2(KEYINPUT112), .A3(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n715), .A2(G29gat), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n719), .ZN(G1328gat));
  NOR3_X1   g519(.A1(new_n701), .A2(G36gat), .A3(new_n314), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT46), .ZN(new_n722));
  OAI21_X1  g521(.A(G36gat), .B1(new_n714), .B2(new_n314), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(G1329gat));
  OAI21_X1  g523(.A(G43gat), .B1(new_n714), .B2(new_n502), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n565), .B1(new_n503), .B2(new_n517), .ZN(new_n726));
  INV_X1    g525(.A(G43gat), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n726), .A2(new_n727), .A3(new_n512), .A4(new_n713), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n725), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT113), .ZN(new_n730));
  AOI21_X1  g529(.A(KEYINPUT47), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT114), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n729), .B(new_n732), .ZN(G1330gat));
  NAND3_X1  g532(.A1(new_n716), .A2(G50gat), .A3(new_n465), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n418), .B1(new_n701), .B2(new_n432), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT48), .ZN(new_n736));
  OAI211_X1 g535(.A(new_n734), .B(new_n735), .C1(KEYINPUT115), .C2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(KEYINPUT115), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n737), .B(new_n738), .ZN(G1331gat));
  AND2_X1   g538(.A1(new_n708), .A2(new_n651), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n609), .A2(new_n614), .A3(new_n676), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n717), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g544(.A1(new_n740), .A2(new_n742), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n746), .A2(new_n314), .ZN(new_n747));
  NOR2_X1   g546(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n748));
  AND2_X1   g547(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n750), .B1(new_n747), .B2(new_n748), .ZN(G1333gat));
  NAND3_X1  g550(.A1(new_n743), .A2(G71gat), .A3(new_n690), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n512), .B(KEYINPUT116), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n746), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n752), .B1(G71gat), .B2(new_n754), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g555(.A1(new_n743), .A2(new_n465), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g557(.A1(new_n648), .A2(new_n650), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n675), .A2(new_n608), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n708), .A2(new_n613), .A3(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT51), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n708), .A2(KEYINPUT51), .A3(new_n613), .A4(new_n760), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n759), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(G85gat), .B1(new_n765), .B2(new_n717), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n712), .A2(new_n651), .A3(new_n760), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n767), .A2(new_n520), .A3(new_n461), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n766), .A2(new_n768), .ZN(G1336gat));
  INV_X1    g568(.A(new_n519), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n770), .B1(new_n767), .B2(new_n314), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT52), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n763), .A2(new_n764), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  OR3_X1    g573(.A1(new_n759), .A2(G92gat), .A3(new_n314), .ZN(new_n775));
  OAI211_X1 g574(.A(new_n771), .B(new_n772), .C1(new_n774), .C2(new_n775), .ZN(new_n776));
  XOR2_X1   g575(.A(new_n775), .B(KEYINPUT117), .Z(new_n777));
  NAND2_X1  g576(.A1(new_n773), .A2(new_n777), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n771), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n776), .B1(new_n779), .B2(new_n772), .ZN(G1337gat));
  AOI21_X1  g579(.A(G99gat), .B1(new_n765), .B2(new_n512), .ZN(new_n781));
  INV_X1    g580(.A(G99gat), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n767), .A2(new_n782), .A3(new_n502), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n781), .A2(new_n783), .ZN(G1338gat));
  INV_X1    g583(.A(KEYINPUT53), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n785), .A2(KEYINPUT118), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n773), .A2(new_n651), .A3(new_n465), .ZN(new_n788));
  INV_X1    g587(.A(G106gat), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n432), .A2(new_n789), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n712), .A2(new_n651), .A3(new_n760), .A4(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n785), .A2(KEYINPUT118), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n787), .B1(new_n790), .B2(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(G106gat), .B1(new_n765), .B2(new_n465), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n792), .A2(new_n793), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n796), .A2(new_n797), .A3(new_n786), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n795), .A2(new_n798), .ZN(G1339gat));
  INV_X1    g598(.A(KEYINPUT119), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n800), .B1(new_n651), .B2(new_n741), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n615), .A2(KEYINPUT119), .A3(new_n676), .A4(new_n759), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n804));
  OAI21_X1  g603(.A(KEYINPUT54), .B1(new_n628), .B2(new_n631), .ZN(new_n805));
  AOI21_X1  g604(.A(KEYINPUT106), .B1(new_n626), .B2(new_n627), .ZN(new_n806));
  INV_X1    g605(.A(new_n627), .ZN(new_n807));
  AOI211_X1 g606(.A(new_n629), .B(new_n807), .C1(new_n624), .C2(new_n625), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n805), .B1(new_n809), .B2(new_n631), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT54), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n642), .B1(new_n645), .B2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n804), .B1(new_n810), .B2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(new_n633), .ZN(new_n815));
  OAI211_X1 g614(.A(KEYINPUT55), .B(new_n812), .C1(new_n815), .C2(new_n805), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n659), .A2(new_n660), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n654), .A2(new_n655), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n670), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n820), .A2(new_n674), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n817), .A2(new_n643), .A3(new_n613), .A4(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n648), .A2(new_n650), .A3(new_n821), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n814), .A2(new_n816), .A3(new_n675), .A4(new_n643), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT120), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n823), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n565), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n825), .B1(new_n823), .B2(new_n824), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n822), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n803), .B1(new_n829), .B2(new_n612), .ZN(new_n830));
  OAI21_X1  g629(.A(KEYINPUT121), .B1(new_n830), .B2(new_n465), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT121), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n823), .A2(new_n824), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(KEYINPUT120), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n834), .A2(new_n565), .A3(new_n826), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n608), .B1(new_n835), .B2(new_n822), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n832), .B(new_n432), .C1(new_n836), .C2(new_n803), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n831), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n315), .A2(new_n461), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n838), .A2(new_n512), .A3(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(G113gat), .B1(new_n840), .B2(new_n676), .ZN(new_n841));
  INV_X1    g640(.A(new_n830), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n505), .A2(new_n507), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n842), .A2(new_n843), .A3(new_n839), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n845), .A2(new_n324), .A3(new_n675), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n841), .A2(new_n846), .ZN(G1340gat));
  OAI21_X1  g646(.A(G120gat), .B1(new_n840), .B2(new_n759), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n845), .A2(new_n322), .A3(new_n651), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(G1341gat));
  NAND2_X1  g649(.A1(new_n608), .A2(G127gat), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n844), .A2(new_n612), .ZN(new_n852));
  OAI22_X1  g651(.A1(new_n840), .A2(new_n851), .B1(new_n852), .B2(G127gat), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT122), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n853), .B(new_n854), .ZN(G1342gat));
  AND2_X1   g654(.A1(new_n842), .A2(new_n843), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n613), .A2(new_n314), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n857), .A2(G134gat), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n856), .A2(new_n717), .A3(new_n858), .ZN(new_n859));
  XOR2_X1   g658(.A(new_n859), .B(KEYINPUT56), .Z(new_n860));
  OAI21_X1  g659(.A(G134gat), .B1(new_n840), .B2(new_n565), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(G1343gat));
  NOR2_X1   g661(.A1(new_n335), .A2(new_n336), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n830), .A2(new_n432), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT57), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n502), .A2(new_n839), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n833), .A2(new_n565), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n608), .B1(new_n868), .B2(new_n822), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n465), .B1(new_n803), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n867), .B1(new_n870), .B2(KEYINPUT57), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n866), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n863), .B1(new_n872), .B2(new_n676), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n830), .A2(new_n432), .A3(new_n690), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(new_n839), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n675), .A2(new_n354), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n873), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(KEYINPUT58), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT58), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n873), .B(new_n879), .C1(new_n875), .C2(new_n876), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n878), .A2(new_n880), .ZN(G1344gat));
  INV_X1    g680(.A(new_n875), .ZN(new_n882));
  OR2_X1    g681(.A1(new_n338), .A2(new_n339), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n882), .A2(new_n883), .A3(new_n651), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT59), .ZN(new_n885));
  OAI21_X1  g684(.A(KEYINPUT57), .B1(new_n830), .B2(new_n432), .ZN(new_n886));
  INV_X1    g685(.A(new_n867), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n651), .A2(new_n741), .ZN(new_n888));
  OAI211_X1 g687(.A(new_n865), .B(new_n465), .C1(new_n869), .C2(new_n888), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n886), .A2(new_n651), .A3(new_n887), .A4(new_n889), .ZN(new_n890));
  OR2_X1    g689(.A1(new_n890), .A2(KEYINPUT123), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n355), .B1(new_n890), .B2(KEYINPUT123), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n885), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n885), .B1(new_n872), .B2(new_n759), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n894), .A2(new_n883), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n884), .B1(new_n893), .B2(new_n895), .ZN(G1345gat));
  AOI21_X1  g695(.A(G155gat), .B1(new_n882), .B2(new_n608), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n872), .A2(new_n348), .A3(new_n612), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n897), .A2(new_n898), .ZN(G1346gat));
  OR3_X1    g698(.A1(new_n872), .A2(KEYINPUT124), .A3(new_n565), .ZN(new_n900));
  OAI21_X1  g699(.A(KEYINPUT124), .B1(new_n872), .B2(new_n565), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n900), .A2(G162gat), .A3(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n874), .A2(new_n349), .A3(new_n717), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n902), .B1(new_n857), .B2(new_n903), .ZN(G1347gat));
  NOR2_X1   g703(.A1(new_n717), .A2(new_n314), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n856), .A2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n907), .A2(new_n245), .A3(new_n675), .ZN(new_n908));
  INV_X1    g707(.A(new_n905), .ZN(new_n909));
  AOI211_X1 g708(.A(new_n753), .B(new_n909), .C1(new_n831), .C2(new_n837), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n910), .A2(new_n675), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n908), .B1(new_n911), .B2(new_n245), .ZN(G1348gat));
  NAND3_X1  g711(.A1(new_n910), .A2(G176gat), .A3(new_n651), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT125), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n910), .A2(KEYINPUT125), .A3(G176gat), .A4(new_n651), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n246), .B1(new_n906), .B2(new_n759), .ZN(new_n917));
  AND3_X1   g716(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(G1349gat));
  INV_X1    g717(.A(new_n753), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n838), .A2(new_n919), .A3(new_n905), .ZN(new_n920));
  OAI21_X1  g719(.A(G183gat), .B1(new_n920), .B2(new_n612), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT60), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n608), .A2(new_n237), .ZN(new_n923));
  OAI211_X1 g722(.A(new_n921), .B(new_n922), .C1(new_n906), .C2(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n223), .B1(new_n910), .B2(new_n608), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n906), .A2(new_n923), .ZN(new_n926));
  OAI21_X1  g725(.A(KEYINPUT60), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n924), .A2(new_n927), .ZN(G1350gat));
  NAND3_X1  g727(.A1(new_n907), .A2(new_n228), .A3(new_n613), .ZN(new_n929));
  NAND4_X1  g728(.A1(new_n838), .A2(new_n613), .A3(new_n919), .A4(new_n905), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT61), .ZN(new_n931));
  AND3_X1   g730(.A1(new_n930), .A2(new_n931), .A3(G190gat), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n931), .B1(new_n930), .B2(G190gat), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n929), .B1(new_n932), .B2(new_n933), .ZN(G1351gat));
  NOR2_X1   g733(.A1(new_n690), .A2(new_n909), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n864), .A2(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(G197gat), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n936), .A2(new_n937), .A3(new_n675), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n886), .A2(new_n889), .ZN(new_n939));
  AND3_X1   g738(.A1(new_n939), .A2(new_n675), .A3(new_n935), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n938), .B1(new_n940), .B2(new_n937), .ZN(G1352gat));
  INV_X1    g740(.A(G204gat), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n936), .A2(new_n942), .A3(new_n651), .ZN(new_n943));
  OR2_X1    g742(.A1(new_n943), .A2(KEYINPUT62), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(KEYINPUT62), .ZN(new_n945));
  AND3_X1   g744(.A1(new_n939), .A2(new_n651), .A3(new_n935), .ZN(new_n946));
  OAI211_X1 g745(.A(new_n944), .B(new_n945), .C1(new_n942), .C2(new_n946), .ZN(G1353gat));
  NAND3_X1  g746(.A1(new_n939), .A2(new_n608), .A3(new_n935), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(G211gat), .ZN(new_n949));
  NAND2_X1  g748(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT126), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT63), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n949), .A2(new_n950), .A3(new_n953), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n936), .A2(new_n210), .A3(new_n608), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n948), .A2(new_n951), .A3(new_n952), .A4(G211gat), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n954), .A2(new_n955), .A3(new_n956), .ZN(G1354gat));
  NAND3_X1  g756(.A1(new_n936), .A2(new_n211), .A3(new_n613), .ZN(new_n958));
  NAND4_X1  g757(.A1(new_n886), .A2(new_n613), .A3(new_n889), .A4(new_n935), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(G218gat), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT127), .ZN(new_n962));
  XNOR2_X1  g761(.A(new_n961), .B(new_n962), .ZN(G1355gat));
endmodule


