//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 1 0 0 1 1 1 1 1 0 0 1 1 1 1 0 0 0 0 1 0 1 1 0 0 0 0 0 0 1 1 0 1 1 1 0 0 1 1 0 1 0 0 1 1 0 1 0 0 0 1 1 0 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:23 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n556, new_n558, new_n559,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n623, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1196,
    new_n1197, new_n1198;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT66), .ZN(new_n460));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  AOI22_X1  g036(.A1(new_n461), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G125), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n465), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n472), .A2(KEYINPUT66), .A3(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n464), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n461), .A2(G137), .A3(new_n463), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n466), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G101), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT67), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n476), .A2(KEYINPUT67), .A3(G101), .ZN(new_n480));
  AND3_X1   g055(.A1(new_n475), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n474), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G160));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n470), .A2(KEYINPUT68), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT68), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n461), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n486), .A2(new_n488), .A3(G2105), .ZN(new_n489));
  INV_X1    g064(.A(G124), .ZN(new_n490));
  INV_X1    g065(.A(G136), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n486), .A2(new_n488), .A3(new_n463), .ZN(new_n492));
  OAI221_X1 g067(.A(new_n485), .B1(new_n489), .B2(new_n490), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  NAND4_X1  g069(.A1(new_n467), .A2(new_n469), .A3(G138), .A4(new_n463), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT71), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n461), .A2(KEYINPUT71), .A3(G138), .A4(new_n463), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n497), .A2(new_n498), .A3(KEYINPUT4), .ZN(new_n499));
  XNOR2_X1  g074(.A(KEYINPUT69), .B(G114), .ZN(new_n500));
  OAI21_X1  g075(.A(KEYINPUT70), .B1(new_n500), .B2(new_n463), .ZN(new_n501));
  OAI21_X1  g076(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT70), .ZN(new_n504));
  INV_X1    g079(.A(G114), .ZN(new_n505));
  AND2_X1   g080(.A1(new_n505), .A2(KEYINPUT69), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(KEYINPUT69), .ZN(new_n507));
  OAI211_X1 g082(.A(new_n504), .B(G2105), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n501), .A2(new_n503), .A3(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT4), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n495), .A2(new_n496), .A3(new_n510), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n461), .A2(G126), .A3(G2105), .ZN(new_n512));
  NAND4_X1  g087(.A1(new_n499), .A2(new_n509), .A3(new_n511), .A4(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(G164));
  XNOR2_X1  g089(.A(KEYINPUT5), .B(G543), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT6), .B(G651), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n515), .A2(new_n516), .A3(G88), .ZN(new_n517));
  AND2_X1   g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  OAI211_X1 g094(.A(G50), .B(G543), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(G75), .A2(G543), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n522), .B1(new_n515), .B2(G62), .ZN(new_n523));
  INV_X1    g098(.A(G651), .ZN(new_n524));
  OAI211_X1 g099(.A(new_n517), .B(new_n520), .C1(new_n523), .C2(new_n524), .ZN(G303));
  INV_X1    g100(.A(G303), .ZN(G166));
  NAND3_X1  g101(.A1(new_n515), .A2(G63), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT72), .ZN(new_n528));
  AND2_X1   g103(.A1(new_n516), .A2(G543), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G51), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT7), .ZN(new_n532));
  INV_X1    g107(.A(G543), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(KEYINPUT5), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT5), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G543), .ZN(new_n536));
  OAI211_X1 g111(.A(new_n534), .B(new_n536), .C1(new_n518), .C2(new_n519), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G89), .ZN(new_n539));
  NAND4_X1  g114(.A1(new_n528), .A2(new_n530), .A3(new_n532), .A4(new_n539), .ZN(G286));
  INV_X1    g115(.A(G286), .ZN(G168));
  AOI22_X1  g116(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(new_n524), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n516), .A2(G543), .ZN(new_n544));
  INV_X1    g119(.A(G52), .ZN(new_n545));
  INV_X1    g120(.A(G90), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n544), .A2(new_n545), .B1(new_n537), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n543), .A2(new_n547), .ZN(G171));
  AOI22_X1  g123(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n549), .A2(new_n524), .ZN(new_n550));
  INV_X1    g125(.A(G43), .ZN(new_n551));
  INV_X1    g126(.A(G81), .ZN(new_n552));
  OAI22_X1  g127(.A1(new_n544), .A2(new_n551), .B1(new_n537), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  AND3_X1   g130(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n556), .A2(new_n559), .ZN(G188));
  NAND3_X1  g135(.A1(new_n529), .A2(KEYINPUT73), .A3(G53), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(KEYINPUT9), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n529), .A2(KEYINPUT73), .A3(new_n563), .A4(G53), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n562), .A2(new_n564), .B1(G91), .B2(new_n538), .ZN(new_n565));
  NAND2_X1  g140(.A1(G78), .A2(G543), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n534), .A2(new_n536), .ZN(new_n567));
  INV_X1    g142(.A(G65), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G651), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT74), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n565), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(KEYINPUT75), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT75), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n565), .A2(new_n571), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n573), .A2(new_n575), .ZN(G299));
  INV_X1    g151(.A(G171), .ZN(G301));
  OAI21_X1  g152(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n515), .A2(new_n516), .A3(G87), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n516), .A2(G49), .A3(G543), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n581), .B(KEYINPUT76), .ZN(G288));
  OAI211_X1 g157(.A(G48), .B(G543), .C1(new_n518), .C2(new_n519), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n534), .A2(new_n536), .A3(G61), .ZN(new_n585));
  NAND2_X1  g160(.A1(G73), .A2(G543), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(KEYINPUT77), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT77), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n588), .A2(G73), .A3(G543), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n585), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n584), .B1(new_n590), .B2(G651), .ZN(new_n591));
  INV_X1    g166(.A(G86), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n537), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n591), .A2(new_n594), .ZN(G305));
  AOI22_X1  g170(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n596), .A2(new_n524), .ZN(new_n597));
  XNOR2_X1  g172(.A(KEYINPUT78), .B(G47), .ZN(new_n598));
  INV_X1    g173(.A(G85), .ZN(new_n599));
  OAI22_X1  g174(.A1(new_n544), .A2(new_n598), .B1(new_n537), .B2(new_n599), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(G290));
  NAND2_X1  g177(.A1(G301), .A2(G868), .ZN(new_n603));
  NAND2_X1  g178(.A1(G79), .A2(G543), .ZN(new_n604));
  INV_X1    g179(.A(G66), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n567), .B2(new_n605), .ZN(new_n606));
  AOI22_X1  g181(.A1(G651), .A2(new_n606), .B1(new_n529), .B2(G54), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT80), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n538), .A2(G92), .ZN(new_n609));
  XOR2_X1   g184(.A(KEYINPUT79), .B(KEYINPUT10), .Z(new_n610));
  XNOR2_X1  g185(.A(new_n609), .B(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n603), .B1(new_n613), .B2(G868), .ZN(G284));
  OAI21_X1  g189(.A(new_n603), .B1(new_n613), .B2(G868), .ZN(G321));
  INV_X1    g190(.A(G299), .ZN(new_n616));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(G168), .A2(G868), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(KEYINPUT81), .Z(G297));
  INV_X1    g196(.A(new_n620), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n613), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n613), .A2(new_n623), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G868), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(G868), .B2(new_n554), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g203(.A(new_n489), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(G123), .ZN(new_n630));
  OAI21_X1  g205(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n631));
  INV_X1    g206(.A(KEYINPUT83), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n632), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n633), .B(new_n634), .C1(G111), .C2(new_n463), .ZN(new_n635));
  AND2_X1   g210(.A1(new_n630), .A2(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(KEYINPUT82), .ZN(new_n637));
  INV_X1    g212(.A(G135), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n637), .B1(new_n492), .B2(new_n638), .ZN(new_n639));
  INV_X1    g214(.A(new_n492), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n640), .A2(KEYINPUT82), .A3(G135), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n636), .A2(new_n639), .A3(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(G2096), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n461), .A2(new_n476), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT12), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT13), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2100), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n644), .A2(new_n648), .ZN(G156));
  XNOR2_X1  g224(.A(KEYINPUT15), .B(G2430), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2435), .ZN(new_n651));
  XOR2_X1   g226(.A(G2427), .B(G2438), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(KEYINPUT14), .ZN(new_n654));
  XOR2_X1   g229(.A(G1341), .B(G1348), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2443), .B(G2446), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2451), .B(G2454), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT16), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT84), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n658), .A2(new_n661), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n662), .A2(G14), .A3(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(KEYINPUT85), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n664), .A2(new_n665), .ZN(new_n667));
  AND2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(G401));
  XNOR2_X1  g243(.A(G2072), .B(G2078), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT17), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2067), .B(G2678), .ZN(new_n671));
  XOR2_X1   g246(.A(G2084), .B(G2090), .Z(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  NOR3_X1   g248(.A1(new_n670), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n673), .B1(new_n671), .B2(new_n669), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(KEYINPUT87), .Z(new_n676));
  NAND2_X1  g251(.A1(new_n670), .A2(new_n671), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n674), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n672), .A2(new_n671), .A3(new_n669), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT86), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT18), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(new_n643), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(G2100), .ZN(G227));
  XNOR2_X1  g259(.A(G1971), .B(G1976), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT88), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT19), .ZN(new_n687));
  XOR2_X1   g262(.A(G1956), .B(G2474), .Z(new_n688));
  XOR2_X1   g263(.A(G1961), .B(G1966), .Z(new_n689));
  AND2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT20), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n688), .A2(new_n689), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n687), .A2(new_n693), .ZN(new_n694));
  OR3_X1    g269(.A1(new_n687), .A2(new_n690), .A3(new_n693), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n692), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT21), .B(G1986), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(G1991), .B(G1996), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT22), .B(G1981), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n700), .B(new_n701), .Z(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(G229));
  INV_X1    g278(.A(G16), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G5), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G171), .B2(new_n704), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(G1961), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT30), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G28), .ZN(new_n709));
  INV_X1    g284(.A(G29), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(new_n708), .B2(G28), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n709), .B1(new_n711), .B2(KEYINPUT101), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(KEYINPUT101), .B2(new_n711), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n707), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT89), .B(G29), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n493), .A2(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(G35), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n716), .B1(new_n717), .B2(new_n715), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(KEYINPUT29), .ZN(new_n719));
  INV_X1    g294(.A(G2090), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT29), .ZN(new_n721));
  OAI211_X1 g296(.A(new_n716), .B(new_n721), .C1(new_n717), .C2(new_n715), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n719), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  OR2_X1    g298(.A1(G104), .A2(G2105), .ZN(new_n724));
  OAI211_X1 g299(.A(new_n724), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT96), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G128), .ZN(new_n728));
  INV_X1    g303(.A(G140), .ZN(new_n729));
  OAI221_X1 g304(.A(new_n727), .B1(new_n489), .B2(new_n728), .C1(new_n729), .C2(new_n492), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G29), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT28), .ZN(new_n732));
  INV_X1    g307(.A(G26), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n732), .B1(new_n715), .B2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(new_n715), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n735), .A2(KEYINPUT28), .A3(G26), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n731), .A2(new_n734), .A3(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(G2067), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND4_X1  g314(.A1(new_n731), .A2(G2067), .A3(new_n734), .A4(new_n736), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT24), .B(G34), .Z(new_n742));
  OAI22_X1  g317(.A1(new_n482), .A2(new_n710), .B1(new_n715), .B2(new_n742), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G2084), .ZN(new_n744));
  AND3_X1   g319(.A1(new_n723), .A2(new_n741), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(KEYINPUT23), .B1(new_n704), .B2(G20), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(G299), .B2(G16), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n704), .A2(KEYINPUT23), .A3(G20), .ZN(new_n748));
  AND3_X1   g323(.A1(new_n747), .A2(G1956), .A3(new_n748), .ZN(new_n749));
  AOI21_X1  g324(.A(G1956), .B1(new_n747), .B2(new_n748), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n714), .B(new_n745), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n640), .A2(G141), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT99), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n476), .A2(G105), .ZN(new_n756));
  NAND3_X1  g331(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT26), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n629), .B2(G129), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n755), .A2(new_n756), .A3(new_n759), .ZN(new_n760));
  MUX2_X1   g335(.A(G32), .B(new_n760), .S(G29), .Z(new_n761));
  XOR2_X1   g336(.A(KEYINPUT27), .B(G1996), .Z(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT100), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n761), .B(new_n763), .Z(new_n764));
  INV_X1    g339(.A(G19), .ZN(new_n765));
  OAI21_X1  g340(.A(KEYINPUT95), .B1(new_n765), .B2(G16), .ZN(new_n766));
  OR3_X1    g341(.A1(new_n765), .A2(KEYINPUT95), .A3(G16), .ZN(new_n767));
  OAI211_X1 g342(.A(new_n766), .B(new_n767), .C1(new_n554), .C2(new_n704), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(G1341), .Z(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT31), .B(G11), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n769), .B(new_n770), .C1(new_n642), .C2(new_n735), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n704), .A2(G21), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G168), .B2(new_n704), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G1966), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n771), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n720), .B1(new_n719), .B2(new_n722), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n476), .A2(G103), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT25), .Z(new_n778));
  INV_X1    g353(.A(G139), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n778), .B1(new_n492), .B2(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT97), .ZN(new_n781));
  AND2_X1   g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n780), .A2(new_n781), .ZN(new_n783));
  AOI22_X1  g358(.A1(new_n461), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n784));
  OAI22_X1  g359(.A1(new_n782), .A2(new_n783), .B1(new_n463), .B2(new_n784), .ZN(new_n785));
  MUX2_X1   g360(.A(G33), .B(new_n785), .S(G29), .Z(new_n786));
  AOI21_X1  g361(.A(new_n776), .B1(new_n786), .B2(G2072), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n752), .A2(new_n764), .A3(new_n775), .A4(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT36), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT94), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT90), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n581), .A2(new_n791), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n578), .A2(new_n579), .A3(new_n580), .A4(KEYINPUT90), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n794), .A2(G16), .ZN(new_n795));
  XOR2_X1   g370(.A(KEYINPUT33), .B(G1976), .Z(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g372(.A1(G16), .A2(G23), .ZN(new_n798));
  INV_X1    g373(.A(new_n798), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n795), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n704), .B1(new_n792), .B2(new_n793), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n796), .B1(new_n801), .B2(new_n798), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT32), .B(G1981), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n704), .B1(new_n591), .B2(new_n594), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n704), .A2(G6), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n804), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(new_n804), .ZN(new_n809));
  AND2_X1   g384(.A1(new_n587), .A2(new_n589), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n524), .B1(new_n810), .B2(new_n585), .ZN(new_n811));
  NOR3_X1   g386(.A1(new_n811), .A2(new_n593), .A3(new_n584), .ZN(new_n812));
  OAI211_X1 g387(.A(new_n809), .B(new_n806), .C1(new_n812), .C2(new_n704), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n808), .A2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n803), .A2(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(G1971), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT92), .ZN(new_n818));
  INV_X1    g393(.A(G22), .ZN(new_n819));
  NOR3_X1   g394(.A1(new_n819), .A2(KEYINPUT91), .A3(G16), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(G303), .B2(G16), .ZN(new_n821));
  OAI21_X1  g396(.A(KEYINPUT91), .B1(new_n819), .B2(G16), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n818), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(G88), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n520), .B1(new_n537), .B2(new_n824), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n534), .A2(new_n536), .A3(G62), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n524), .B1(new_n826), .B2(new_n521), .ZN(new_n827));
  OAI21_X1  g402(.A(G16), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(new_n820), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n828), .A2(new_n818), .A3(new_n822), .A4(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n817), .B1(new_n823), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n828), .A2(new_n822), .A3(new_n829), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(KEYINPUT92), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n834), .A2(G1971), .A3(new_n830), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  NOR3_X1   g411(.A1(new_n816), .A2(new_n836), .A3(KEYINPUT93), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT93), .ZN(new_n838));
  AND3_X1   g413(.A1(new_n834), .A2(G1971), .A3(new_n830), .ZN(new_n839));
  AOI21_X1  g414(.A(G1971), .B1(new_n834), .B2(new_n830), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n814), .B1(new_n802), .B2(new_n800), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n838), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(KEYINPUT34), .B1(new_n837), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(KEYINPUT93), .B1(new_n816), .B2(new_n836), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT34), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n841), .A2(new_n842), .A3(new_n838), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n844), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n735), .A2(G25), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n629), .A2(G119), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n640), .A2(G131), .ZN(new_n852));
  OR2_X1    g427(.A1(G95), .A2(G2105), .ZN(new_n853));
  OAI211_X1 g428(.A(new_n853), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n851), .A2(new_n852), .A3(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n850), .B1(new_n856), .B2(new_n735), .ZN(new_n857));
  XNOR2_X1  g432(.A(KEYINPUT35), .B(G1991), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n857), .B(new_n859), .ZN(new_n860));
  NOR2_X1   g435(.A1(G16), .A2(G24), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n861), .B1(new_n601), .B2(G16), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n862), .B(G1986), .Z(new_n863));
  NAND2_X1  g438(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n790), .B1(new_n849), .B2(new_n865), .ZN(new_n866));
  AOI211_X1 g441(.A(KEYINPUT94), .B(new_n864), .C1(new_n844), .C2(new_n848), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n789), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  AND3_X1   g443(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n846), .B1(new_n845), .B2(new_n847), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n865), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(KEYINPUT94), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n849), .A2(new_n790), .A3(new_n865), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n872), .A2(KEYINPUT36), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n788), .B1(new_n868), .B2(new_n874), .ZN(new_n875));
  NOR2_X1   g450(.A1(G4), .A2(G16), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n876), .B1(new_n613), .B2(G16), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(G1348), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n786), .A2(G2072), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT98), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n735), .A2(G27), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n883), .B1(G164), .B2(new_n735), .ZN(new_n884));
  INV_X1    g459(.A(G2078), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n884), .B(new_n885), .ZN(new_n886));
  NAND4_X1  g461(.A1(new_n875), .A2(new_n879), .A3(new_n882), .A4(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(G311));
  NAND2_X1  g463(.A1(new_n887), .A2(KEYINPUT102), .ZN(new_n889));
  INV_X1    g464(.A(new_n886), .ZN(new_n890));
  AOI211_X1 g465(.A(new_n890), .B(new_n788), .C1(new_n868), .C2(new_n874), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT102), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n891), .A2(new_n892), .A3(new_n879), .A4(new_n882), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n889), .A2(new_n893), .ZN(G150));
  NAND2_X1  g469(.A1(new_n529), .A2(G55), .ZN(new_n895));
  AOI22_X1  g470(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n896));
  XNOR2_X1  g471(.A(KEYINPUT103), .B(G93), .ZN(new_n897));
  OAI221_X1 g472(.A(new_n895), .B1(new_n524), .B2(new_n896), .C1(new_n537), .C2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(G860), .ZN(new_n899));
  XOR2_X1   g474(.A(new_n899), .B(KEYINPUT37), .Z(new_n900));
  XNOR2_X1  g475(.A(new_n898), .B(new_n554), .ZN(new_n901));
  XOR2_X1   g476(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n902));
  XNOR2_X1  g477(.A(new_n901), .B(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n612), .A2(new_n623), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n903), .B(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n900), .B1(new_n905), .B2(G860), .ZN(G145));
  XOR2_X1   g481(.A(new_n760), .B(new_n730), .Z(new_n907));
  XNOR2_X1  g482(.A(new_n785), .B(G164), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n629), .A2(G130), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n640), .A2(G142), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n463), .A2(G118), .ZN(new_n912));
  XOR2_X1   g487(.A(new_n912), .B(KEYINPUT105), .Z(new_n913));
  OAI211_X1 g488(.A(new_n913), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n910), .A2(new_n911), .A3(new_n914), .ZN(new_n915));
  XOR2_X1   g490(.A(new_n915), .B(new_n646), .Z(new_n916));
  XNOR2_X1  g491(.A(new_n916), .B(new_n855), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n760), .B(new_n730), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n785), .B(new_n513), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n909), .A2(new_n917), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(KEYINPUT106), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n909), .A2(new_n920), .ZN(new_n923));
  INV_X1    g498(.A(new_n917), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n922), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n493), .B(KEYINPUT104), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n927), .B(new_n482), .ZN(new_n928));
  INV_X1    g503(.A(new_n642), .ZN(new_n929));
  OR2_X1    g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n928), .A2(new_n929), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n930), .A2(KEYINPUT107), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(KEYINPUT107), .B1(new_n930), .B2(new_n931), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n923), .A2(KEYINPUT106), .A3(new_n924), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n926), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(G37), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n925), .A2(new_n921), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n930), .A2(new_n931), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n936), .A2(new_n937), .A3(new_n940), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n941), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g517(.A1(new_n616), .A2(new_n613), .ZN(new_n943));
  NAND2_X1  g518(.A1(G299), .A2(new_n612), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT41), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n625), .B(new_n901), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n943), .A2(KEYINPUT41), .A3(new_n944), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  OR2_X1    g525(.A1(new_n948), .A2(new_n945), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(KEYINPUT108), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT108), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n812), .B(G303), .ZN(new_n956));
  XNOR2_X1  g531(.A(G290), .B(new_n794), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n956), .B1(new_n957), .B2(KEYINPUT109), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n958), .B1(KEYINPUT109), .B2(new_n957), .ZN(new_n959));
  INV_X1    g534(.A(new_n957), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT109), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n960), .A2(new_n961), .A3(new_n956), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n963), .B(KEYINPUT42), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n953), .A2(new_n955), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n965), .B1(new_n953), .B2(new_n955), .ZN(new_n967));
  OAI21_X1  g542(.A(G868), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n898), .A2(new_n617), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(G295));
  NAND2_X1  g545(.A1(new_n968), .A2(new_n969), .ZN(G331));
  INV_X1    g546(.A(KEYINPUT110), .ZN(new_n972));
  NAND2_X1  g547(.A1(G301), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(G171), .A2(KEYINPUT110), .ZN(new_n974));
  NAND3_X1  g549(.A1(G168), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(G286), .A2(new_n972), .A3(G301), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n901), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n901), .A2(new_n975), .A3(new_n976), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(KEYINPUT111), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n979), .A2(KEYINPUT111), .A3(new_n981), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n947), .A2(new_n983), .A3(new_n949), .A4(new_n984), .ZN(new_n985));
  AND2_X1   g560(.A1(new_n943), .A2(new_n944), .ZN(new_n986));
  OR3_X1    g561(.A1(new_n977), .A2(new_n978), .A3(KEYINPUT112), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n979), .A2(KEYINPUT112), .A3(new_n981), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n986), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n963), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n985), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n992), .A2(new_n937), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n963), .B(KEYINPUT113), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n947), .A2(new_n949), .A3(new_n987), .A4(new_n988), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n983), .A2(new_n984), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(new_n986), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n995), .A2(new_n999), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n993), .A2(KEYINPUT43), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n994), .B1(new_n985), .B2(new_n990), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(KEYINPUT43), .B1(new_n1003), .B2(new_n993), .ZN(new_n1004));
  OAI21_X1  g579(.A(KEYINPUT44), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT43), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n993), .A2(new_n1006), .A3(new_n1000), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n992), .A2(new_n937), .ZN(new_n1008));
  OAI21_X1  g583(.A(KEYINPUT43), .B1(new_n1008), .B2(new_n1002), .ZN(new_n1009));
  AND2_X1   g584(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1005), .B1(KEYINPUT44), .B2(new_n1010), .ZN(G397));
  INV_X1    g586(.A(G1384), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n513), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(KEYINPUT50), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n475), .A2(new_n479), .A3(G40), .A4(new_n480), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1015), .B1(new_n464), .B2(new_n473), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT50), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n513), .A2(new_n1017), .A3(new_n1012), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1014), .A2(new_n1016), .A3(new_n1018), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1019), .A2(G2090), .ZN(new_n1020));
  AND4_X1   g595(.A1(G40), .A2(new_n475), .A3(new_n479), .A4(new_n480), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n474), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT45), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1022), .B1(new_n1013), .B2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n513), .A2(KEYINPUT45), .A3(new_n1012), .ZN(new_n1025));
  AOI21_X1  g600(.A(G1971), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(G8), .B1(new_n1020), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(G303), .A2(G8), .ZN(new_n1028));
  XOR2_X1   g603(.A(new_n1028), .B(KEYINPUT55), .Z(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g606(.A1(G305), .A2(G1981), .ZN(new_n1032));
  INV_X1    g607(.A(G1981), .ZN(new_n1033));
  XOR2_X1   g608(.A(KEYINPUT116), .B(G86), .Z(new_n1034));
  NAND2_X1  g609(.A1(new_n538), .A2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1033), .B1(new_n591), .B2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1032), .A2(new_n1036), .ZN(new_n1037));
  OR2_X1    g612(.A1(new_n1037), .A2(KEYINPUT49), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1016), .A2(new_n513), .A3(new_n1012), .ZN(new_n1039));
  AND2_X1   g614(.A1(new_n1039), .A2(G8), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1037), .A2(KEYINPUT49), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1038), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n794), .A2(G1976), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1039), .A2(new_n1043), .A3(G8), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1045), .A2(KEYINPUT115), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1044), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(G1976), .ZN(new_n1049));
  NAND3_X1  g624(.A1(G288), .A2(new_n1045), .A3(new_n1049), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1039), .A2(new_n1043), .A3(G8), .A4(new_n1046), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1048), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  AND2_X1   g627(.A1(new_n1042), .A2(new_n1052), .ZN(new_n1053));
  OAI211_X1 g628(.A(G8), .B(new_n1029), .C1(new_n1020), .C2(new_n1026), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1031), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(G2084), .ZN(new_n1056));
  AND4_X1   g631(.A1(new_n1056), .A2(new_n1014), .A3(new_n1016), .A4(new_n1018), .ZN(new_n1057));
  AOI21_X1  g632(.A(G1966), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1058));
  OAI21_X1  g633(.A(G8), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(G286), .A2(G8), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1059), .A2(KEYINPUT51), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT51), .ZN(new_n1062));
  AND3_X1   g637(.A1(new_n513), .A2(KEYINPUT45), .A3(new_n1012), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT45), .B1(new_n513), .B2(new_n1012), .ZN(new_n1064));
  NOR3_X1   g639(.A1(new_n1063), .A2(new_n1064), .A3(new_n1022), .ZN(new_n1065));
  OAI22_X1  g640(.A1(new_n1065), .A2(G1966), .B1(new_n1019), .B2(G2084), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n1062), .B(G8), .C1(new_n1066), .C2(G286), .ZN(new_n1067));
  AND2_X1   g642(.A1(new_n1061), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1060), .ZN(new_n1069));
  AOI21_X1  g644(.A(KEYINPUT120), .B1(new_n1066), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1066), .A2(KEYINPUT120), .A3(new_n1069), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1055), .B1(new_n1068), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT54), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT53), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1013), .A2(new_n1023), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1077), .A2(new_n885), .A3(new_n1016), .A4(new_n1025), .ZN(new_n1078));
  INV_X1    g653(.A(G1961), .ZN(new_n1079));
  AOI22_X1  g654(.A1(new_n1076), .A2(new_n1078), .B1(new_n1019), .B2(new_n1079), .ZN(new_n1080));
  AND2_X1   g655(.A1(new_n1025), .A2(new_n885), .ZN(new_n1081));
  AND2_X1   g656(.A1(new_n472), .A2(KEYINPUT122), .ZN(new_n1082));
  OAI21_X1  g657(.A(G2105), .B1(new_n472), .B2(KEYINPUT122), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1021), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT123), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1021), .B(KEYINPUT123), .C1(new_n1083), .C2(new_n1082), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1081), .A2(KEYINPUT53), .A3(new_n1077), .A4(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(KEYINPUT124), .B1(new_n1080), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1078), .A2(new_n1076), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1019), .A2(new_n1079), .ZN(new_n1092));
  AND4_X1   g667(.A1(KEYINPUT124), .A2(new_n1091), .A3(new_n1092), .A4(new_n1089), .ZN(new_n1093));
  OAI21_X1  g668(.A(G171), .B1(new_n1090), .B2(new_n1093), .ZN(new_n1094));
  OR2_X1    g669(.A1(new_n1078), .A2(KEYINPUT121), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1078), .A2(KEYINPUT121), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1095), .A2(KEYINPUT53), .A3(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1097), .A2(G301), .A3(new_n1080), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1075), .B1(new_n1094), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(G301), .B1(new_n1097), .B2(new_n1080), .ZN(new_n1100));
  AND3_X1   g675(.A1(new_n1080), .A2(G301), .A3(new_n1089), .ZN(new_n1101));
  NOR3_X1   g676(.A1(new_n1100), .A2(KEYINPUT54), .A3(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1074), .B1(new_n1099), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT125), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT125), .ZN(new_n1105));
  OAI211_X1 g680(.A(new_n1074), .B(new_n1105), .C1(new_n1099), .C2(new_n1102), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT57), .ZN(new_n1107));
  XNOR2_X1  g682(.A(new_n572), .B(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g683(.A(KEYINPUT56), .B(G2072), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1065), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(G1956), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1019), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1108), .A2(new_n1110), .A3(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1108), .B1(new_n1112), .B2(new_n1110), .ZN(new_n1114));
  INV_X1    g689(.A(G1348), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1039), .ZN(new_n1116));
  AOI22_X1  g691(.A1(new_n1019), .A2(new_n1115), .B1(new_n738), .B2(new_n1116), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1117), .A2(new_n612), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1113), .B1(new_n1114), .B2(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g694(.A(new_n1119), .B(KEYINPUT119), .ZN(new_n1120));
  INV_X1    g695(.A(G1996), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1065), .A2(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g697(.A(KEYINPUT58), .B(G1341), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1122), .B1(new_n1116), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(new_n554), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(KEYINPUT59), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT59), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1124), .A2(new_n1127), .A3(new_n554), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1108), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(new_n1113), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT61), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1117), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1136), .A2(new_n613), .ZN(new_n1137));
  OAI21_X1  g712(.A(KEYINPUT60), .B1(new_n1137), .B2(new_n1118), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1132), .A2(KEYINPUT61), .A3(new_n1113), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1129), .A2(new_n1135), .A3(new_n1138), .A4(new_n1139), .ZN(new_n1140));
  NOR3_X1   g715(.A1(new_n1136), .A2(KEYINPUT60), .A3(new_n612), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1120), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1104), .A2(new_n1106), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1072), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1067), .B(new_n1061), .C1(new_n1144), .C2(new_n1070), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1055), .B1(new_n1145), .B2(KEYINPUT62), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT62), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1068), .A2(new_n1073), .A3(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1146), .A2(new_n1148), .A3(new_n1100), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1054), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(new_n1053), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n1032), .B(KEYINPUT117), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1042), .A2(new_n1049), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1152), .B1(new_n1153), .B2(G288), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(new_n1040), .ZN(new_n1155));
  AND3_X1   g730(.A1(new_n1149), .A2(new_n1151), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1059), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1031), .A2(new_n1053), .A3(new_n1054), .A4(new_n1157), .ZN(new_n1158));
  OR2_X1    g733(.A1(new_n1158), .A2(G286), .ZN(new_n1159));
  AOI21_X1  g734(.A(KEYINPUT63), .B1(new_n1159), .B2(KEYINPUT118), .ZN(new_n1160));
  OAI211_X1 g735(.A(KEYINPUT118), .B(KEYINPUT63), .C1(new_n1158), .C2(G286), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1143), .A2(new_n1156), .A3(new_n1163), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n760), .B(new_n1121), .ZN(new_n1165));
  XNOR2_X1  g740(.A(new_n730), .B(new_n738), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n855), .B(new_n858), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n1168), .B(KEYINPUT114), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n601), .B(G1986), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1077), .A2(new_n1022), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1164), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1166), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1173), .B1(new_n1176), .B2(new_n760), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT46), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1173), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1178), .B1(new_n1179), .B2(G1996), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1173), .A2(KEYINPUT46), .A3(new_n1121), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1177), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g757(.A(new_n1182), .B(KEYINPUT47), .ZN(new_n1183));
  NOR3_X1   g758(.A1(new_n1179), .A2(G1986), .A3(G290), .ZN(new_n1184));
  XNOR2_X1  g759(.A(new_n1184), .B(KEYINPUT127), .ZN(new_n1185));
  XNOR2_X1  g760(.A(new_n1185), .B(KEYINPUT48), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n1170), .A2(new_n1179), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1183), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  AOI211_X1 g763(.A(new_n858), .B(new_n855), .C1(new_n1167), .C2(new_n1173), .ZN(new_n1189));
  NOR2_X1   g764(.A1(new_n730), .A2(G2067), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  XNOR2_X1  g766(.A(new_n1191), .B(KEYINPUT126), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1188), .B1(new_n1192), .B2(new_n1173), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1175), .A2(new_n1193), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g769(.A(G227), .B1(new_n666), .B2(new_n667), .ZN(new_n1196));
  AND2_X1   g770(.A1(new_n941), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g771(.A(new_n458), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1198));
  AND3_X1   g772(.A1(new_n1197), .A2(new_n1198), .A3(new_n702), .ZN(G308));
  NAND3_X1  g773(.A1(new_n1197), .A2(new_n1198), .A3(new_n702), .ZN(G225));
endmodule


