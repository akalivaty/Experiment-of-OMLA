

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597;

  XNOR2_X1 U323 ( .A(n401), .B(n400), .ZN(n405) );
  XNOR2_X1 U324 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U325 ( .A(n472), .B(n471), .ZN(n560) );
  XNOR2_X1 U326 ( .A(n486), .B(n485), .ZN(n520) );
  XOR2_X1 U327 ( .A(n457), .B(n456), .Z(n545) );
  XOR2_X1 U328 ( .A(n415), .B(n414), .Z(n535) );
  XOR2_X1 U329 ( .A(n360), .B(n419), .Z(n291) );
  XNOR2_X1 U330 ( .A(KEYINPUT45), .B(KEYINPUT112), .ZN(n292) );
  XNOR2_X1 U331 ( .A(n417), .B(KEYINPUT54), .ZN(n293) );
  OR2_X1 U332 ( .A1(n560), .A2(n473), .ZN(n474) );
  XNOR2_X1 U333 ( .A(n368), .B(n367), .ZN(n369) );
  INV_X1 U334 ( .A(KEYINPUT95), .ZN(n398) );
  XNOR2_X1 U335 ( .A(n370), .B(n369), .ZN(n376) );
  XNOR2_X1 U336 ( .A(KEYINPUT19), .B(KEYINPUT86), .ZN(n410) );
  XNOR2_X1 U337 ( .A(n411), .B(KEYINPUT85), .ZN(n412) );
  INV_X1 U338 ( .A(KEYINPUT26), .ZN(n471) );
  XNOR2_X1 U339 ( .A(n413), .B(n412), .ZN(n455) );
  INV_X1 U340 ( .A(KEYINPUT121), .ZN(n494) );
  XNOR2_X1 U341 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n386) );
  XNOR2_X1 U342 ( .A(n497), .B(KEYINPUT126), .ZN(n498) );
  XNOR2_X1 U343 ( .A(n590), .B(n386), .ZN(n565) );
  INV_X1 U344 ( .A(G50GAT), .ZN(n487) );
  INV_X1 U345 ( .A(G43GAT), .ZN(n490) );
  XNOR2_X1 U346 ( .A(n499), .B(n498), .ZN(n501) );
  XNOR2_X1 U347 ( .A(n459), .B(G190GAT), .ZN(n460) );
  XNOR2_X1 U348 ( .A(n487), .B(KEYINPUT108), .ZN(n488) );
  XNOR2_X1 U349 ( .A(n490), .B(KEYINPUT40), .ZN(n491) );
  XNOR2_X1 U350 ( .A(n461), .B(n460), .ZN(G1351GAT) );
  XNOR2_X1 U351 ( .A(n489), .B(n488), .ZN(G1331GAT) );
  INV_X1 U352 ( .A(KEYINPUT8), .ZN(n294) );
  NAND2_X1 U353 ( .A1(G43GAT), .A2(n294), .ZN(n296) );
  NAND2_X1 U354 ( .A1(n490), .A2(KEYINPUT8), .ZN(n295) );
  NAND2_X1 U355 ( .A1(n296), .A2(n295), .ZN(n298) );
  XNOR2_X1 U356 ( .A(G29GAT), .B(KEYINPUT7), .ZN(n297) );
  XNOR2_X1 U357 ( .A(n298), .B(n297), .ZN(n360) );
  XOR2_X1 U358 ( .A(KEYINPUT76), .B(G134GAT), .Z(n419) );
  NAND2_X1 U359 ( .A1(G232GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U360 ( .A(n291), .B(n299), .ZN(n300) );
  XNOR2_X1 U361 ( .A(n300), .B(KEYINPUT75), .ZN(n303) );
  XNOR2_X1 U362 ( .A(G218GAT), .B(G36GAT), .ZN(n301) );
  XNOR2_X1 U363 ( .A(n301), .B(G190GAT), .ZN(n401) );
  XOR2_X1 U364 ( .A(n401), .B(KEYINPUT9), .Z(n302) );
  NAND2_X1 U365 ( .A1(n303), .A2(n302), .ZN(n305) );
  OR2_X1 U366 ( .A1(n303), .A2(n302), .ZN(n304) );
  NAND2_X1 U367 ( .A1(n305), .A2(n304), .ZN(n309) );
  XOR2_X1 U368 ( .A(G92GAT), .B(G106GAT), .Z(n307) );
  XNOR2_X1 U369 ( .A(KEYINPUT10), .B(KEYINPUT11), .ZN(n306) );
  XNOR2_X1 U370 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U371 ( .A(n309), .B(n308), .Z(n311) );
  XOR2_X1 U372 ( .A(G162GAT), .B(G50GAT), .Z(n318) );
  XOR2_X1 U373 ( .A(G85GAT), .B(G99GAT), .Z(n368) );
  XNOR2_X1 U374 ( .A(n318), .B(n368), .ZN(n310) );
  XNOR2_X2 U375 ( .A(n311), .B(n310), .ZN(n571) );
  XOR2_X1 U376 ( .A(KEYINPUT21), .B(G197GAT), .Z(n402) );
  XOR2_X1 U377 ( .A(n402), .B(G204GAT), .Z(n313) );
  XOR2_X1 U378 ( .A(G155GAT), .B(G22GAT), .Z(n332) );
  XNOR2_X1 U379 ( .A(G218GAT), .B(n332), .ZN(n312) );
  XNOR2_X1 U380 ( .A(n313), .B(n312), .ZN(n317) );
  XOR2_X1 U381 ( .A(KEYINPUT90), .B(KEYINPUT24), .Z(n315) );
  NAND2_X1 U382 ( .A1(G228GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U383 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U384 ( .A(n317), .B(n316), .Z(n320) );
  XNOR2_X1 U385 ( .A(n318), .B(G211GAT), .ZN(n319) );
  XNOR2_X1 U386 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U387 ( .A(KEYINPUT88), .B(KEYINPUT23), .Z(n322) );
  XNOR2_X1 U388 ( .A(KEYINPUT22), .B(KEYINPUT89), .ZN(n321) );
  XNOR2_X1 U389 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U390 ( .A(n324), .B(n323), .ZN(n329) );
  XNOR2_X1 U391 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n325) );
  XNOR2_X1 U392 ( .A(n325), .B(KEYINPUT2), .ZN(n418) );
  XOR2_X1 U393 ( .A(KEYINPUT71), .B(G78GAT), .Z(n327) );
  XNOR2_X1 U394 ( .A(G148GAT), .B(G106GAT), .ZN(n326) );
  XNOR2_X1 U395 ( .A(n327), .B(n326), .ZN(n381) );
  XNOR2_X1 U396 ( .A(n418), .B(n381), .ZN(n328) );
  XNOR2_X1 U397 ( .A(n329), .B(n328), .ZN(n468) );
  XNOR2_X1 U398 ( .A(KEYINPUT113), .B(KEYINPUT48), .ZN(n397) );
  XOR2_X1 U399 ( .A(KEYINPUT78), .B(KEYINPUT14), .Z(n331) );
  XNOR2_X1 U400 ( .A(G1GAT), .B(KEYINPUT15), .ZN(n330) );
  XNOR2_X1 U401 ( .A(n331), .B(n330), .ZN(n348) );
  XOR2_X1 U402 ( .A(G64GAT), .B(G78GAT), .Z(n334) );
  XOR2_X1 U403 ( .A(G127GAT), .B(G15GAT), .Z(n443) );
  XNOR2_X1 U404 ( .A(n443), .B(n332), .ZN(n333) );
  XNOR2_X1 U405 ( .A(n334), .B(n333), .ZN(n344) );
  XOR2_X1 U406 ( .A(G8GAT), .B(KEYINPUT77), .Z(n336) );
  XNOR2_X1 U407 ( .A(G183GAT), .B(G211GAT), .ZN(n335) );
  XNOR2_X1 U408 ( .A(n336), .B(n335), .ZN(n407) );
  XOR2_X1 U409 ( .A(KEYINPUT68), .B(KEYINPUT13), .Z(n338) );
  XNOR2_X1 U410 ( .A(G57GAT), .B(G71GAT), .ZN(n337) );
  XNOR2_X1 U411 ( .A(n338), .B(n337), .ZN(n370) );
  XNOR2_X1 U412 ( .A(n407), .B(n370), .ZN(n342) );
  XOR2_X1 U413 ( .A(KEYINPUT80), .B(KEYINPUT79), .Z(n340) );
  XNOR2_X1 U414 ( .A(KEYINPUT12), .B(KEYINPUT81), .ZN(n339) );
  XNOR2_X1 U415 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U416 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U417 ( .A(n344), .B(n343), .Z(n346) );
  NAND2_X1 U418 ( .A1(G231GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U419 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U420 ( .A(n348), .B(n347), .ZN(n596) );
  XOR2_X1 U421 ( .A(KEYINPUT111), .B(n596), .Z(n583) );
  XOR2_X1 U422 ( .A(G169GAT), .B(G15GAT), .Z(n350) );
  XNOR2_X1 U423 ( .A(G113GAT), .B(G141GAT), .ZN(n349) );
  XNOR2_X1 U424 ( .A(n350), .B(n349), .ZN(n364) );
  XOR2_X1 U425 ( .A(G36GAT), .B(G50GAT), .Z(n352) );
  NAND2_X1 U426 ( .A1(G229GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U427 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U428 ( .A(KEYINPUT66), .B(KEYINPUT67), .Z(n354) );
  XNOR2_X1 U429 ( .A(KEYINPUT29), .B(KEYINPUT30), .ZN(n353) );
  XNOR2_X1 U430 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U431 ( .A(n356), .B(n355), .Z(n362) );
  XOR2_X1 U432 ( .A(G197GAT), .B(G22GAT), .Z(n358) );
  XNOR2_X1 U433 ( .A(G1GAT), .B(G8GAT), .ZN(n357) );
  XNOR2_X1 U434 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U435 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U436 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U437 ( .A(n364), .B(n363), .ZN(n585) );
  INV_X1 U438 ( .A(n585), .ZN(n574) );
  XOR2_X1 U439 ( .A(KEYINPUT31), .B(KEYINPUT72), .Z(n366) );
  XNOR2_X1 U440 ( .A(G120GAT), .B(KEYINPUT70), .ZN(n365) );
  XNOR2_X1 U441 ( .A(n366), .B(n365), .ZN(n385) );
  AND2_X1 U442 ( .A1(G230GAT), .A2(G233GAT), .ZN(n367) );
  INV_X1 U443 ( .A(n376), .ZN(n374) );
  XOR2_X1 U444 ( .A(KEYINPUT73), .B(KEYINPUT69), .Z(n372) );
  XNOR2_X1 U445 ( .A(KEYINPUT33), .B(KEYINPUT32), .ZN(n371) );
  XOR2_X1 U446 ( .A(n372), .B(n371), .Z(n375) );
  INV_X1 U447 ( .A(n375), .ZN(n373) );
  NAND2_X1 U448 ( .A1(n374), .A2(n373), .ZN(n378) );
  NAND2_X1 U449 ( .A1(n376), .A2(n375), .ZN(n377) );
  NAND2_X1 U450 ( .A1(n378), .A2(n377), .ZN(n383) );
  XOR2_X1 U451 ( .A(G204GAT), .B(G176GAT), .Z(n380) );
  XNOR2_X1 U452 ( .A(G92GAT), .B(G64GAT), .ZN(n379) );
  XNOR2_X1 U453 ( .A(n380), .B(n379), .ZN(n406) );
  XNOR2_X1 U454 ( .A(n406), .B(n381), .ZN(n382) );
  XNOR2_X1 U455 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U456 ( .A(n385), .B(n384), .Z(n590) );
  NOR2_X1 U457 ( .A1(n574), .A2(n565), .ZN(n387) );
  XNOR2_X1 U458 ( .A(n387), .B(KEYINPUT46), .ZN(n388) );
  NOR2_X1 U459 ( .A1(n583), .A2(n388), .ZN(n389) );
  NAND2_X1 U460 ( .A1(n389), .A2(n571), .ZN(n390) );
  XNOR2_X1 U461 ( .A(n390), .B(KEYINPUT47), .ZN(n395) );
  XOR2_X1 U462 ( .A(KEYINPUT36), .B(n571), .Z(n496) );
  AND2_X1 U463 ( .A1(n496), .A2(n596), .ZN(n391) );
  XNOR2_X1 U464 ( .A(n391), .B(n292), .ZN(n393) );
  NOR2_X1 U465 ( .A1(n590), .A2(n585), .ZN(n392) );
  AND2_X1 U466 ( .A1(n393), .A2(n392), .ZN(n394) );
  NOR2_X1 U467 ( .A1(n395), .A2(n394), .ZN(n396) );
  XNOR2_X1 U468 ( .A(n397), .B(n396), .ZN(n543) );
  INV_X1 U469 ( .A(n543), .ZN(n416) );
  NAND2_X1 U470 ( .A1(G226GAT), .A2(G233GAT), .ZN(n399) );
  XNOR2_X1 U471 ( .A(n402), .B(KEYINPUT93), .ZN(n403) );
  XNOR2_X1 U472 ( .A(n403), .B(KEYINPUT94), .ZN(n404) );
  XOR2_X1 U473 ( .A(n405), .B(n404), .Z(n409) );
  XNOR2_X1 U474 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U475 ( .A(n409), .B(n408), .ZN(n415) );
  XNOR2_X1 U476 ( .A(n410), .B(G169GAT), .ZN(n413) );
  XNOR2_X1 U477 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n411) );
  INV_X1 U478 ( .A(n455), .ZN(n414) );
  NOR2_X1 U479 ( .A1(n416), .A2(n535), .ZN(n417) );
  XOR2_X1 U480 ( .A(n419), .B(n418), .Z(n421) );
  NAND2_X1 U481 ( .A1(G225GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U482 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U483 ( .A(n422), .B(KEYINPUT92), .Z(n426) );
  XOR2_X1 U484 ( .A(G113GAT), .B(G120GAT), .Z(n424) );
  XNOR2_X1 U485 ( .A(KEYINPUT0), .B(KEYINPUT82), .ZN(n423) );
  XNOR2_X1 U486 ( .A(n424), .B(n423), .ZN(n447) );
  XNOR2_X1 U487 ( .A(n447), .B(KEYINPUT4), .ZN(n425) );
  XNOR2_X1 U488 ( .A(n426), .B(n425), .ZN(n430) );
  XOR2_X1 U489 ( .A(G127GAT), .B(G85GAT), .Z(n428) );
  XNOR2_X1 U490 ( .A(G29GAT), .B(G162GAT), .ZN(n427) );
  XNOR2_X1 U491 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U492 ( .A(n430), .B(n429), .Z(n438) );
  XOR2_X1 U493 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n432) );
  XNOR2_X1 U494 ( .A(KEYINPUT5), .B(KEYINPUT91), .ZN(n431) );
  XNOR2_X1 U495 ( .A(n432), .B(n431), .ZN(n436) );
  XOR2_X1 U496 ( .A(G57GAT), .B(G1GAT), .Z(n434) );
  XNOR2_X1 U497 ( .A(G148GAT), .B(G155GAT), .ZN(n433) );
  XNOR2_X1 U498 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U499 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U500 ( .A(n438), .B(n437), .ZN(n533) );
  NAND2_X1 U501 ( .A1(n293), .A2(n533), .ZN(n493) );
  NOR2_X1 U502 ( .A1(n468), .A2(n493), .ZN(n440) );
  INV_X1 U503 ( .A(KEYINPUT55), .ZN(n439) );
  XNOR2_X1 U504 ( .A(n440), .B(n439), .ZN(n458) );
  XOR2_X1 U505 ( .A(G71GAT), .B(G183GAT), .Z(n442) );
  XNOR2_X1 U506 ( .A(G99GAT), .B(G43GAT), .ZN(n441) );
  XNOR2_X1 U507 ( .A(n442), .B(n441), .ZN(n444) );
  XOR2_X1 U508 ( .A(n444), .B(n443), .Z(n446) );
  XNOR2_X1 U509 ( .A(G134GAT), .B(G190GAT), .ZN(n445) );
  XNOR2_X1 U510 ( .A(n446), .B(n445), .ZN(n451) );
  XOR2_X1 U511 ( .A(n447), .B(KEYINPUT83), .Z(n449) );
  NAND2_X1 U512 ( .A1(G227GAT), .A2(G233GAT), .ZN(n448) );
  XNOR2_X1 U513 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U514 ( .A(n451), .B(n450), .Z(n457) );
  XOR2_X1 U515 ( .A(KEYINPUT84), .B(KEYINPUT87), .Z(n453) );
  XNOR2_X1 U516 ( .A(G176GAT), .B(KEYINPUT20), .ZN(n452) );
  XNOR2_X1 U517 ( .A(n453), .B(n452), .ZN(n454) );
  XOR2_X1 U518 ( .A(n455), .B(n454), .Z(n456) );
  INV_X1 U519 ( .A(n545), .ZN(n469) );
  NAND2_X1 U520 ( .A1(n458), .A2(n469), .ZN(n581) );
  NOR2_X1 U521 ( .A1(n571), .A2(n581), .ZN(n461) );
  INV_X1 U522 ( .A(KEYINPUT58), .ZN(n459) );
  XNOR2_X1 U523 ( .A(n535), .B(KEYINPUT27), .ZN(n473) );
  NOR2_X1 U524 ( .A1(n473), .A2(n533), .ZN(n462) );
  XNOR2_X1 U525 ( .A(n462), .B(KEYINPUT96), .ZN(n542) );
  XNOR2_X1 U526 ( .A(n468), .B(KEYINPUT65), .ZN(n463) );
  XNOR2_X1 U527 ( .A(KEYINPUT28), .B(n463), .ZN(n546) );
  NAND2_X1 U528 ( .A1(n542), .A2(n546), .ZN(n464) );
  NOR2_X1 U529 ( .A1(n469), .A2(n464), .ZN(n465) );
  XNOR2_X1 U530 ( .A(n465), .B(KEYINPUT97), .ZN(n479) );
  NOR2_X1 U531 ( .A1(n535), .A2(n545), .ZN(n466) );
  NOR2_X1 U532 ( .A1(n468), .A2(n466), .ZN(n467) );
  XNOR2_X1 U533 ( .A(n467), .B(KEYINPUT25), .ZN(n475) );
  INV_X1 U534 ( .A(n468), .ZN(n470) );
  NOR2_X1 U535 ( .A1(n470), .A2(n469), .ZN(n472) );
  NAND2_X1 U536 ( .A1(n475), .A2(n474), .ZN(n476) );
  NAND2_X1 U537 ( .A1(n533), .A2(n476), .ZN(n477) );
  XNOR2_X1 U538 ( .A(KEYINPUT98), .B(n477), .ZN(n478) );
  NAND2_X1 U539 ( .A1(n479), .A2(n478), .ZN(n480) );
  XNOR2_X1 U540 ( .A(n480), .B(KEYINPUT99), .ZN(n504) );
  NOR2_X1 U541 ( .A1(n504), .A2(n596), .ZN(n481) );
  XNOR2_X1 U542 ( .A(KEYINPUT104), .B(n481), .ZN(n482) );
  NAND2_X1 U543 ( .A1(n482), .A2(n496), .ZN(n483) );
  XNOR2_X1 U544 ( .A(n483), .B(KEYINPUT37), .ZN(n532) );
  NOR2_X1 U545 ( .A1(n590), .A2(n574), .ZN(n484) );
  XNOR2_X1 U546 ( .A(n484), .B(KEYINPUT74), .ZN(n505) );
  NAND2_X1 U547 ( .A1(n532), .A2(n505), .ZN(n486) );
  XOR2_X1 U548 ( .A(KEYINPUT38), .B(KEYINPUT105), .Z(n485) );
  NOR2_X1 U549 ( .A1(n520), .A2(n546), .ZN(n489) );
  NOR2_X1 U550 ( .A1(n520), .A2(n545), .ZN(n492) );
  XNOR2_X1 U551 ( .A(n492), .B(n491), .ZN(G1330GAT) );
  NOR2_X1 U552 ( .A1(n493), .A2(n560), .ZN(n495) );
  XNOR2_X1 U553 ( .A(n495), .B(n494), .ZN(n595) );
  NAND2_X1 U554 ( .A1(n595), .A2(n496), .ZN(n499) );
  XOR2_X1 U555 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n497) );
  XOR2_X1 U556 ( .A(G218GAT), .B(KEYINPUT125), .Z(n500) );
  XNOR2_X1 U557 ( .A(n501), .B(n500), .ZN(G1355GAT) );
  XNOR2_X1 U558 ( .A(KEYINPUT34), .B(KEYINPUT101), .ZN(n508) );
  NAND2_X1 U559 ( .A1(n571), .A2(n596), .ZN(n502) );
  XNOR2_X1 U560 ( .A(KEYINPUT16), .B(n502), .ZN(n503) );
  NOR2_X1 U561 ( .A1(n504), .A2(n503), .ZN(n523) );
  NAND2_X1 U562 ( .A1(n505), .A2(n523), .ZN(n506) );
  XNOR2_X1 U563 ( .A(n506), .B(KEYINPUT100), .ZN(n515) );
  NOR2_X1 U564 ( .A1(n533), .A2(n515), .ZN(n507) );
  XNOR2_X1 U565 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U566 ( .A(G1GAT), .B(n509), .ZN(G1324GAT) );
  NOR2_X1 U567 ( .A1(n535), .A2(n515), .ZN(n510) );
  XOR2_X1 U568 ( .A(G8GAT), .B(n510), .Z(G1325GAT) );
  NOR2_X1 U569 ( .A1(n545), .A2(n515), .ZN(n514) );
  XOR2_X1 U570 ( .A(KEYINPUT102), .B(KEYINPUT35), .Z(n512) );
  XNOR2_X1 U571 ( .A(G15GAT), .B(KEYINPUT103), .ZN(n511) );
  XNOR2_X1 U572 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U573 ( .A(n514), .B(n513), .ZN(G1326GAT) );
  NOR2_X1 U574 ( .A1(n515), .A2(n546), .ZN(n516) );
  XOR2_X1 U575 ( .A(G22GAT), .B(n516), .Z(G1327GAT) );
  NOR2_X1 U576 ( .A1(n520), .A2(n533), .ZN(n519) );
  XNOR2_X1 U577 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n517) );
  XNOR2_X1 U578 ( .A(n517), .B(KEYINPUT106), .ZN(n518) );
  XNOR2_X1 U579 ( .A(n519), .B(n518), .ZN(G1328GAT) );
  XNOR2_X1 U580 ( .A(G36GAT), .B(KEYINPUT107), .ZN(n522) );
  NOR2_X1 U581 ( .A1(n535), .A2(n520), .ZN(n521) );
  XNOR2_X1 U582 ( .A(n522), .B(n521), .ZN(G1329GAT) );
  XOR2_X1 U583 ( .A(n565), .B(KEYINPUT109), .Z(n576) );
  NOR2_X1 U584 ( .A1(n576), .A2(n585), .ZN(n531) );
  NAND2_X1 U585 ( .A1(n531), .A2(n523), .ZN(n528) );
  NOR2_X1 U586 ( .A1(n533), .A2(n528), .ZN(n524) );
  XOR2_X1 U587 ( .A(G57GAT), .B(n524), .Z(n525) );
  XNOR2_X1 U588 ( .A(KEYINPUT42), .B(n525), .ZN(G1332GAT) );
  NOR2_X1 U589 ( .A1(n535), .A2(n528), .ZN(n526) );
  XOR2_X1 U590 ( .A(G64GAT), .B(n526), .Z(G1333GAT) );
  NOR2_X1 U591 ( .A1(n545), .A2(n528), .ZN(n527) );
  XOR2_X1 U592 ( .A(G71GAT), .B(n527), .Z(G1334GAT) );
  NOR2_X1 U593 ( .A1(n546), .A2(n528), .ZN(n530) );
  XNOR2_X1 U594 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n529) );
  XNOR2_X1 U595 ( .A(n530), .B(n529), .ZN(G1335GAT) );
  NAND2_X1 U596 ( .A1(n532), .A2(n531), .ZN(n538) );
  NOR2_X1 U597 ( .A1(n533), .A2(n538), .ZN(n534) );
  XOR2_X1 U598 ( .A(G85GAT), .B(n534), .Z(G1336GAT) );
  NOR2_X1 U599 ( .A1(n535), .A2(n538), .ZN(n536) );
  XOR2_X1 U600 ( .A(G92GAT), .B(n536), .Z(G1337GAT) );
  NOR2_X1 U601 ( .A1(n545), .A2(n538), .ZN(n537) );
  XOR2_X1 U602 ( .A(G99GAT), .B(n537), .Z(G1338GAT) );
  NOR2_X1 U603 ( .A1(n546), .A2(n538), .ZN(n540) );
  XNOR2_X1 U604 ( .A(KEYINPUT44), .B(KEYINPUT110), .ZN(n539) );
  XNOR2_X1 U605 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U606 ( .A(G106GAT), .B(n541), .Z(G1339GAT) );
  NAND2_X1 U607 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U608 ( .A(KEYINPUT114), .B(n544), .ZN(n559) );
  NOR2_X1 U609 ( .A1(n559), .A2(n545), .ZN(n547) );
  NAND2_X1 U610 ( .A1(n547), .A2(n546), .ZN(n556) );
  NOR2_X1 U611 ( .A1(n574), .A2(n556), .ZN(n549) );
  XNOR2_X1 U612 ( .A(G113GAT), .B(KEYINPUT115), .ZN(n548) );
  XNOR2_X1 U613 ( .A(n549), .B(n548), .ZN(G1340GAT) );
  NOR2_X1 U614 ( .A1(n576), .A2(n556), .ZN(n551) );
  XNOR2_X1 U615 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n551), .B(n550), .ZN(G1341GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n554) );
  INV_X1 U618 ( .A(n556), .ZN(n552) );
  NAND2_X1 U619 ( .A1(n552), .A2(n583), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n554), .B(n553), .ZN(n555) );
  XOR2_X1 U621 ( .A(G127GAT), .B(n555), .Z(G1342GAT) );
  NOR2_X1 U622 ( .A1(n571), .A2(n556), .ZN(n558) );
  XNOR2_X1 U623 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(G1343GAT) );
  XOR2_X1 U625 ( .A(G141GAT), .B(KEYINPUT117), .Z(n562) );
  NOR2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n568) );
  NAND2_X1 U627 ( .A1(n568), .A2(n585), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(G1344GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n564) );
  XNOR2_X1 U630 ( .A(G148GAT), .B(KEYINPUT118), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(n567) );
  INV_X1 U632 ( .A(n568), .ZN(n570) );
  NOR2_X1 U633 ( .A1(n565), .A2(n570), .ZN(n566) );
  XOR2_X1 U634 ( .A(n567), .B(n566), .Z(G1345GAT) );
  NAND2_X1 U635 ( .A1(n596), .A2(n568), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n569), .B(G155GAT), .ZN(G1346GAT) );
  NOR2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n573) );
  XNOR2_X1 U638 ( .A(G162GAT), .B(KEYINPUT119), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(G1347GAT) );
  NOR2_X1 U640 ( .A1(n574), .A2(n581), .ZN(n575) );
  XOR2_X1 U641 ( .A(G169GAT), .B(n575), .Z(G1348GAT) );
  XNOR2_X1 U642 ( .A(KEYINPUT120), .B(KEYINPUT57), .ZN(n580) );
  NOR2_X1 U643 ( .A1(n576), .A2(n581), .ZN(n578) );
  XNOR2_X1 U644 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n577) );
  XNOR2_X1 U645 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n580), .B(n579), .ZN(G1349GAT) );
  INV_X1 U647 ( .A(n581), .ZN(n582) );
  NAND2_X1 U648 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n584), .B(G183GAT), .ZN(G1350GAT) );
  AND2_X1 U650 ( .A1(n585), .A2(n595), .ZN(n589) );
  XNOR2_X1 U651 ( .A(G197GAT), .B(KEYINPUT122), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n586), .B(KEYINPUT60), .ZN(n587) );
  XNOR2_X1 U653 ( .A(KEYINPUT59), .B(n587), .ZN(n588) );
  XNOR2_X1 U654 ( .A(n589), .B(n588), .ZN(G1352GAT) );
  AND2_X1 U655 ( .A1(n595), .A2(n590), .ZN(n594) );
  XOR2_X1 U656 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n592) );
  XNOR2_X1 U657 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n591) );
  XNOR2_X1 U658 ( .A(n592), .B(n591), .ZN(n593) );
  XNOR2_X1 U659 ( .A(n594), .B(n593), .ZN(G1353GAT) );
  AND2_X1 U660 ( .A1(n596), .A2(n595), .ZN(n597) );
  XOR2_X1 U661 ( .A(G211GAT), .B(n597), .Z(G1354GAT) );
endmodule

