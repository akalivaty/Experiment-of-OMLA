//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 1 1 1 1 0 1 0 0 0 0 1 1 1 1 1 0 1 0 1 0 0 0 1 0 0 0 0 1 0 1 1 0 0 1 0 0 1 0 1 0 1 1 0 0 0 1 0 0 0 0 1 1 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:42 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n545, new_n546, new_n547, new_n548, new_n549, new_n552,
    new_n553, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n607, new_n610, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n846, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n946, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT64), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT65), .Z(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  XOR2_X1   g031(.A(G325), .B(KEYINPUT66), .Z(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  XNOR2_X1  g036(.A(KEYINPUT67), .B(G2105), .ZN(new_n462));
  OR2_X1    g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n462), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n465), .A2(new_n462), .A3(G137), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n468), .A2(new_n473), .ZN(G160));
  AND2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NOR2_X1   g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n477), .A2(new_n462), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n477), .A2(G2105), .ZN(new_n479));
  AOI22_X1  g054(.A1(G124), .A2(new_n478), .B1(new_n479), .B2(G136), .ZN(new_n480));
  OAI221_X1 g055(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n462), .C2(G112), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT68), .ZN(G162));
  AND2_X1   g058(.A1(G126), .A2(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n484), .B1(new_n475), .B2(new_n476), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n470), .A2(G114), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g063(.A(G138), .B1(new_n475), .B2(new_n476), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n470), .A2(KEYINPUT67), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT67), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(KEYINPUT4), .B1(new_n489), .B2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n465), .A2(new_n462), .A3(new_n495), .A4(G138), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n488), .B1(new_n494), .B2(new_n496), .ZN(G164));
  OR2_X1    g072(.A1(KEYINPUT5), .A2(G543), .ZN(new_n498));
  NAND2_X1  g073(.A1(KEYINPUT5), .A2(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n500), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n501));
  INV_X1    g076(.A(G651), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OR2_X1    g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n500), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G88), .ZN(new_n508));
  INV_X1    g083(.A(G50), .ZN(new_n509));
  AND2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  OAI21_X1  g086(.A(G543), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  OAI22_X1  g087(.A1(new_n507), .A2(new_n508), .B1(new_n509), .B2(new_n512), .ZN(new_n513));
  OR2_X1    g088(.A1(new_n503), .A2(new_n513), .ZN(G303));
  INV_X1    g089(.A(G303), .ZN(G166));
  XNOR2_X1  g090(.A(KEYINPUT70), .B(G89), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n506), .A2(new_n516), .B1(G63), .B2(G651), .ZN(new_n517));
  AND2_X1   g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  NOR2_X1   g093(.A1(KEYINPUT5), .A2(G543), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  OR2_X1    g095(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT69), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n512), .A2(new_n522), .ZN(new_n523));
  OAI211_X1 g098(.A(KEYINPUT69), .B(G543), .C1(new_n510), .C2(new_n511), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G51), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  AND3_X1   g103(.A1(new_n521), .A2(new_n526), .A3(new_n528), .ZN(G168));
  INV_X1    g104(.A(KEYINPUT71), .ZN(new_n530));
  INV_X1    g105(.A(G64), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n531), .B1(new_n498), .B2(new_n499), .ZN(new_n532));
  NAND2_X1  g107(.A1(G77), .A2(G543), .ZN(new_n533));
  INV_X1    g108(.A(new_n533), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n530), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  OAI211_X1 g110(.A(KEYINPUT71), .B(new_n533), .C1(new_n520), .C2(new_n531), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n535), .A2(G651), .A3(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT72), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g114(.A1(new_n535), .A2(new_n536), .A3(KEYINPUT72), .A4(G651), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n498), .A2(new_n499), .B1(new_n504), .B2(new_n505), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n525), .A2(G52), .B1(G90), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n539), .A2(new_n540), .A3(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  NAND2_X1  g119(.A1(new_n525), .A2(G43), .ZN(new_n545));
  NAND2_X1  g120(.A1(G68), .A2(G543), .ZN(new_n546));
  INV_X1    g121(.A(G56), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n520), .B2(new_n547), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n548), .A2(G651), .B1(new_n541), .B2(G81), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n545), .A2(new_n549), .A3(G860), .ZN(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(G188));
  INV_X1    g129(.A(G65), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n555), .B1(new_n498), .B2(new_n499), .ZN(new_n556));
  AND2_X1   g131(.A1(G78), .A2(G543), .ZN(new_n557));
  OAI21_X1  g132(.A(G651), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n541), .A2(G91), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT9), .ZN(new_n560));
  INV_X1    g135(.A(G543), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n561), .B1(new_n504), .B2(new_n505), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n560), .B1(new_n562), .B2(G53), .ZN(new_n563));
  OAI211_X1 g138(.A(G53), .B(G543), .C1(new_n510), .C2(new_n511), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n564), .A2(KEYINPUT9), .ZN(new_n565));
  OAI211_X1 g140(.A(new_n558), .B(new_n559), .C1(new_n563), .C2(new_n565), .ZN(G299));
  NAND3_X1  g141(.A1(new_n521), .A2(new_n526), .A3(new_n528), .ZN(G286));
  OAI21_X1  g142(.A(G651), .B1(new_n500), .B2(G74), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n562), .A2(G49), .ZN(new_n569));
  INV_X1    g144(.A(G87), .ZN(new_n570));
  OAI211_X1 g145(.A(new_n568), .B(new_n569), .C1(new_n570), .C2(new_n507), .ZN(G288));
  NAND2_X1  g146(.A1(G73), .A2(G543), .ZN(new_n572));
  INV_X1    g147(.A(G61), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n520), .B2(new_n573), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n574), .A2(G651), .B1(G48), .B2(new_n562), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n541), .A2(G86), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(G305));
  INV_X1    g152(.A(G60), .ZN(new_n578));
  INV_X1    g153(.A(G72), .ZN(new_n579));
  OAI22_X1  g154(.A1(new_n520), .A2(new_n578), .B1(new_n579), .B2(new_n561), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n502), .B1(new_n580), .B2(KEYINPUT73), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n581), .B1(KEYINPUT73), .B2(new_n580), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n525), .A2(G47), .B1(G85), .B2(new_n541), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(G290));
  NAND2_X1  g159(.A1(G301), .A2(G868), .ZN(new_n585));
  AOI21_X1  g160(.A(KEYINPUT10), .B1(new_n541), .B2(G92), .ZN(new_n586));
  AND4_X1   g161(.A1(KEYINPUT10), .A2(new_n500), .A3(new_n506), .A4(G92), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g163(.A(KEYINPUT69), .B1(new_n506), .B2(G543), .ZN(new_n589));
  INV_X1    g164(.A(new_n524), .ZN(new_n590));
  OAI21_X1  g165(.A(G54), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  OAI21_X1  g166(.A(G66), .B1(new_n518), .B2(new_n519), .ZN(new_n592));
  NAND2_X1  g167(.A1(G79), .A2(G543), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n502), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n591), .A2(KEYINPUT74), .A3(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT74), .ZN(new_n597));
  INV_X1    g172(.A(G54), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n598), .B1(new_n523), .B2(new_n524), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n597), .B1(new_n599), .B2(new_n594), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n588), .B1(new_n596), .B2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT75), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n601), .B(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n585), .B1(new_n603), .B2(G868), .ZN(G284));
  OAI21_X1  g179(.A(new_n585), .B1(new_n603), .B2(G868), .ZN(G321));
  INV_X1    g180(.A(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(G299), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n607), .B1(G168), .B2(new_n606), .ZN(G297));
  OAI21_X1  g183(.A(new_n607), .B1(G168), .B2(new_n606), .ZN(G280));
  INV_X1    g184(.A(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n603), .B1(new_n610), .B2(G860), .ZN(G148));
  NAND2_X1  g186(.A1(new_n545), .A2(new_n549), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n603), .A2(new_n610), .ZN(new_n613));
  MUX2_X1   g188(.A(new_n612), .B(new_n613), .S(G868), .Z(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g190(.A1(new_n465), .A2(new_n471), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT12), .ZN(new_n617));
  XNOR2_X1  g192(.A(KEYINPUT76), .B(KEYINPUT13), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n619), .A2(G2100), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(G2100), .ZN(new_n621));
  INV_X1    g196(.A(G111), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT77), .ZN(new_n623));
  OAI21_X1  g198(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n624));
  AOI22_X1  g199(.A1(new_n493), .A2(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(new_n623), .B2(new_n624), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n479), .A2(G135), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n478), .A2(G123), .ZN(new_n628));
  AND3_X1   g203(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2096), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n620), .A2(new_n621), .A3(new_n630), .ZN(G156));
  INV_X1    g206(.A(G14), .ZN(new_n632));
  XOR2_X1   g207(.A(KEYINPUT15), .B(G2435), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2438), .ZN(new_n634));
  XOR2_X1   g209(.A(G2427), .B(G2430), .Z(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT79), .B(KEYINPUT14), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n634), .A2(new_n635), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n639), .B(new_n640), .Z(new_n641));
  XOR2_X1   g216(.A(G2451), .B(G2454), .Z(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n641), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G1341), .B(G1348), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT80), .Z(new_n647));
  AOI21_X1  g222(.A(new_n632), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(KEYINPUT81), .ZN(new_n649));
  AND2_X1   g224(.A1(new_n641), .A2(new_n644), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n641), .A2(new_n644), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(new_n647), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n649), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NOR3_X1   g229(.A1(new_n645), .A2(KEYINPUT81), .A3(new_n647), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n648), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(KEYINPUT82), .ZN(new_n657));
  INV_X1    g232(.A(KEYINPUT82), .ZN(new_n658));
  OAI211_X1 g233(.A(new_n648), .B(new_n658), .C1(new_n654), .C2(new_n655), .ZN(new_n659));
  AND2_X1   g234(.A1(new_n657), .A2(new_n659), .ZN(G401));
  INV_X1    g235(.A(KEYINPUT18), .ZN(new_n661));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  XNOR2_X1  g237(.A(G2067), .B(G2678), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n664), .A2(KEYINPUT17), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n662), .A2(new_n663), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n661), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(G2100), .ZN(new_n668));
  XOR2_X1   g243(.A(G2072), .B(G2078), .Z(new_n669));
  AOI21_X1  g244(.A(new_n669), .B1(new_n664), .B2(KEYINPUT18), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G2096), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n668), .B(new_n671), .ZN(G227));
  XNOR2_X1  g247(.A(G1991), .B(G1996), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(G1986), .ZN(new_n675));
  XOR2_X1   g250(.A(G1971), .B(G1976), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT19), .ZN(new_n677));
  XOR2_X1   g252(.A(G1956), .B(G2474), .Z(new_n678));
  XOR2_X1   g253(.A(G1961), .B(G1966), .Z(new_n679));
  AND2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT20), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n678), .A2(new_n679), .ZN(new_n684));
  OR3_X1    g259(.A1(new_n677), .A2(new_n680), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n677), .A2(new_n684), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(G1981), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n688), .A2(new_n689), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n675), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n692), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n694), .A2(new_n690), .A3(G1986), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT83), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n693), .A2(new_n695), .A3(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n698), .B1(new_n693), .B2(new_n695), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n674), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n693), .A2(new_n695), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(new_n697), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n704), .A2(new_n699), .A3(new_n673), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n702), .A2(new_n705), .ZN(G229));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G22), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(G166), .B2(new_n707), .ZN(new_n709));
  INV_X1    g284(.A(G1971), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n707), .A2(G6), .ZN(new_n712));
  INV_X1    g287(.A(G305), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n712), .B1(new_n713), .B2(new_n707), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT32), .B(G1981), .Z(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  NOR2_X1   g291(.A1(G16), .A2(G23), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT88), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT89), .ZN(new_n719));
  NAND2_X1  g294(.A1(G288), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n541), .A2(G87), .ZN(new_n721));
  NAND4_X1  g296(.A1(new_n721), .A2(KEYINPUT89), .A3(new_n568), .A4(new_n569), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n718), .B1(new_n723), .B2(new_n707), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT33), .B(G1976), .Z(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n711), .A2(new_n716), .A3(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT34), .ZN(new_n728));
  INV_X1    g303(.A(G29), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(G25), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n478), .A2(G119), .ZN(new_n731));
  OAI221_X1 g306(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n462), .C2(G107), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n479), .A2(G131), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT84), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n730), .B1(new_n737), .B2(new_n729), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT35), .B(G1991), .Z(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT85), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n738), .B(new_n740), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n741), .A2(KEYINPUT86), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n741), .A2(KEYINPUT86), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n707), .A2(G24), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT87), .Z(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(G290), .B2(G16), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(new_n675), .ZN(new_n747));
  NOR4_X1   g322(.A1(new_n728), .A2(new_n742), .A3(new_n743), .A4(new_n747), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT36), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n729), .A2(G35), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G162), .B2(new_n729), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT29), .Z(new_n752));
  INV_X1    g327(.A(G2090), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n752), .A2(new_n753), .ZN(new_n755));
  NOR2_X1   g330(.A1(G171), .A2(new_n707), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G5), .B2(new_n707), .ZN(new_n757));
  INV_X1    g332(.A(G1961), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n755), .A2(new_n759), .ZN(new_n760));
  AOI211_X1 g335(.A(new_n754), .B(new_n760), .C1(new_n758), .C2(new_n757), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n729), .A2(G26), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT28), .Z(new_n763));
  AOI22_X1  g338(.A1(G128), .A2(new_n478), .B1(new_n479), .B2(G140), .ZN(new_n764));
  OAI221_X1 g339(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n462), .C2(G116), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n763), .B1(new_n766), .B2(G29), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G2067), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT30), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT96), .ZN(new_n770));
  AND3_X1   g345(.A1(new_n770), .A2(new_n769), .A3(G28), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n770), .B1(new_n769), .B2(G28), .ZN(new_n772));
  OAI221_X1 g347(.A(new_n729), .B1(new_n769), .B2(G28), .C1(new_n771), .C2(new_n772), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT31), .B(G11), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n629), .A2(G29), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n775), .B1(new_n776), .B2(KEYINPUT95), .ZN(new_n777));
  OAI211_X1 g352(.A(new_n768), .B(new_n777), .C1(KEYINPUT95), .C2(new_n776), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n729), .A2(G32), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n479), .A2(G141), .B1(G105), .B2(new_n471), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n478), .A2(G129), .ZN(new_n781));
  NAND3_X1  g356(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT26), .Z(new_n783));
  NAND3_X1  g358(.A1(new_n780), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n779), .B1(new_n785), .B2(new_n729), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT27), .B(G1996), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n786), .B(new_n787), .Z(new_n788));
  NAND2_X1  g363(.A1(new_n729), .A2(G27), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT98), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G164), .B2(new_n729), .ZN(new_n791));
  INV_X1    g366(.A(G2078), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT99), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT24), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n729), .B1(new_n796), .B2(G34), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(new_n796), .B2(G34), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G160), .B2(G29), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n799), .A2(G2084), .ZN(new_n800));
  NOR4_X1   g375(.A1(new_n778), .A2(new_n788), .A3(new_n795), .A4(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n799), .A2(G2084), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT97), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n707), .A2(G21), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G168), .B2(new_n707), .ZN(new_n805));
  INV_X1    g380(.A(G1966), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n707), .A2(G20), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT23), .ZN(new_n809));
  INV_X1    g384(.A(G299), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n809), .B1(new_n810), .B2(new_n707), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(G1956), .Z(new_n812));
  NAND4_X1  g387(.A1(new_n801), .A2(new_n803), .A3(new_n807), .A4(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(G2072), .ZN(new_n814));
  AOI22_X1  g389(.A1(new_n465), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n815), .A2(new_n462), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT25), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n817), .A2(new_n818), .ZN(new_n820));
  AOI22_X1  g395(.A1(new_n819), .A2(new_n820), .B1(G139), .B2(new_n479), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT92), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n821), .A2(new_n822), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n816), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n825), .A2(KEYINPUT93), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT93), .ZN(new_n827));
  AOI211_X1 g402(.A(new_n827), .B(new_n816), .C1(new_n823), .C2(new_n824), .ZN(new_n828));
  OAI21_X1  g403(.A(G29), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n729), .A2(G33), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n814), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  MUX2_X1   g406(.A(G19), .B(new_n612), .S(G16), .Z(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT91), .ZN(new_n833));
  XOR2_X1   g408(.A(KEYINPUT90), .B(G1341), .Z(new_n834));
  AOI22_X1  g409(.A1(new_n833), .A2(new_n834), .B1(new_n794), .B2(new_n793), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(new_n834), .B2(new_n833), .ZN(new_n836));
  NOR3_X1   g411(.A1(new_n813), .A2(new_n831), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n707), .A2(G4), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n838), .B1(new_n603), .B2(new_n707), .ZN(new_n839));
  INV_X1    g414(.A(G1348), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n829), .A2(new_n814), .A3(new_n830), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT94), .Z(new_n843));
  NAND4_X1  g418(.A1(new_n761), .A2(new_n837), .A3(new_n841), .A4(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n749), .A2(new_n844), .ZN(G311));
  INV_X1    g420(.A(KEYINPUT36), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n748), .B(new_n846), .ZN(new_n847));
  AND2_X1   g422(.A1(new_n843), .A2(new_n841), .ZN(new_n848));
  NAND4_X1  g423(.A1(new_n847), .A2(new_n761), .A3(new_n837), .A4(new_n848), .ZN(G150));
  NAND2_X1  g424(.A1(G80), .A2(G543), .ZN(new_n850));
  INV_X1    g425(.A(G67), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n850), .B1(new_n520), .B2(new_n851), .ZN(new_n852));
  AOI22_X1  g427(.A1(new_n852), .A2(G651), .B1(new_n541), .B2(G93), .ZN(new_n853));
  OAI21_X1  g428(.A(G55), .B1(new_n589), .B2(new_n590), .ZN(new_n854));
  AND3_X1   g429(.A1(new_n853), .A2(new_n854), .A3(KEYINPUT100), .ZN(new_n855));
  AOI21_X1  g430(.A(KEYINPUT100), .B1(new_n853), .B2(new_n854), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n612), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n545), .A2(new_n549), .A3(new_n853), .A4(new_n854), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT38), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n603), .A2(G559), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n860), .B(new_n861), .Z(new_n862));
  AND2_X1   g437(.A1(new_n862), .A2(KEYINPUT39), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n862), .A2(KEYINPUT39), .ZN(new_n864));
  NOR3_X1   g439(.A1(new_n863), .A2(new_n864), .A3(G860), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n855), .A2(new_n856), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(G860), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT37), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n865), .A2(new_n868), .ZN(G145));
  XNOR2_X1  g444(.A(G162), .B(G160), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n870), .B(new_n629), .Z(new_n871));
  OR2_X1    g446(.A1(new_n825), .A2(KEYINPUT93), .ZN(new_n872));
  INV_X1    g447(.A(new_n828), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n785), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NOR3_X1   g449(.A1(new_n826), .A2(new_n828), .A3(new_n784), .ZN(new_n875));
  AOI22_X1  g450(.A1(G130), .A2(new_n478), .B1(new_n479), .B2(G142), .ZN(new_n876));
  OAI221_X1 g451(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n462), .C2(G118), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(new_n617), .ZN(new_n879));
  NOR3_X1   g454(.A1(new_n874), .A2(new_n875), .A3(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n879), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n872), .A2(new_n873), .A3(new_n785), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n784), .B1(new_n826), .B2(new_n828), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n494), .A2(new_n496), .ZN(new_n885));
  INV_X1    g460(.A(new_n488), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n766), .B(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(new_n734), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  NOR3_X1   g465(.A1(new_n880), .A2(new_n884), .A3(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n879), .B1(new_n874), .B2(new_n875), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n882), .A2(new_n883), .A3(new_n881), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n889), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n871), .B1(new_n891), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n890), .B1(new_n880), .B2(new_n884), .ZN(new_n896));
  INV_X1    g471(.A(new_n871), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n892), .A2(new_n889), .A3(new_n893), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n895), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(KEYINPUT101), .B(G37), .ZN(new_n901));
  AOI21_X1  g476(.A(KEYINPUT40), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT40), .ZN(new_n903));
  INV_X1    g478(.A(new_n901), .ZN(new_n904));
  AOI211_X1 g479(.A(new_n903), .B(new_n904), .C1(new_n895), .C2(new_n899), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n902), .A2(new_n905), .ZN(G395));
  NAND3_X1  g481(.A1(new_n603), .A2(new_n610), .A3(new_n859), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n588), .ZN(new_n909));
  AOI21_X1  g484(.A(KEYINPUT74), .B1(new_n591), .B2(new_n595), .ZN(new_n910));
  NOR3_X1   g485(.A1(new_n599), .A2(new_n597), .A3(new_n594), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(G299), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n601), .A2(new_n810), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n913), .A2(KEYINPUT102), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(KEYINPUT102), .B1(new_n913), .B2(new_n914), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n859), .B1(new_n603), .B2(new_n610), .ZN(new_n918));
  OR3_X1    g493(.A1(new_n908), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n596), .A2(new_n600), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n810), .B1(new_n920), .B2(new_n909), .ZN(new_n921));
  AOI211_X1 g496(.A(G299), .B(new_n588), .C1(new_n596), .C2(new_n600), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT41), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n923), .A2(KEYINPUT103), .A3(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(KEYINPUT41), .B1(new_n921), .B2(new_n922), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n913), .A2(new_n924), .A3(new_n914), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT103), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  OAI211_X1 g504(.A(new_n925), .B(new_n929), .C1(new_n908), .C2(new_n918), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n723), .A2(new_n713), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n720), .A2(G305), .A3(new_n722), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(G166), .A2(G290), .ZN(new_n934));
  NAND3_X1  g509(.A1(G303), .A2(new_n582), .A3(new_n583), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n934), .A2(new_n935), .A3(new_n931), .A4(new_n932), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n939), .B(KEYINPUT42), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n919), .A2(new_n930), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n940), .B1(new_n919), .B2(new_n930), .ZN(new_n942));
  OAI21_X1  g517(.A(G868), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n866), .A2(new_n606), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(G331));
  INV_X1    g520(.A(KEYINPUT104), .ZN(new_n946));
  XNOR2_X1  g521(.A(G331), .B(new_n946), .ZN(G295));
  NAND2_X1  g522(.A1(G301), .A2(G168), .ZN(new_n948));
  NAND4_X1  g523(.A1(G286), .A2(new_n539), .A3(new_n540), .A4(new_n542), .ZN(new_n949));
  AND4_X1   g524(.A1(new_n857), .A2(new_n948), .A3(new_n858), .A4(new_n949), .ZN(new_n950));
  AOI22_X1  g525(.A1(new_n948), .A2(new_n949), .B1(new_n857), .B2(new_n858), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n952), .A2(new_n929), .A3(new_n925), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n923), .B1(new_n950), .B2(new_n951), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n953), .A2(new_n939), .A3(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT43), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n939), .B1(new_n953), .B2(new_n954), .ZN(new_n958));
  NOR3_X1   g533(.A1(new_n957), .A2(G37), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n948), .A2(new_n949), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n960), .B(new_n859), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n939), .B1(new_n961), .B2(new_n917), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n952), .A2(new_n927), .A3(new_n926), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n904), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n956), .B1(new_n964), .B2(new_n955), .ZN(new_n965));
  OAI21_X1  g540(.A(KEYINPUT44), .B1(new_n959), .B2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT44), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n964), .A2(new_n956), .A3(new_n955), .ZN(new_n968));
  AND3_X1   g543(.A1(new_n953), .A2(new_n939), .A3(new_n954), .ZN(new_n969));
  NOR3_X1   g544(.A1(new_n969), .A2(new_n958), .A3(G37), .ZN(new_n970));
  OAI211_X1 g545(.A(new_n967), .B(new_n968), .C1(new_n970), .C2(new_n956), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT105), .ZN(new_n972));
  AND3_X1   g547(.A1(new_n966), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n972), .B1(new_n966), .B2(new_n971), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n973), .A2(new_n974), .ZN(G397));
  XOR2_X1   g550(.A(KEYINPUT106), .B(G1384), .Z(new_n976));
  AOI21_X1  g551(.A(new_n976), .B1(new_n885), .B2(new_n886), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n977), .A2(KEYINPUT45), .ZN(new_n978));
  INV_X1    g553(.A(G125), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n467), .B1(new_n477), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n493), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n981), .A2(G40), .A3(new_n472), .A4(new_n469), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n978), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G2067), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n766), .B(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(G1996), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n784), .B(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n984), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  XOR2_X1   g564(.A(new_n989), .B(KEYINPUT107), .Z(new_n990));
  XNOR2_X1  g565(.A(new_n734), .B(new_n740), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n990), .B1(new_n984), .B2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(new_n984), .ZN(new_n993));
  XNOR2_X1  g568(.A(G290), .B(G1986), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n992), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT45), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n996), .B1(G164), .B2(G1384), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(KEYINPUT108), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n982), .B1(new_n977), .B2(KEYINPUT45), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT108), .ZN(new_n1000));
  OAI211_X1 g575(.A(new_n1000), .B(new_n996), .C1(G164), .C2(G1384), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n998), .A2(new_n999), .A3(new_n792), .A4(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT53), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NOR3_X1   g579(.A1(G164), .A2(new_n996), .A3(G1384), .ZN(new_n1005));
  OR2_X1    g580(.A1(new_n1005), .A2(KEYINPUT114), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n997), .A2(new_n983), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1003), .A2(G2078), .ZN(new_n1008));
  INV_X1    g583(.A(G1384), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n887), .A2(KEYINPUT114), .A3(KEYINPUT45), .A4(new_n1009), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .A4(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT50), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n887), .A2(new_n1012), .A3(new_n1009), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1013), .A2(new_n1014), .A3(new_n983), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(new_n758), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1004), .A2(new_n1011), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(G171), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT122), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT122), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1017), .A2(new_n1020), .A3(G171), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n999), .B(new_n1008), .C1(KEYINPUT45), .C2(new_n977), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1004), .A2(new_n1016), .A3(new_n1022), .ZN(new_n1023));
  OR2_X1    g598(.A1(new_n1023), .A2(G171), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1019), .A2(new_n1021), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT123), .ZN(new_n1026));
  XOR2_X1   g601(.A(KEYINPUT121), .B(KEYINPUT54), .Z(new_n1027));
  AND3_X1   g602(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1026), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n998), .A2(new_n999), .A3(new_n1001), .ZN(new_n1031));
  AND3_X1   g606(.A1(new_n1013), .A2(new_n1014), .A3(new_n983), .ZN(new_n1032));
  AOI22_X1  g607(.A1(new_n1031), .A2(new_n710), .B1(new_n1032), .B2(new_n753), .ZN(new_n1033));
  INV_X1    g608(.A(G8), .ZN(new_n1034));
  NAND2_X1  g609(.A1(G303), .A2(G8), .ZN(new_n1035));
  XNOR2_X1  g610(.A(KEYINPUT109), .B(KEYINPUT55), .ZN(new_n1036));
  XNOR2_X1  g611(.A(new_n1035), .B(new_n1036), .ZN(new_n1037));
  OR3_X1    g612(.A1(new_n1033), .A2(new_n1034), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT111), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1039), .B1(G305), .B2(G1981), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n575), .A2(KEYINPUT111), .A3(new_n689), .A4(new_n576), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  XNOR2_X1  g617(.A(KEYINPUT112), .B(G86), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n575), .B1(new_n507), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(G1981), .ZN(new_n1045));
  AOI21_X1  g620(.A(KEYINPUT49), .B1(new_n1042), .B2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(G164), .A2(G1384), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n983), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(G8), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1046), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1042), .A2(KEYINPUT49), .A3(new_n1045), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n720), .A2(G1976), .A3(new_n722), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1048), .A2(new_n1052), .A3(G8), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT110), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT52), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(KEYINPUT52), .A2(G1976), .ZN(new_n1058));
  AOI22_X1  g633(.A1(new_n1053), .A2(new_n1057), .B1(G288), .B2(new_n1058), .ZN(new_n1059));
  OR2_X1    g634(.A1(new_n1053), .A2(new_n1057), .ZN(new_n1060));
  AOI22_X1  g635(.A1(new_n1050), .A2(new_n1051), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1037), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1038), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  OR2_X1    g638(.A1(new_n1017), .A2(G171), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT54), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1065), .B1(new_n1023), .B2(G171), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1063), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1010), .A2(new_n983), .A3(new_n997), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1005), .A2(KEYINPUT114), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n806), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(G2084), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1032), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT119), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(G286), .A2(G8), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1070), .A2(new_n1072), .A3(KEYINPUT119), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1075), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(KEYINPUT51), .A2(G8), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1075), .A2(new_n1078), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1080), .B1(new_n1081), .B2(G168), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1073), .A2(G8), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1077), .A2(KEYINPUT51), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1083), .A2(KEYINPUT120), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT120), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1034), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1084), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1086), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1085), .A2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1079), .B1(new_n1082), .B2(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g666(.A(KEYINPUT56), .B(G2072), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n998), .A2(new_n999), .A3(new_n1001), .A4(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g668(.A(KEYINPUT115), .B(G1956), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1015), .A2(new_n1094), .ZN(new_n1095));
  XOR2_X1   g670(.A(G299), .B(KEYINPUT57), .Z(new_n1096));
  NAND3_X1  g671(.A1(new_n1093), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  NOR2_X1   g672(.A1(KEYINPUT118), .A2(KEYINPUT61), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1096), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1093), .A2(new_n1095), .A3(KEYINPUT61), .A4(new_n1096), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1099), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT60), .ZN(new_n1105));
  NOR4_X1   g680(.A1(new_n982), .A2(G164), .A3(G1384), .A4(G2067), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1106), .B1(new_n1015), .B2(new_n840), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1105), .B1(new_n1107), .B2(new_n601), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1108), .B1(new_n601), .B2(new_n1107), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1107), .A2(new_n1105), .A3(new_n601), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1104), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n998), .A2(new_n999), .A3(new_n987), .A4(new_n1001), .ZN(new_n1112));
  XOR2_X1   g687(.A(KEYINPUT58), .B(G1341), .Z(new_n1113));
  AOI22_X1  g688(.A1(new_n1112), .A2(KEYINPUT117), .B1(new_n1048), .B2(new_n1113), .ZN(new_n1114));
  AND2_X1   g689(.A1(new_n998), .A2(new_n999), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT117), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1115), .A2(new_n1116), .A3(new_n987), .A4(new_n1001), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n612), .B1(new_n1114), .B2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1118), .A2(KEYINPUT59), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT59), .ZN(new_n1120));
  AOI211_X1 g695(.A(new_n1120), .B(new_n612), .C1(new_n1114), .C2(new_n1117), .ZN(new_n1121));
  NOR3_X1   g696(.A1(new_n1111), .A2(new_n1119), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1097), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1107), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(new_n601), .ZN(new_n1125));
  OR2_X1    g700(.A1(new_n1125), .A2(KEYINPUT116), .ZN(new_n1126));
  AOI22_X1  g701(.A1(new_n1125), .A2(KEYINPUT116), .B1(new_n1101), .B2(new_n1100), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1123), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1067), .B(new_n1091), .C1(new_n1122), .C2(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1030), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1131));
  NOR2_X1   g706(.A1(G288), .A2(G1976), .ZN(new_n1132));
  AOI22_X1  g707(.A1(new_n1131), .A2(new_n1132), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1133));
  XOR2_X1   g708(.A(new_n1049), .B(KEYINPUT113), .Z(new_n1134));
  INV_X1    g709(.A(new_n1061), .ZN(new_n1135));
  OAI22_X1  g710(.A1(new_n1133), .A2(new_n1134), .B1(new_n1135), .B2(new_n1038), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1083), .A2(G286), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1137), .A2(KEYINPUT63), .A3(new_n1038), .A4(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT63), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1138), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1140), .B1(new_n1063), .B2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1136), .B1(new_n1139), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT62), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1079), .B(new_n1144), .C1(new_n1082), .C2(new_n1090), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1063), .B1(new_n1021), .B2(new_n1019), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(G286), .B1(new_n1075), .B2(new_n1078), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n1089), .B(new_n1085), .C1(new_n1148), .C2(new_n1080), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1144), .B1(new_n1149), .B2(new_n1079), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1143), .B1(new_n1147), .B2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n995), .B1(new_n1130), .B2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n984), .B1(new_n986), .B2(new_n785), .ZN(new_n1153));
  OR3_X1    g728(.A1(new_n984), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1154));
  OAI21_X1  g729(.A(KEYINPUT46), .B1(new_n984), .B2(G1996), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1153), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g731(.A(KEYINPUT126), .B(KEYINPUT47), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n1156), .B(new_n1157), .ZN(new_n1158));
  NOR3_X1   g733(.A1(new_n984), .A2(G1986), .A3(G290), .ZN(new_n1159));
  XOR2_X1   g734(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n1160));
  XNOR2_X1  g735(.A(new_n1159), .B(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1158), .B1(new_n992), .B2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n766), .A2(G2067), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n737), .A2(new_n740), .ZN(new_n1164));
  XOR2_X1   g739(.A(new_n1164), .B(KEYINPUT124), .Z(new_n1165));
  AOI21_X1  g740(.A(new_n1163), .B1(new_n990), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT125), .ZN(new_n1167));
  OR2_X1    g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n984), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1162), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1152), .A2(new_n1170), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g746(.A1(new_n900), .A2(new_n901), .ZN(new_n1173));
  NOR2_X1   g747(.A1(G227), .A2(new_n460), .ZN(new_n1174));
  NAND3_X1  g748(.A1(new_n702), .A2(new_n705), .A3(new_n1174), .ZN(new_n1175));
  AOI21_X1  g749(.A(new_n1175), .B1(new_n657), .B2(new_n659), .ZN(new_n1176));
  OAI21_X1  g750(.A(new_n968), .B1(new_n970), .B2(new_n956), .ZN(new_n1177));
  AND3_X1   g751(.A1(new_n1173), .A2(new_n1176), .A3(new_n1177), .ZN(G308));
  NAND3_X1  g752(.A1(new_n1173), .A2(new_n1176), .A3(new_n1177), .ZN(G225));
endmodule


