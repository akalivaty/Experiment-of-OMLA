//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 0 0 1 0 0 0 0 0 1 0 0 1 0 1 1 0 0 0 0 0 1 1 1 1 0 0 0 1 1 1 1 1 0 1 1 1 1 0 0 1 1 1 1 0 0 1 0 1 0 1 1 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:38 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1298, new_n1299, new_n1300, new_n1301, new_n1302, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1377,
    new_n1378, new_n1379, new_n1380, new_n1381;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n206), .A2(new_n207), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  INV_X1    g0016(.A(G20), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n220), .B1(new_n202), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n211), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n214), .B(new_n219), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XOR2_X1   g0030(.A(G250), .B(G257), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT65), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  INV_X1    g0035(.A(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(KEYINPUT2), .B(G226), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n234), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT66), .ZN(new_n242));
  XOR2_X1   g0042(.A(G107), .B(G116), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  NAND2_X1  g0048(.A1(new_n208), .A2(G20), .ZN(new_n249));
  NOR2_X1   g0049(.A1(G20), .A2(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G150), .ZN(new_n251));
  XNOR2_X1  g0051(.A(KEYINPUT8), .B(G58), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n217), .A2(G33), .ZN(new_n253));
  OAI211_X1 g0053(.A(new_n249), .B(new_n251), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(new_n216), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G1), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n258), .A2(G13), .A3(G20), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT67), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND4_X1  g0061(.A1(new_n258), .A2(KEYINPUT67), .A3(G13), .A4(G20), .ZN(new_n262));
  AND2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(new_n207), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n263), .A2(new_n256), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n258), .A2(G20), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n265), .A2(G50), .A3(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n257), .A2(new_n264), .A3(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT9), .ZN(new_n270));
  INV_X1    g0070(.A(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(KEYINPUT3), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT3), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G1698), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AOI22_X1  g0077(.A1(new_n277), .A2(G223), .B1(G77), .B2(new_n275), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT3), .B(G33), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n279), .A2(G222), .A3(new_n276), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G41), .ZN(new_n284));
  INV_X1    g0084(.A(G45), .ZN(new_n285));
  AOI21_X1  g0085(.A(G1), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(G33), .A2(G41), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n287), .A2(G1), .A3(G13), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n286), .A2(new_n288), .A3(G274), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n282), .A2(new_n286), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n290), .B1(G226), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n283), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G200), .ZN(new_n294));
  INV_X1    g0094(.A(new_n293), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G190), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT9), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n268), .A2(new_n297), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n270), .A2(new_n294), .A3(new_n296), .A4(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT10), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n300), .B1(new_n294), .B2(KEYINPUT70), .ZN(new_n301));
  OR2_X1    g0101(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n299), .A2(new_n301), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G169), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n269), .B1(new_n305), .B2(new_n293), .ZN(new_n306));
  OR2_X1    g0106(.A1(new_n306), .A2(KEYINPUT68), .ZN(new_n307));
  INV_X1    g0107(.A(G179), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n306), .A2(KEYINPUT68), .B1(new_n308), .B2(new_n295), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  AND2_X1   g0110(.A1(new_n304), .A2(new_n310), .ZN(new_n311));
  OR2_X1    g0111(.A1(G226), .A2(G1698), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n236), .A2(G1698), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n279), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT71), .ZN(new_n315));
  NAND2_X1  g0115(.A1(G33), .A2(G97), .ZN(new_n316));
  AND3_X1   g0116(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n315), .B1(new_n314), .B2(new_n316), .ZN(new_n318));
  NOR3_X1   g0118(.A1(new_n317), .A2(new_n318), .A3(new_n288), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n258), .B1(G41), .B2(G45), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n288), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n289), .B1(new_n221), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(KEYINPUT72), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT72), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n289), .B(new_n324), .C1(new_n221), .C2(new_n321), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(KEYINPUT13), .B1(new_n319), .B2(new_n326), .ZN(new_n327));
  AND2_X1   g0127(.A1(new_n323), .A2(new_n325), .ZN(new_n328));
  INV_X1    g0128(.A(new_n318), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n329), .A2(new_n282), .A3(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT13), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n328), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n327), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G169), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(KEYINPUT14), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n327), .A2(new_n333), .A3(G179), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT14), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n334), .A2(new_n338), .A3(G169), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n336), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n261), .A2(new_n202), .A3(new_n262), .ZN(new_n341));
  XNOR2_X1  g0141(.A(new_n341), .B(KEYINPUT12), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n261), .A2(new_n262), .ZN(new_n344));
  INV_X1    g0144(.A(new_n256), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n344), .A2(new_n345), .A3(G68), .A4(new_n266), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n250), .A2(G50), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n202), .A2(G20), .ZN(new_n348));
  INV_X1    g0148(.A(G77), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n347), .B(new_n348), .C1(new_n349), .C2(new_n253), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT11), .ZN(new_n351));
  AND3_X1   g0151(.A1(new_n350), .A2(new_n351), .A3(new_n256), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n351), .B1(new_n350), .B2(new_n256), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n346), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(KEYINPUT73), .B1(new_n343), .B2(new_n354), .ZN(new_n355));
  OR2_X1    g0155(.A1(new_n352), .A2(new_n353), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT73), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n356), .A2(new_n357), .A3(new_n342), .A4(new_n346), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n340), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT74), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n327), .A2(new_n333), .A3(G190), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n359), .ZN(new_n364));
  INV_X1    g0164(.A(G200), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n365), .B1(new_n327), .B2(new_n333), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n362), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n366), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n368), .A2(KEYINPUT74), .A3(new_n359), .A4(new_n363), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n252), .ZN(new_n371));
  AOI22_X1  g0171(.A1(new_n371), .A2(new_n250), .B1(G20), .B2(G77), .ZN(new_n372));
  XNOR2_X1  g0172(.A(KEYINPUT15), .B(G87), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n372), .B1(new_n253), .B2(new_n373), .ZN(new_n374));
  AOI22_X1  g0174(.A1(new_n374), .A2(new_n256), .B1(new_n349), .B2(new_n263), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n265), .A2(G77), .A3(new_n266), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n290), .B1(G244), .B2(new_n291), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n279), .A2(G232), .A3(new_n276), .ZN(new_n380));
  XNOR2_X1  g0180(.A(KEYINPUT69), .B(G107), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n380), .B1(new_n279), .B2(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n382), .B1(G238), .B2(new_n277), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n379), .B1(new_n383), .B2(new_n288), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(G200), .ZN(new_n385));
  INV_X1    g0185(.A(G190), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n378), .B(new_n385), .C1(new_n386), .C2(new_n384), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n384), .A2(new_n305), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n388), .B(new_n377), .C1(G179), .C2(new_n384), .ZN(new_n389));
  AND2_X1   g0189(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n311), .A2(new_n361), .A3(new_n370), .A4(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n252), .B1(new_n258), .B2(G20), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n265), .A2(new_n392), .B1(new_n263), .B2(new_n252), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT75), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n272), .A2(new_n274), .A3(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT76), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT7), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n397), .A2(G20), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n271), .A2(KEYINPUT75), .A3(KEYINPUT3), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n395), .A2(new_n396), .A3(new_n398), .A4(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n397), .B1(new_n279), .B2(G20), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n399), .A2(new_n398), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n396), .B1(new_n404), .B2(new_n395), .ZN(new_n405));
  OAI21_X1  g0205(.A(G68), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n203), .B(new_n205), .C1(new_n201), .C2(new_n202), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n407), .A2(G20), .B1(G159), .B2(new_n250), .ZN(new_n408));
  AOI21_X1  g0208(.A(KEYINPUT16), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n275), .A2(new_n217), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n410), .A2(new_n397), .B1(new_n275), .B2(new_n398), .ZN(new_n411));
  OAI211_X1 g0211(.A(KEYINPUT16), .B(new_n408), .C1(new_n411), .C2(new_n202), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n256), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n393), .B1(new_n409), .B2(new_n413), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n272), .A2(new_n274), .A3(G223), .A4(new_n276), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n272), .A2(new_n274), .A3(G226), .A4(G1698), .ZN(new_n416));
  NAND2_X1  g0216(.A1(G33), .A2(G87), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n282), .ZN(new_n419));
  INV_X1    g0219(.A(G274), .ZN(new_n420));
  INV_X1    g0220(.A(new_n216), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n420), .B1(new_n421), .B2(new_n287), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n291), .A2(G232), .B1(new_n422), .B2(new_n286), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n419), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(G169), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(new_n308), .B2(new_n424), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n414), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(KEYINPUT18), .ZN(new_n428));
  OR2_X1    g0228(.A1(new_n409), .A2(new_n413), .ZN(new_n429));
  AND3_X1   g0229(.A1(new_n419), .A2(new_n423), .A3(G190), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n365), .B1(new_n419), .B2(new_n423), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n429), .A2(KEYINPUT17), .A3(new_n393), .A4(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT18), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n414), .A2(new_n426), .A3(new_n434), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n432), .B(new_n393), .C1(new_n409), .C2(new_n413), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT17), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n428), .A2(new_n433), .A3(new_n435), .A4(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n391), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT77), .ZN(new_n441));
  INV_X1    g0241(.A(new_n381), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n441), .B(new_n442), .C1(new_n402), .C2(new_n405), .ZN(new_n443));
  INV_X1    g0243(.A(G107), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n444), .A2(KEYINPUT6), .A3(G97), .ZN(new_n445));
  INV_X1    g0245(.A(G97), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n446), .A2(new_n444), .ZN(new_n447));
  NOR2_X1   g0247(.A1(G97), .A2(G107), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n445), .B1(new_n449), .B2(KEYINPUT6), .ZN(new_n450));
  AOI22_X1  g0250(.A1(new_n450), .A2(G20), .B1(G77), .B2(new_n250), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n443), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n395), .ZN(new_n453));
  OAI21_X1  g0253(.A(KEYINPUT76), .B1(new_n453), .B2(new_n403), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n454), .A2(new_n401), .A3(new_n400), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n441), .B1(new_n455), .B2(new_n442), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n256), .B1(new_n452), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n344), .A2(new_n446), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n271), .A2(G1), .ZN(new_n459));
  AOI211_X1 g0259(.A(new_n459), .B(new_n256), .C1(new_n261), .C2(new_n262), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n458), .B1(new_n460), .B2(new_n446), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n272), .A2(new_n274), .A3(G244), .A4(new_n276), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT4), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G250), .A2(G1698), .ZN(new_n465));
  NAND2_X1  g0265(.A1(KEYINPUT4), .A2(G244), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n465), .B1(new_n466), .B2(G1698), .ZN(new_n467));
  AOI22_X1  g0267(.A1(new_n279), .A2(new_n467), .B1(G33), .B2(G283), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n288), .B1(new_n464), .B2(new_n468), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n258), .B(G45), .C1(new_n284), .C2(KEYINPUT5), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT5), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n471), .A2(G41), .ZN(new_n472));
  OAI211_X1 g0272(.A(G257), .B(new_n288), .C1(new_n470), .C2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n288), .A2(G274), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT78), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n475), .B1(new_n471), .B2(G41), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n284), .A2(KEYINPUT78), .A3(KEYINPUT5), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n285), .A2(G1), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n471), .A2(G41), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n476), .A2(new_n477), .A3(new_n478), .A4(new_n479), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n473), .B1(new_n474), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n469), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n386), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n483), .B1(G200), .B2(new_n482), .ZN(new_n484));
  AND3_X1   g0284(.A1(new_n457), .A2(new_n461), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n464), .A2(new_n468), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n282), .ZN(new_n487));
  INV_X1    g0287(.A(new_n481), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n487), .A2(new_n488), .A3(G179), .ZN(new_n489));
  OAI21_X1  g0289(.A(G169), .B1(new_n469), .B2(new_n481), .ZN(new_n490));
  AND2_X1   g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n491), .B1(new_n457), .B2(new_n461), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n272), .A2(new_n274), .A3(new_n217), .A4(G68), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n253), .A2(new_n446), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n493), .B1(KEYINPUT19), .B2(new_n494), .ZN(new_n495));
  NOR2_X1   g0295(.A1(G87), .A2(G97), .ZN(new_n496));
  NAND3_X1  g0296(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n381), .A2(new_n496), .B1(new_n217), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n256), .B1(new_n495), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n263), .A2(new_n373), .ZN(new_n500));
  INV_X1    g0300(.A(new_n459), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n344), .A2(new_n345), .A3(G87), .A4(new_n501), .ZN(new_n502));
  AND3_X1   g0302(.A1(new_n499), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n272), .A2(new_n274), .A3(G244), .A4(G1698), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n272), .A2(new_n274), .A3(G238), .A4(new_n276), .ZN(new_n505));
  NAND2_X1  g0305(.A1(G33), .A2(G116), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n282), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n223), .B1(new_n285), .B2(G1), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n258), .A2(new_n420), .A3(G45), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n288), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(G200), .ZN(new_n513));
  INV_X1    g0313(.A(new_n511), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n514), .B1(new_n507), .B2(new_n282), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(G190), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n503), .A2(new_n513), .A3(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n373), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n344), .A2(new_n345), .A3(new_n518), .A4(new_n501), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n499), .A2(new_n500), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n515), .A2(new_n308), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n520), .B(new_n521), .C1(G169), .C2(new_n515), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n517), .A2(new_n522), .ZN(new_n523));
  NOR3_X1   g0323(.A1(new_n485), .A2(new_n492), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n460), .A2(G107), .ZN(new_n525));
  OAI211_X1 g0325(.A(KEYINPUT81), .B(KEYINPUT25), .C1(new_n344), .C2(G107), .ZN(new_n526));
  XOR2_X1   g0326(.A(KEYINPUT81), .B(KEYINPUT25), .Z(new_n527));
  NAND3_X1  g0327(.A1(new_n263), .A2(new_n444), .A3(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n525), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT24), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n272), .A2(new_n274), .A3(new_n217), .A4(G87), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(KEYINPUT22), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT22), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n279), .A2(new_n533), .A3(new_n217), .A4(G87), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT23), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n536), .A2(new_n444), .A3(G20), .ZN(new_n537));
  INV_X1    g0337(.A(G116), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n537), .B1(new_n538), .B2(new_n253), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n381), .A2(G20), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n539), .B1(new_n540), .B2(KEYINPUT23), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n530), .B1(new_n535), .B2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n535), .A2(new_n541), .A3(new_n530), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n529), .B1(new_n545), .B2(new_n256), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n272), .A2(new_n274), .A3(G257), .A4(G1698), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n272), .A2(new_n274), .A3(G250), .A4(new_n276), .ZN(new_n548));
  NAND2_X1  g0348(.A1(G33), .A2(G294), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n282), .ZN(new_n551));
  OR2_X1    g0351(.A1(new_n480), .A2(new_n474), .ZN(new_n552));
  OAI211_X1 g0352(.A(G264), .B(new_n288), .C1(new_n470), .C2(new_n472), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT82), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n554), .A2(new_n555), .A3(G169), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n555), .B1(new_n554), .B2(G169), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT83), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n551), .A2(new_n560), .A3(new_n553), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n560), .B1(new_n551), .B2(new_n553), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n563), .A2(G179), .A3(new_n552), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n546), .B1(new_n559), .B2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n544), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n256), .B1(new_n566), .B2(new_n542), .ZN(new_n567));
  INV_X1    g0367(.A(new_n529), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n551), .A2(new_n553), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(KEYINPUT83), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n551), .A2(new_n560), .A3(new_n553), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n571), .A2(new_n552), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n365), .ZN(new_n574));
  INV_X1    g0374(.A(new_n554), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n386), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n569), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n565), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n263), .A2(new_n538), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n344), .A2(new_n345), .A3(G116), .A4(new_n501), .ZN(new_n580));
  AND2_X1   g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n255), .A2(new_n216), .B1(G20), .B2(new_n538), .ZN(new_n582));
  AOI21_X1  g0382(.A(G20), .B1(G33), .B2(G283), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(G33), .B2(new_n446), .ZN(new_n584));
  AND3_X1   g0384(.A1(new_n582), .A2(new_n584), .A3(KEYINPUT20), .ZN(new_n585));
  AOI21_X1  g0385(.A(KEYINPUT20), .B1(new_n582), .B2(new_n584), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n581), .A2(new_n588), .A3(KEYINPUT79), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT79), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n579), .A2(new_n580), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n590), .B1(new_n591), .B2(new_n587), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n288), .B1(new_n470), .B2(new_n472), .ZN(new_n594));
  INV_X1    g0394(.A(G270), .ZN(new_n595));
  OAI22_X1  g0395(.A1(new_n594), .A2(new_n595), .B1(new_n480), .B2(new_n474), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n272), .A2(new_n274), .A3(G264), .A4(G1698), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n272), .A2(new_n274), .A3(G257), .A4(new_n276), .ZN(new_n598));
  INV_X1    g0398(.A(G303), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n597), .B(new_n598), .C1(new_n599), .C2(new_n279), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n596), .B1(new_n282), .B2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n602), .A2(new_n386), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n601), .A2(new_n365), .ZN(new_n604));
  NOR3_X1   g0404(.A1(new_n593), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n600), .A2(new_n282), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  OAI211_X1 g0407(.A(KEYINPUT21), .B(G169), .C1(new_n607), .C2(new_n596), .ZN(new_n608));
  OR2_X1    g0408(.A1(new_n594), .A2(new_n595), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n606), .A2(G179), .A3(new_n552), .A4(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  AND2_X1   g0411(.A1(new_n611), .A2(new_n593), .ZN(new_n612));
  XNOR2_X1  g0412(.A(KEYINPUT80), .B(KEYINPUT21), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n601), .A2(new_n305), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n614), .B1(new_n593), .B2(new_n615), .ZN(new_n616));
  NOR3_X1   g0416(.A1(new_n605), .A2(new_n612), .A3(new_n616), .ZN(new_n617));
  AND4_X1   g0417(.A1(new_n440), .A2(new_n524), .A3(new_n578), .A4(new_n617), .ZN(G372));
  INV_X1    g0418(.A(new_n558), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n619), .B(new_n556), .C1(new_n573), .C2(new_n308), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n569), .ZN(new_n621));
  AOI21_X1  g0421(.A(KEYINPUT79), .B1(new_n581), .B2(new_n588), .ZN(new_n622));
  NOR3_X1   g0422(.A1(new_n591), .A2(new_n587), .A3(new_n590), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n615), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n624), .A2(new_n613), .B1(new_n611), .B2(new_n593), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n485), .A2(new_n492), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n577), .A2(new_n523), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n517), .A2(new_n522), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n492), .A2(KEYINPUT26), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n457), .A2(new_n461), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT85), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n489), .A2(new_n633), .A3(new_n490), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n633), .B1(new_n489), .B2(new_n490), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n630), .A2(new_n632), .A3(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n631), .B1(new_n637), .B2(KEYINPUT26), .ZN(new_n638));
  XNOR2_X1  g0438(.A(new_n522), .B(KEYINPUT84), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n629), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n440), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g0441(.A(new_n436), .B(KEYINPUT17), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n368), .A2(new_n359), .A3(new_n363), .ZN(new_n644));
  INV_X1    g0444(.A(new_n389), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n643), .B1(new_n361), .B2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n435), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n434), .B1(new_n414), .B2(new_n426), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n304), .B1(new_n647), .B2(new_n651), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n652), .A2(new_n310), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n641), .A2(new_n653), .ZN(G369));
  NAND3_X1  g0454(.A1(new_n258), .A2(new_n217), .A3(G13), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n655), .A2(KEYINPUT27), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(KEYINPUT27), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n656), .A2(G213), .A3(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(G343), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n593), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g0461(.A(new_n661), .B(KEYINPUT86), .ZN(new_n662));
  INV_X1    g0462(.A(new_n617), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT87), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n662), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n617), .A2(KEYINPUT87), .ZN(new_n666));
  INV_X1    g0466(.A(new_n625), .ZN(new_n667));
  AOI22_X1  g0467(.A1(new_n665), .A2(new_n666), .B1(new_n667), .B2(new_n662), .ZN(new_n668));
  INV_X1    g0468(.A(G330), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n660), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n578), .B1(new_n546), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n565), .A2(new_n660), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n667), .A2(new_n672), .ZN(new_n678));
  NOR3_X1   g0478(.A1(new_n678), .A2(new_n577), .A3(new_n565), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n621), .A2(new_n660), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n677), .A2(new_n681), .ZN(G399));
  NAND3_X1  g0482(.A1(new_n212), .A2(KEYINPUT88), .A3(new_n284), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(KEYINPUT88), .B1(new_n212), .B2(new_n284), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n381), .A2(new_n538), .A3(new_n496), .ZN(new_n687));
  NOR3_X1   g0487(.A1(new_n686), .A2(new_n258), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n688), .B1(new_n215), .B2(new_n686), .ZN(new_n689));
  XOR2_X1   g0489(.A(new_n689), .B(KEYINPUT28), .Z(new_n690));
  INV_X1    g0490(.A(KEYINPUT92), .ZN(new_n691));
  INV_X1    g0491(.A(new_n639), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n457), .A2(new_n461), .A3(new_n484), .ZN(new_n693));
  INV_X1    g0493(.A(new_n461), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n442), .B1(new_n402), .B2(new_n405), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(KEYINPUT77), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n696), .A2(new_n443), .A3(new_n451), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n694), .B1(new_n697), .B2(new_n256), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n693), .B1(new_n698), .B2(new_n491), .ZN(new_n699));
  AOI22_X1  g0499(.A1(new_n573), .A2(new_n365), .B1(new_n386), .B2(new_n575), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n630), .B1(new_n700), .B2(new_n569), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n692), .B1(new_n702), .B2(new_n626), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n632), .A2(new_n630), .A3(new_n636), .A4(KEYINPUT26), .ZN(new_n704));
  NOR3_X1   g0504(.A1(new_n698), .A2(new_n491), .A3(new_n523), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n704), .B1(new_n705), .B2(KEYINPUT26), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n660), .B1(new_n703), .B2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT91), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n707), .A2(new_n708), .A3(KEYINPUT29), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n629), .A2(new_n706), .A3(new_n639), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n710), .A2(KEYINPUT29), .A3(new_n672), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(KEYINPUT91), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n640), .A2(new_n672), .ZN(new_n713));
  XOR2_X1   g0513(.A(KEYINPUT90), .B(KEYINPUT29), .Z(new_n714));
  AOI22_X1  g0514(.A1(new_n709), .A2(new_n712), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n524), .A2(new_n617), .A3(new_n578), .A4(new_n672), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n487), .A2(new_n488), .A3(new_n515), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(new_n610), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n718), .A2(new_n563), .A3(KEYINPUT30), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n482), .A2(G179), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n573), .A2(new_n512), .A3(new_n602), .A4(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(KEYINPUT30), .B1(new_n718), .B2(new_n563), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT89), .ZN(new_n723));
  OAI211_X1 g0523(.A(new_n719), .B(new_n721), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT30), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n601), .A2(new_n482), .A3(G179), .A4(new_n515), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n571), .A2(new_n572), .ZN(new_n727));
  OAI211_X1 g0527(.A(new_n723), .B(new_n725), .C1(new_n726), .C2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n660), .B1(new_n724), .B2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT31), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n721), .A2(new_n733), .A3(new_n719), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n734), .A2(KEYINPUT31), .A3(new_n660), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n716), .A2(new_n732), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(G330), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n691), .B1(new_n715), .B2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR3_X1   g0540(.A1(new_n715), .A2(new_n691), .A3(new_n738), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n690), .B1(new_n743), .B2(G1), .ZN(G364));
  AND2_X1   g0544(.A1(new_n217), .A2(G13), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n258), .B1(new_n745), .B2(G45), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n686), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n670), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n665), .A2(new_n666), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n662), .A2(new_n667), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(G330), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(G13), .A2(G33), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(G20), .ZN(new_n757));
  XOR2_X1   g0557(.A(new_n757), .B(KEYINPUT98), .Z(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n668), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n279), .A2(new_n212), .ZN(new_n761));
  INV_X1    g0561(.A(G355), .ZN(new_n762));
  OAI22_X1  g0562(.A1(new_n761), .A2(new_n762), .B1(G116), .B2(new_n212), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n247), .A2(G45), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n275), .A2(new_n212), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n765), .B1(new_n215), .B2(new_n285), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n763), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n216), .B1(G20), .B2(new_n305), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n757), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n748), .B1(new_n767), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n217), .A2(G179), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G190), .A2(G200), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G159), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT94), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n777), .B(KEYINPUT32), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n386), .A2(G200), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n217), .B1(new_n779), .B2(new_n308), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n446), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n772), .A2(new_n386), .A3(G200), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n444), .ZN(new_n783));
  NAND2_X1  g0583(.A1(G20), .A2(G179), .ZN(new_n784));
  XOR2_X1   g0584(.A(new_n784), .B(KEYINPUT93), .Z(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(new_n779), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI211_X1 g0587(.A(new_n781), .B(new_n783), .C1(new_n787), .C2(G58), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n785), .A2(new_n773), .ZN(new_n789));
  OAI211_X1 g0589(.A(new_n778), .B(new_n788), .C1(new_n349), .C2(new_n789), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n772), .A2(G190), .A3(G200), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n279), .B1(new_n791), .B2(new_n222), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT95), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n785), .A2(G200), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n386), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n794), .A2(G190), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n793), .B1(new_n796), .B2(new_n207), .C1(new_n202), .C2(new_n798), .ZN(new_n799));
  OR2_X1    g0599(.A1(new_n774), .A2(KEYINPUT97), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n774), .A2(KEYINPUT97), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n789), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n803), .A2(G329), .B1(new_n804), .B2(G311), .ZN(new_n805));
  INV_X1    g0605(.A(G322), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n805), .B1(new_n806), .B2(new_n786), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n795), .A2(G326), .ZN(new_n808));
  XNOR2_X1  g0608(.A(KEYINPUT33), .B(G317), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n797), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n791), .B(KEYINPUT96), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(G303), .ZN(new_n812));
  INV_X1    g0612(.A(G294), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n275), .B1(new_n780), .B2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n782), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n814), .B1(G283), .B2(new_n815), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n808), .A2(new_n810), .A3(new_n812), .A4(new_n816), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n790), .A2(new_n799), .B1(new_n807), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n771), .B1(new_n818), .B2(new_n768), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n749), .A2(new_n754), .B1(new_n760), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(G396));
  NOR2_X1   g0621(.A1(new_n389), .A2(new_n660), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n377), .A2(new_n660), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n387), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n822), .B1(new_n389), .B2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT99), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(new_n713), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n390), .A2(new_n672), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n829), .B1(new_n703), .B2(new_n638), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n748), .B1(new_n832), .B2(new_n737), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n833), .B1(new_n737), .B2(new_n832), .ZN(new_n834));
  OR2_X1    g0634(.A1(new_n768), .A2(new_n755), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n748), .B1(G77), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(G311), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n802), .A2(new_n837), .B1(new_n789), .B2(new_n538), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n838), .B1(G294), .B2(new_n787), .ZN(new_n839));
  AOI22_X1  g0639(.A1(G283), .A2(new_n797), .B1(new_n795), .B2(G303), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n782), .A2(new_n222), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n275), .B1(new_n780), .B2(new_n446), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n841), .B(new_n842), .C1(new_n811), .C2(G107), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n839), .A2(new_n840), .A3(new_n843), .ZN(new_n844));
  AOI22_X1  g0644(.A1(G143), .A2(new_n787), .B1(new_n804), .B2(G159), .ZN(new_n845));
  INV_X1    g0645(.A(G150), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n845), .B1(new_n846), .B2(new_n798), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n847), .B1(G137), .B2(new_n795), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT34), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n811), .A2(G50), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n279), .B1(new_n782), .B2(new_n202), .ZN(new_n851));
  INV_X1    g0651(.A(new_n780), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n851), .B1(G58), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(G132), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n850), .B(new_n853), .C1(new_n854), .C2(new_n802), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n844), .B1(new_n849), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n836), .B1(new_n856), .B2(new_n768), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n857), .B1(new_n756), .B2(new_n825), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n834), .A2(new_n858), .ZN(new_n859));
  XOR2_X1   g0659(.A(new_n859), .B(KEYINPUT100), .Z(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(G384));
  NAND2_X1  g0661(.A1(new_n715), .A2(new_n440), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n653), .ZN(new_n863));
  OAI22_X1  g0663(.A1(new_n364), .A2(new_n366), .B1(new_n359), .B2(new_n672), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n864), .B1(new_n340), .B2(new_n360), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n360), .A2(new_n660), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n340), .B1(new_n367), .B2(new_n369), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n869), .B1(new_n830), .B2(new_n822), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT38), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT37), .ZN(new_n873));
  OR2_X1    g0673(.A1(new_n411), .A2(new_n202), .ZN(new_n874));
  AOI21_X1  g0674(.A(KEYINPUT16), .B1(new_n874), .B2(new_n408), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n393), .B1(new_n875), .B2(new_n413), .ZN(new_n876));
  INV_X1    g0676(.A(new_n658), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n876), .B1(new_n426), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n873), .B1(new_n878), .B2(new_n436), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n427), .A2(new_n436), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT101), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n414), .A2(new_n881), .A3(new_n877), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n414), .A2(new_n877), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(KEYINPUT101), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n880), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n879), .B1(new_n885), .B2(new_n873), .ZN(new_n886));
  AND2_X1   g0686(.A1(new_n876), .A2(new_n877), .ZN(new_n887));
  AND2_X1   g0687(.A1(new_n439), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n872), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n879), .ZN(new_n890));
  AND3_X1   g0690(.A1(new_n414), .A2(new_n881), .A3(new_n877), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n881), .B1(new_n414), .B2(new_n877), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n427), .B(new_n436), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n890), .B1(new_n893), .B2(KEYINPUT37), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n439), .A2(new_n887), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n894), .A2(KEYINPUT38), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n889), .A2(new_n896), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n871), .A2(new_n897), .B1(new_n651), .B2(new_n658), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n885), .A2(new_n873), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n884), .A2(new_n882), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n900), .B1(new_n650), .B2(new_n642), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n893), .A2(KEYINPUT37), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n872), .B(new_n899), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n896), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT39), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n340), .A2(new_n360), .A3(new_n672), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n889), .A2(KEYINPUT39), .A3(new_n896), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n906), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n898), .A2(new_n910), .ZN(new_n911));
  XOR2_X1   g0711(.A(new_n863), .B(new_n911), .Z(new_n912));
  INV_X1    g0712(.A(new_n340), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n370), .ZN(new_n914));
  INV_X1    g0714(.A(new_n867), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n865), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n825), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI211_X1 g0718(.A(KEYINPUT31), .B(new_n660), .C1(new_n724), .C2(new_n729), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n733), .A2(KEYINPUT89), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n921), .A2(new_n728), .A3(new_n719), .A4(new_n721), .ZN(new_n922));
  AOI21_X1  g0722(.A(KEYINPUT31), .B1(new_n922), .B2(new_n660), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(KEYINPUT102), .B1(new_n924), .B2(new_n716), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n716), .A2(new_n732), .A3(KEYINPUT102), .A4(new_n919), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n918), .B(new_n904), .C1(new_n925), .C2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(KEYINPUT40), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n867), .B1(new_n913), .B2(new_n370), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n825), .B1(new_n930), .B2(new_n865), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n716), .A2(new_n732), .A3(new_n919), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT102), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n931), .B1(new_n934), .B2(new_n926), .ZN(new_n935));
  AOI21_X1  g0735(.A(KEYINPUT40), .B1(new_n889), .B2(new_n896), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n929), .A2(new_n937), .ZN(new_n938));
  AOI211_X1 g0738(.A(new_n439), .B(new_n391), .C1(new_n934), .C2(new_n926), .ZN(new_n939));
  AND2_X1   g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n938), .A2(new_n939), .ZN(new_n941));
  NOR3_X1   g0741(.A1(new_n940), .A2(new_n941), .A3(new_n669), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n912), .A2(new_n942), .B1(new_n258), .B2(new_n745), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n943), .B1(new_n912), .B2(new_n942), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n450), .A2(KEYINPUT35), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n450), .A2(KEYINPUT35), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n945), .A2(G116), .A3(new_n218), .A4(new_n946), .ZN(new_n947));
  XOR2_X1   g0747(.A(new_n947), .B(KEYINPUT36), .Z(new_n948));
  OAI211_X1 g0748(.A(new_n215), .B(G77), .C1(new_n201), .C2(new_n202), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n207), .A2(G68), .ZN(new_n950));
  AOI211_X1 g0750(.A(new_n258), .B(G13), .C1(new_n949), .C2(new_n950), .ZN(new_n951));
  OR3_X1    g0751(.A1(new_n944), .A2(new_n948), .A3(new_n951), .ZN(G367));
  NOR2_X1   g0752(.A1(new_n234), .A2(new_n765), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n769), .B1(new_n212), .B2(new_n373), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n748), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(G317), .ZN(new_n956));
  OAI221_X1 g0756(.A(new_n275), .B1(new_n774), .B2(new_n956), .C1(new_n446), .C2(new_n782), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n957), .B1(new_n442), .B2(new_n852), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n796), .B2(new_n837), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n811), .A2(KEYINPUT46), .A3(G116), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n798), .B2(new_n813), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT46), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n791), .B2(new_n538), .ZN(new_n963));
  INV_X1    g0763(.A(G283), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n963), .B1(new_n786), .B2(new_n599), .C1(new_n964), .C2(new_n789), .ZN(new_n965));
  NOR3_X1   g0765(.A1(new_n959), .A2(new_n961), .A3(new_n965), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n966), .B(KEYINPUT109), .Z(new_n967));
  NAND2_X1  g0767(.A1(new_n852), .A2(G68), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n786), .B2(new_n846), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n969), .B(KEYINPUT110), .Z(new_n970));
  AOI21_X1  g0770(.A(new_n275), .B1(new_n775), .B2(G137), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n971), .B1(new_n201), .B2(new_n791), .C1(new_n349), .C2(new_n782), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n972), .B1(G50), .B2(new_n804), .ZN(new_n973));
  AOI22_X1  g0773(.A1(G143), .A2(new_n795), .B1(new_n797), .B2(G159), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n970), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n967), .A2(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT47), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n955), .B1(new_n977), .B2(new_n768), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n503), .A2(new_n672), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n630), .A2(new_n979), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n980), .A2(KEYINPUT103), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n639), .A2(new_n979), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n980), .A2(KEYINPUT103), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n981), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT104), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n759), .ZN(new_n986));
  AND2_X1   g0786(.A1(new_n978), .A2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n627), .B1(new_n698), .B2(new_n672), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n632), .A2(new_n636), .A3(new_n660), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  NOR3_X1   g0792(.A1(new_n992), .A2(new_n679), .A3(new_n680), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT45), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n681), .A2(new_n991), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT44), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(new_n677), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT106), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n675), .A2(new_n999), .A3(new_n678), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n673), .A2(new_n674), .A3(new_n678), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(KEYINPUT106), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n679), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT107), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n752), .A2(new_n1004), .A3(G330), .ZN(new_n1005));
  OAI21_X1  g0805(.A(KEYINPUT107), .B1(new_n668), .B2(new_n669), .ZN(new_n1006));
  AND3_X1   g0806(.A1(new_n1003), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1005), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n741), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1009), .B1(new_n1010), .B2(new_n739), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n998), .B1(new_n1011), .B2(KEYINPUT108), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n740), .B2(new_n741), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT108), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n743), .B1(new_n1012), .B2(new_n1016), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n686), .B(KEYINPUT41), .Z(new_n1018));
  INV_X1    g0818(.A(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n747), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n991), .A2(new_n679), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT42), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n492), .B1(new_n991), .B2(new_n565), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1023), .A2(new_n660), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT43), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n1022), .A2(new_n1024), .B1(new_n1025), .B2(new_n985), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n985), .A2(new_n1025), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1026), .B(new_n1027), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n677), .A2(new_n992), .ZN(new_n1029));
  AND2_X1   g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n1030), .A2(KEYINPUT105), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1028), .A2(KEYINPUT105), .A3(new_n1029), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n988), .B1(new_n1020), .B2(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT111), .ZN(G387));
  NAND3_X1  g0836(.A1(new_n1010), .A2(new_n1009), .A3(new_n739), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1014), .A2(new_n1037), .A3(new_n686), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n675), .A2(new_n759), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n687), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n1040), .A2(new_n761), .B1(G107), .B2(new_n212), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT112), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n239), .A2(new_n285), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT113), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n285), .B1(new_n202), .B2(new_n349), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n252), .A2(G50), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT114), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n687), .B(new_n1045), .C1(new_n1047), .C2(KEYINPUT50), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n1047), .A2(KEYINPUT50), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n765), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1042), .B1(new_n1044), .B2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n748), .B1(new_n1051), .B2(new_n770), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(G303), .A2(new_n804), .B1(new_n787), .B2(G317), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n806), .B2(new_n796), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(G311), .B2(new_n797), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n1055), .A2(KEYINPUT48), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(KEYINPUT48), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n791), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n852), .A2(G283), .B1(new_n1058), .B2(G294), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1056), .A2(new_n1057), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT49), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n782), .A2(new_n538), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n279), .B(new_n1064), .C1(G326), .C2(new_n775), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1062), .A2(new_n1063), .A3(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n780), .A2(new_n373), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n279), .B1(new_n774), .B2(new_n846), .C1(new_n446), .C2(new_n782), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n1067), .B(new_n1068), .C1(G77), .C2(new_n1058), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(G50), .A2(new_n787), .B1(new_n804), .B2(G68), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(G159), .A2(new_n795), .B1(new_n797), .B2(new_n371), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1066), .A2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1052), .B1(new_n1073), .B2(new_n768), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n1013), .A2(new_n747), .B1(new_n1039), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1038), .A2(new_n1075), .ZN(G393));
  NAND2_X1  g0876(.A1(new_n998), .A2(new_n747), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n244), .A2(new_n765), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n769), .B1(new_n446), .B2(new_n212), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n748), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT115), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n787), .A2(G159), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n796), .B2(new_n846), .ZN(new_n1083));
  XOR2_X1   g0883(.A(new_n1083), .B(KEYINPUT51), .Z(new_n1084));
  AOI211_X1 g0884(.A(new_n275), .B(new_n841), .C1(G143), .C2(new_n775), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n780), .A2(new_n349), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(G68), .B2(new_n1058), .ZN(new_n1087));
  AND2_X1   g0887(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n1088), .B1(new_n207), .B2(new_n798), .C1(new_n252), .C2(new_n789), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1084), .A2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n275), .B1(new_n774), .B2(new_n806), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n780), .A2(new_n538), .B1(new_n791), .B2(new_n964), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n1091), .B(new_n1092), .C1(G107), .C2(new_n815), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1093), .B1(new_n813), .B2(new_n789), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n796), .A2(new_n956), .B1(new_n786), .B2(new_n837), .ZN(new_n1095));
  XOR2_X1   g0895(.A(new_n1095), .B(KEYINPUT52), .Z(new_n1096));
  AOI211_X1 g0896(.A(new_n1094), .B(new_n1096), .C1(G303), .C2(new_n797), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1090), .B1(new_n1098), .B2(KEYINPUT116), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(KEYINPUT116), .B2(new_n1098), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1081), .B1(new_n1100), .B2(new_n768), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n757), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1101), .B1(new_n991), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1077), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n997), .B(new_n676), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT117), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1106), .A2(new_n1014), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1107), .B1(new_n1106), .B2(new_n1014), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n686), .B1(new_n1012), .B2(new_n1016), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1105), .B1(new_n1111), .B2(new_n1112), .ZN(G390));
  INV_X1    g0913(.A(new_n829), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n822), .B1(new_n640), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n669), .B1(new_n934), .B2(new_n926), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n918), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n916), .B1(new_n737), .B2(new_n917), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1115), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(G330), .B1(new_n925), .B2(new_n927), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n827), .B1(new_n1121), .B2(KEYINPUT119), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT119), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1116), .A2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n869), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n738), .A2(new_n825), .A3(new_n869), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n824), .A2(new_n389), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n710), .A2(new_n672), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n822), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1126), .A2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1120), .B1(new_n1125), .B2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n907), .B1(new_n1115), .B2(new_n916), .ZN(new_n1134));
  AND3_X1   g0934(.A1(new_n889), .A2(KEYINPUT39), .A3(new_n896), .ZN(new_n1135));
  AOI21_X1  g0935(.A(KEYINPUT39), .B1(new_n903), .B2(new_n896), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1134), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n916), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n908), .B1(new_n903), .B2(new_n896), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1117), .B1(new_n1137), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT118), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n906), .A2(new_n909), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n1144), .A2(new_n1134), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n1142), .A2(new_n1143), .B1(new_n1145), .B2(new_n1126), .ZN(new_n1146));
  OAI21_X1  g0946(.A(KEYINPUT118), .B1(new_n1145), .B2(new_n1117), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n440), .A2(new_n1116), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n862), .A2(new_n653), .A3(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1133), .A2(new_n1146), .A3(new_n1147), .A4(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n827), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1152), .B1(new_n1116), .B2(new_n1123), .ZN(new_n1153));
  AOI211_X1 g0953(.A(KEYINPUT119), .B(new_n669), .C1(new_n934), .C2(new_n926), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n916), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1132), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1119), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1121), .A2(new_n931), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n906), .A2(new_n909), .B1(new_n870), .B2(new_n907), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n904), .A2(new_n907), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1160), .A2(new_n1138), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1143), .B(new_n1158), .C1(new_n1159), .C2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1137), .A2(new_n1141), .A3(new_n1126), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1137), .A2(new_n1141), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1143), .B1(new_n1165), .B2(new_n1158), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n1157), .A2(new_n1149), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1151), .A2(new_n1167), .A3(new_n686), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1144), .A2(new_n755), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n748), .B1(new_n371), .B2(new_n835), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n802), .A2(new_n813), .B1(new_n789), .B2(new_n446), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(G116), .B2(new_n787), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(G283), .A2(new_n795), .B1(new_n797), .B2(new_n442), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n275), .B1(new_n782), .B2(new_n202), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n1086), .B(new_n1175), .C1(new_n811), .C2(G87), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1173), .A2(new_n1174), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n787), .A2(G132), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT53), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n791), .A2(new_n846), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(KEYINPUT54), .B(G143), .ZN(new_n1181));
  OAI221_X1 g0981(.A(new_n1178), .B1(new_n1179), .B2(new_n1180), .C1(new_n789), .C2(new_n1181), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(G128), .A2(new_n795), .B1(new_n797), .B2(G137), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n782), .A2(new_n207), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n275), .B(new_n1184), .C1(G159), .C2(new_n852), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n803), .A2(G125), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1183), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1177), .B1(new_n1182), .B2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1171), .B1(new_n1188), .B2(new_n768), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n1169), .A2(new_n747), .B1(new_n1170), .B2(new_n1189), .ZN(new_n1190));
  AND3_X1   g0990(.A1(new_n1168), .A2(KEYINPUT120), .A3(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(KEYINPUT120), .B1(new_n1168), .B2(new_n1190), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1191), .A2(new_n1192), .ZN(G378));
  NOR2_X1   g0993(.A1(new_n269), .A2(new_n658), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(new_n304), .B2(new_n310), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n304), .A2(new_n310), .A3(new_n1195), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1199));
  AND3_X1   g0999(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1199), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n938), .B2(G330), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n928), .A2(KEYINPUT40), .B1(new_n935), .B2(new_n936), .ZN(new_n1205));
  NOR3_X1   g1005(.A1(new_n1205), .A2(new_n669), .A3(new_n1202), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n911), .B1(new_n1204), .B2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n938), .A2(G330), .A3(new_n1203), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1202), .B1(new_n1205), .B2(new_n669), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n911), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1208), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1207), .A2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1202), .A2(new_n755), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n748), .B1(G50), .B2(new_n835), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n444), .A2(new_n786), .B1(new_n789), .B2(new_n373), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n815), .A2(G58), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(new_n1216), .B(KEYINPUT122), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1058), .A2(G77), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n279), .A2(G41), .ZN(new_n1219));
  AND4_X1   g1019(.A1(new_n968), .A2(new_n1217), .A3(new_n1218), .A4(new_n1219), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1220), .B1(new_n446), .B2(new_n798), .C1(new_n538), .C2(new_n796), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1215), .B(new_n1221), .C1(G283), .C2(new_n803), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(KEYINPUT58), .ZN(new_n1223));
  AOI211_X1 g1023(.A(G50), .B(new_n1219), .C1(new_n271), .C2(new_n284), .ZN(new_n1224));
  XOR2_X1   g1024(.A(new_n1224), .B(KEYINPUT121), .Z(new_n1225));
  AND2_X1   g1025(.A1(new_n1223), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n787), .A2(G128), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n852), .A2(G150), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1181), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1058), .A2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1227), .A2(new_n1228), .A3(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n795), .A2(G125), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1232), .B1(new_n798), .B2(new_n854), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n1231), .B(new_n1233), .C1(G137), .C2(new_n804), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1235), .A2(KEYINPUT59), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(KEYINPUT59), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n815), .A2(G159), .ZN(new_n1238));
  AOI211_X1 g1038(.A(G33), .B(G41), .C1(new_n775), .C2(G124), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1237), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  OAI221_X1 g1040(.A(new_n1226), .B1(KEYINPUT58), .B2(new_n1222), .C1(new_n1236), .C2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1214), .B1(new_n1241), .B2(new_n768), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n1212), .A2(new_n747), .B1(new_n1213), .B2(new_n1242), .ZN(new_n1243));
  AND3_X1   g1043(.A1(new_n1208), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1210), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1245));
  OAI21_X1  g1045(.A(KEYINPUT57), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1149), .B1(new_n1169), .B2(new_n1133), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n686), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1147), .A2(new_n1163), .A3(new_n1162), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1150), .B1(new_n1249), .B2(new_n1157), .ZN(new_n1250));
  AOI21_X1  g1050(.A(KEYINPUT57), .B1(new_n1250), .B2(new_n1212), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1243), .B1(new_n1248), .B2(new_n1251), .ZN(G375));
  NAND2_X1  g1052(.A1(new_n1121), .A2(KEYINPUT119), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1253), .A2(new_n1152), .A3(new_n1124), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1132), .B1(new_n1254), .B2(new_n916), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1150), .B1(new_n1255), .B2(new_n1119), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1120), .B(new_n1149), .C1(new_n1125), .C2(new_n1132), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1256), .A2(new_n1019), .A3(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n916), .A2(new_n755), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n748), .B1(G68), .B2(new_n835), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n803), .A2(G303), .B1(new_n804), .B2(new_n442), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1261), .B1(new_n964), .B2(new_n786), .ZN(new_n1262));
  AOI211_X1 g1062(.A(new_n279), .B(new_n1067), .C1(G77), .C2(new_n815), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n797), .A2(G116), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n795), .A2(G294), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n811), .A2(G97), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1263), .A2(new_n1264), .A3(new_n1265), .A4(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n795), .A2(G132), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n797), .A2(new_n1229), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n811), .A2(G159), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1217), .A2(new_n1268), .A3(new_n1269), .A4(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n803), .A2(G128), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n787), .A2(G137), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n275), .B1(new_n852), .B2(G50), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n804), .A2(G150), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1272), .A2(new_n1273), .A3(new_n1274), .A4(new_n1275), .ZN(new_n1276));
  OAI22_X1  g1076(.A1(new_n1262), .A2(new_n1267), .B1(new_n1271), .B2(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1260), .B1(new_n1277), .B2(new_n768), .ZN(new_n1278));
  AOI22_X1  g1078(.A1(new_n1133), .A2(new_n747), .B1(new_n1259), .B2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1258), .A2(new_n1279), .ZN(G381));
  NAND3_X1  g1080(.A1(new_n1038), .A2(new_n820), .A3(new_n1075), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(G384), .A2(new_n1281), .ZN(new_n1282));
  XNOR2_X1  g1082(.A(new_n1282), .B(KEYINPUT123), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1168), .A2(new_n1190), .ZN(new_n1284));
  NOR3_X1   g1084(.A1(G390), .A2(new_n1284), .A3(G381), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1212), .A2(new_n747), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1213), .A2(new_n1242), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1250), .A2(new_n1212), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT57), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n686), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1290), .B1(new_n1207), .B2(new_n1211), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1292), .B1(new_n1293), .B2(new_n1250), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1288), .B1(new_n1291), .B2(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1283), .A2(new_n1285), .A3(new_n1295), .ZN(new_n1296));
  OR2_X1    g1096(.A1(G387), .A2(new_n1296), .ZN(G407));
  INV_X1    g1097(.A(new_n1284), .ZN(new_n1298));
  INV_X1    g1098(.A(G213), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1299), .A2(G343), .ZN(new_n1300));
  XOR2_X1   g1100(.A(new_n1300), .B(KEYINPUT124), .Z(new_n1301));
  NAND3_X1  g1101(.A1(new_n1295), .A2(new_n1298), .A3(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(G407), .A2(G213), .A3(new_n1302), .ZN(G409));
  NAND2_X1  g1103(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n746), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1034), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n987), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1112), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1110), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(new_n1108), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1308), .A2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(G393), .A2(G396), .ZN(new_n1312));
  AOI22_X1  g1112(.A1(new_n1311), .A2(new_n1105), .B1(new_n1281), .B2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT111), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1314), .B1(new_n1312), .B2(new_n1281), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(G390), .A2(new_n1315), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1307), .B1(new_n1313), .B2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1312), .A2(new_n1281), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(G390), .A2(new_n1318), .ZN(new_n1319));
  OAI211_X1 g1119(.A(new_n1035), .B(new_n1319), .C1(G390), .C2(new_n1315), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1317), .A2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT125), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT60), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1257), .A2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1325), .A2(KEYINPUT60), .A3(new_n1120), .A4(new_n1149), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1324), .A2(new_n686), .A3(new_n1256), .A4(new_n1326), .ZN(new_n1327));
  AND3_X1   g1127(.A1(new_n1327), .A2(new_n860), .A3(new_n1279), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n860), .B1(new_n1327), .B2(new_n1279), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1322), .B1(new_n1328), .B2(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1327), .A2(new_n1279), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1331), .A2(G384), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1327), .A2(new_n860), .A3(new_n1279), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1332), .A2(KEYINPUT125), .A3(new_n1333), .ZN(new_n1334));
  AND2_X1   g1134(.A1(new_n1300), .A2(G2897), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1335), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1330), .A2(new_n1334), .A3(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT127), .ZN(new_n1338));
  NOR2_X1   g1138(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1339), .A2(G2897), .A3(new_n1301), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1337), .A2(new_n1338), .A3(new_n1340), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1341), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1338), .B1(new_n1337), .B2(new_n1340), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1250), .A2(new_n1212), .A3(new_n1019), .ZN(new_n1344));
  AOI21_X1  g1144(.A(new_n1284), .B1(new_n1243), .B2(new_n1344), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n1345), .B1(G378), .B2(new_n1295), .ZN(new_n1346));
  NOR2_X1   g1146(.A1(new_n1346), .A2(new_n1301), .ZN(new_n1347));
  NOR3_X1   g1147(.A1(new_n1342), .A2(new_n1343), .A3(new_n1347), .ZN(new_n1348));
  INV_X1    g1148(.A(KEYINPUT61), .ZN(new_n1349));
  AND2_X1   g1149(.A1(new_n1330), .A2(new_n1334), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1243), .A2(new_n1344), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1351), .A2(new_n1298), .ZN(new_n1352));
  INV_X1    g1152(.A(KEYINPUT120), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1284), .A2(new_n1353), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1168), .A2(KEYINPUT120), .A3(new_n1190), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1354), .A2(new_n1355), .ZN(new_n1356));
  OAI21_X1  g1156(.A(new_n1352), .B1(new_n1356), .B2(G375), .ZN(new_n1357));
  INV_X1    g1157(.A(KEYINPUT62), .ZN(new_n1358));
  INV_X1    g1158(.A(new_n1300), .ZN(new_n1359));
  NAND4_X1  g1159(.A1(new_n1350), .A2(new_n1357), .A3(new_n1358), .A4(new_n1359), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1330), .A2(new_n1334), .ZN(new_n1361));
  NOR3_X1   g1161(.A1(new_n1346), .A2(new_n1361), .A3(new_n1301), .ZN(new_n1362));
  OAI211_X1 g1162(.A(new_n1349), .B(new_n1360), .C1(new_n1362), .C2(new_n1358), .ZN(new_n1363));
  OAI21_X1  g1163(.A(new_n1321), .B1(new_n1348), .B2(new_n1363), .ZN(new_n1364));
  NAND3_X1  g1164(.A1(new_n1317), .A2(new_n1349), .A3(new_n1320), .ZN(new_n1365));
  AOI21_X1  g1165(.A(new_n1365), .B1(KEYINPUT63), .B2(new_n1362), .ZN(new_n1366));
  NOR3_X1   g1166(.A1(new_n1346), .A2(new_n1361), .A3(new_n1300), .ZN(new_n1367));
  OR2_X1    g1167(.A1(new_n1367), .A2(KEYINPUT63), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1337), .A2(new_n1340), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1369), .A2(KEYINPUT127), .ZN(new_n1370));
  OAI21_X1  g1170(.A(KEYINPUT126), .B1(new_n1346), .B2(new_n1300), .ZN(new_n1371));
  INV_X1    g1171(.A(KEYINPUT126), .ZN(new_n1372));
  NAND3_X1  g1172(.A1(new_n1357), .A2(new_n1372), .A3(new_n1359), .ZN(new_n1373));
  NAND4_X1  g1173(.A1(new_n1370), .A2(new_n1341), .A3(new_n1371), .A4(new_n1373), .ZN(new_n1374));
  NAND3_X1  g1174(.A1(new_n1366), .A2(new_n1368), .A3(new_n1374), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(new_n1364), .A2(new_n1375), .ZN(G405));
  NAND2_X1  g1176(.A1(G378), .A2(new_n1295), .ZN(new_n1377));
  NAND2_X1  g1177(.A1(G375), .A2(new_n1298), .ZN(new_n1378));
  NAND2_X1  g1178(.A1(new_n1377), .A2(new_n1378), .ZN(new_n1379));
  NOR2_X1   g1179(.A1(new_n1379), .A2(new_n1339), .ZN(new_n1380));
  AOI21_X1  g1180(.A(new_n1380), .B1(new_n1361), .B2(new_n1379), .ZN(new_n1381));
  XNOR2_X1  g1181(.A(new_n1381), .B(new_n1321), .ZN(G402));
endmodule


