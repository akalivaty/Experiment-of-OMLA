//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 0 0 0 0 0 0 0 1 0 1 0 0 1 0 1 0 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 1 1 0 0 0 0 0 0 0 1 0 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:45 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n208,
    new_n209, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1197, new_n1198, new_n1199, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1265, new_n1266, new_n1267, new_n1268;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0007(.A1(G97), .A2(G107), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n209), .A2(G87), .ZN(G355));
  NAND2_X1  g0010(.A1(new_n206), .A2(G50), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT67), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(KEYINPUT66), .ZN(new_n214));
  INV_X1    g0014(.A(KEYINPUT66), .ZN(new_n215));
  NAND3_X1  g0015(.A1(new_n215), .A2(G1), .A3(G13), .ZN(new_n216));
  AND2_X1   g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(G20), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n212), .A2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(KEYINPUT1), .ZN(new_n221));
  INV_X1    g0021(.A(G1), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n222), .A2(new_n218), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT68), .Z(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n228));
  AND3_X1   g0028(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n223), .B1(new_n225), .B2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n220), .B1(new_n221), .B2(new_n230), .ZN(new_n231));
  INV_X1    g0031(.A(G13), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n223), .A2(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  OAI211_X1 g0034(.A(new_n234), .B(G250), .C1(G257), .C2(G264), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n235), .B(KEYINPUT65), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT0), .ZN(new_n237));
  AOI211_X1 g0037(.A(new_n231), .B(new_n237), .C1(new_n221), .C2(new_n230), .ZN(G361));
  XOR2_X1   g0038(.A(G238), .B(G244), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G232), .ZN(new_n240));
  XOR2_X1   g0040(.A(KEYINPUT2), .B(G226), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G264), .B(G270), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G358));
  XNOR2_X1  g0046(.A(G50), .B(G68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n247), .B(new_n248), .Z(new_n249));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XOR2_X1   g0050(.A(G107), .B(G116), .Z(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n249), .B(new_n252), .Z(G351));
  INV_X1    g0053(.A(KEYINPUT18), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n218), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G159), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G58), .A2(G68), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n203), .A2(new_n205), .A3(new_n259), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n258), .B1(new_n260), .B2(G20), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT3), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G33), .ZN(new_n264));
  AOI21_X1  g0064(.A(G20), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT7), .ZN(new_n266));
  OAI21_X1  g0066(.A(G68), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n262), .A2(new_n264), .ZN(new_n268));
  XNOR2_X1  g0068(.A(KEYINPUT75), .B(KEYINPUT7), .ZN(new_n269));
  AND3_X1   g0069(.A1(new_n268), .A2(new_n269), .A3(new_n218), .ZN(new_n270));
  OAI211_X1 g0070(.A(KEYINPUT16), .B(new_n261), .C1(new_n267), .C2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n223), .A2(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n217), .A2(new_n272), .ZN(new_n273));
  AND2_X1   g0073(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT16), .ZN(new_n275));
  XNOR2_X1  g0075(.A(KEYINPUT3), .B(G33), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n269), .B1(new_n276), .B2(G20), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n268), .A2(KEYINPUT7), .A3(new_n218), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n202), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n260), .A2(G20), .ZN(new_n280));
  INV_X1    g0080(.A(new_n258), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n275), .B1(new_n279), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(KEYINPUT76), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT76), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n285), .B(new_n275), .C1(new_n279), .C2(new_n282), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n274), .A2(new_n284), .A3(new_n286), .ZN(new_n287));
  NOR3_X1   g0087(.A1(new_n232), .A2(new_n218), .A3(G1), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n217), .A2(new_n289), .A3(new_n272), .ZN(new_n290));
  XNOR2_X1  g0090(.A(KEYINPUT8), .B(G58), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n222), .A2(G20), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  OAI22_X1  g0094(.A1(new_n290), .A2(new_n294), .B1(new_n289), .B2(new_n292), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT77), .ZN(new_n296));
  XNOR2_X1  g0096(.A(new_n295), .B(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n287), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(G33), .A2(G41), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n299), .A2(G1), .A3(G13), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n222), .B1(G41), .B2(G45), .ZN(new_n301));
  AND3_X1   g0101(.A1(new_n300), .A2(G232), .A3(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT69), .ZN(new_n303));
  AND2_X1   g0103(.A1(G33), .A2(G41), .ZN(new_n304));
  OAI21_X1  g0104(.A(G274), .B1(new_n304), .B2(new_n213), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n303), .B1(new_n305), .B2(new_n301), .ZN(new_n306));
  INV_X1    g0106(.A(new_n301), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n307), .A2(new_n300), .A3(KEYINPUT69), .A4(G274), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n302), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n262), .A2(new_n264), .A3(G226), .A4(G1698), .ZN(new_n310));
  INV_X1    g0110(.A(G1698), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n262), .A2(new_n264), .A3(G223), .A4(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(G33), .A2(G87), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n310), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n304), .B1(new_n214), .B2(new_n216), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AND3_X1   g0116(.A1(new_n309), .A2(G179), .A3(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G169), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n318), .B1(new_n309), .B2(new_n316), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n254), .B1(new_n298), .B2(new_n321), .ZN(new_n322));
  AOI211_X1 g0122(.A(KEYINPUT18), .B(new_n320), .C1(new_n287), .C2(new_n297), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g0124(.A(new_n295), .B(KEYINPUT77), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n271), .A2(new_n273), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n326), .B1(KEYINPUT76), .B2(new_n283), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n325), .B1(new_n327), .B2(new_n286), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT79), .ZN(new_n329));
  AOI21_X1  g0129(.A(G200), .B1(new_n309), .B2(new_n316), .ZN(new_n330));
  INV_X1    g0130(.A(G190), .ZN(new_n331));
  AND3_X1   g0131(.A1(new_n309), .A2(new_n331), .A3(new_n316), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT78), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n330), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n306), .A2(new_n308), .ZN(new_n335));
  INV_X1    g0135(.A(new_n302), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n316), .A2(new_n335), .A3(new_n331), .A4(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(KEYINPUT78), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n329), .B1(new_n334), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n309), .A2(new_n316), .ZN(new_n340));
  INV_X1    g0140(.A(G200), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n309), .A2(new_n333), .A3(new_n316), .A4(new_n331), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n338), .A2(new_n342), .A3(new_n329), .A4(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n328), .B1(new_n339), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT17), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n338), .A2(new_n342), .A3(new_n343), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(KEYINPUT79), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n344), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n351), .A2(KEYINPUT17), .A3(new_n328), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n324), .A2(new_n348), .A3(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n293), .A2(G50), .ZN(new_n355));
  OAI22_X1  g0155(.A1(new_n290), .A2(new_n355), .B1(G50), .B2(new_n289), .ZN(new_n356));
  XNOR2_X1  g0156(.A(new_n356), .B(KEYINPUT70), .ZN(new_n357));
  OAI21_X1  g0157(.A(G20), .B1(new_n206), .B2(G50), .ZN(new_n358));
  INV_X1    g0158(.A(G150), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n218), .A2(G33), .ZN(new_n360));
  OAI221_X1 g0160(.A(new_n358), .B1(new_n359), .B2(new_n256), .C1(new_n291), .C2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n273), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n357), .A2(new_n362), .ZN(new_n363));
  XOR2_X1   g0163(.A(new_n363), .B(KEYINPUT9), .Z(new_n364));
  NOR2_X1   g0164(.A1(new_n268), .A2(G1698), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(G222), .ZN(new_n366));
  INV_X1    g0166(.A(G77), .ZN(new_n367));
  INV_X1    g0167(.A(G223), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n276), .A2(G1698), .ZN(new_n369));
  OAI221_X1 g0169(.A(new_n366), .B1(new_n367), .B2(new_n276), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n315), .ZN(new_n371));
  INV_X1    g0171(.A(new_n335), .ZN(new_n372));
  AND2_X1   g0172(.A1(new_n300), .A2(new_n301), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n372), .B1(G226), .B2(new_n373), .ZN(new_n374));
  AND2_X1   g0174(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(KEYINPUT72), .B1(new_n375), .B2(G190), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n376), .B1(new_n341), .B2(new_n375), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n364), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT10), .ZN(new_n379));
  XNOR2_X1  g0179(.A(new_n378), .B(new_n379), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n375), .A2(G169), .ZN(new_n381));
  INV_X1    g0181(.A(G179), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n381), .B1(new_n382), .B2(new_n375), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n363), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n380), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(G238), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n387), .B1(new_n373), .B2(KEYINPUT73), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(KEYINPUT73), .B2(new_n373), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n276), .A2(G232), .A3(G1698), .ZN(new_n390));
  NAND2_X1  g0190(.A1(G33), .A2(G97), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n276), .A2(new_n311), .ZN(new_n392));
  INV_X1    g0192(.A(G226), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n390), .B(new_n391), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(new_n315), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n389), .A2(new_n395), .A3(new_n335), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(KEYINPUT13), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n396), .A2(KEYINPUT13), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(KEYINPUT14), .B1(new_n400), .B2(new_n318), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(G179), .ZN(new_n402));
  INV_X1    g0202(.A(new_n399), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n397), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT14), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n404), .A2(new_n405), .A3(G169), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n401), .A2(new_n402), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(KEYINPUT74), .B1(new_n288), .B2(new_n202), .ZN(new_n408));
  XNOR2_X1  g0208(.A(new_n408), .B(KEYINPUT12), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n202), .A2(G20), .ZN(new_n410));
  INV_X1    g0210(.A(G50), .ZN(new_n411));
  OAI221_X1 g0211(.A(new_n410), .B1(new_n360), .B2(new_n367), .C1(new_n411), .C2(new_n256), .ZN(new_n412));
  AND2_X1   g0212(.A1(new_n273), .A2(new_n412), .ZN(new_n413));
  OR2_X1    g0213(.A1(new_n413), .A2(KEYINPUT11), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(KEYINPUT11), .ZN(new_n415));
  INV_X1    g0215(.A(new_n290), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n416), .A2(G68), .A3(new_n293), .ZN(new_n417));
  AND4_X1   g0217(.A1(new_n409), .A2(new_n414), .A3(new_n415), .A4(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n407), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n418), .B1(new_n404), .B2(new_n331), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n400), .A2(new_n341), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n420), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n416), .A2(G77), .A3(new_n293), .ZN(new_n427));
  XOR2_X1   g0227(.A(new_n427), .B(KEYINPUT71), .Z(new_n428));
  NAND2_X1  g0228(.A1(G20), .A2(G77), .ZN(new_n429));
  XNOR2_X1  g0229(.A(KEYINPUT15), .B(G87), .ZN(new_n430));
  OAI221_X1 g0230(.A(new_n429), .B1(new_n291), .B2(new_n256), .C1(new_n360), .C2(new_n430), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n431), .A2(new_n273), .B1(new_n367), .B2(new_n288), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n372), .B1(G244), .B2(new_n373), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n276), .A2(G232), .A3(new_n311), .ZN(new_n435));
  INV_X1    g0235(.A(G107), .ZN(new_n436));
  OAI221_X1 g0236(.A(new_n435), .B1(new_n436), .B2(new_n276), .C1(new_n369), .C2(new_n387), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(new_n315), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(new_n382), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n439), .A2(new_n318), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n433), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n428), .B(new_n432), .C1(new_n331), .C2(new_n439), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n440), .A2(new_n341), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  AND4_X1   g0248(.A1(new_n354), .A2(new_n386), .A3(new_n426), .A4(new_n448), .ZN(new_n449));
  XNOR2_X1  g0249(.A(KEYINPUT5), .B(G41), .ZN(new_n450));
  INV_X1    g0250(.A(G45), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n451), .A2(G1), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n453), .A2(new_n305), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n453), .A2(new_n300), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n454), .B1(new_n455), .B2(G264), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n276), .A2(G257), .A3(G1698), .ZN(new_n457));
  NAND2_X1  g0257(.A1(G33), .A2(G294), .ZN(new_n458));
  INV_X1    g0258(.A(G250), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n457), .B(new_n458), .C1(new_n392), .C2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(new_n315), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n456), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(G169), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n463), .B(KEYINPUT84), .C1(new_n382), .C2(new_n462), .ZN(new_n464));
  OR3_X1    g0264(.A1(new_n462), .A2(KEYINPUT84), .A3(new_n382), .ZN(new_n465));
  INV_X1    g0265(.A(new_n273), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT24), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n276), .A2(new_n218), .A3(G87), .ZN(new_n468));
  XNOR2_X1  g0268(.A(new_n468), .B(KEYINPUT22), .ZN(new_n469));
  INV_X1    g0269(.A(G116), .ZN(new_n470));
  NOR3_X1   g0270(.A1(new_n255), .A2(new_n470), .A3(G20), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT23), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n472), .B1(new_n218), .B2(G107), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n436), .A2(KEYINPUT23), .A3(G20), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n471), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n467), .B1(new_n469), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n469), .A2(new_n467), .A3(new_n475), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n466), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n290), .B1(new_n222), .B2(G33), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT25), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n481), .B1(new_n289), .B2(G107), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n288), .A2(KEYINPUT25), .A3(new_n436), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n480), .A2(G107), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n464), .B(new_n465), .C1(new_n479), .C2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n478), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n273), .B1(new_n487), .B2(new_n476), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n456), .A2(new_n461), .A3(G190), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n462), .A2(G200), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n488), .A2(new_n484), .A3(new_n489), .A4(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n486), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(KEYINPUT85), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT85), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n486), .A2(new_n494), .A3(new_n491), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(G244), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(G1698), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n498), .B1(G238), .B2(G1698), .ZN(new_n499));
  OAI22_X1  g0299(.A1(new_n499), .A2(new_n268), .B1(new_n255), .B2(new_n470), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n315), .ZN(new_n501));
  INV_X1    g0301(.A(G274), .ZN(new_n502));
  INV_X1    g0302(.A(new_n213), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n502), .B1(new_n503), .B2(new_n299), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n459), .B1(new_n222), .B2(G45), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n504), .A2(new_n452), .B1(new_n300), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n501), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n318), .ZN(new_n508));
  NOR2_X1   g0308(.A1(G238), .A2(G1698), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n509), .B1(new_n497), .B2(G1698), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n510), .A2(new_n276), .B1(G33), .B2(G116), .ZN(new_n511));
  INV_X1    g0311(.A(new_n315), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n506), .B(new_n382), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(KEYINPUT80), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT80), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n501), .A2(new_n515), .A3(new_n382), .A4(new_n506), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n508), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT81), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n508), .A2(new_n514), .A3(KEYINPUT81), .A4(new_n516), .ZN(new_n520));
  INV_X1    g0320(.A(new_n430), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n480), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT19), .ZN(new_n523));
  INV_X1    g0323(.A(G97), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n523), .B1(new_n360), .B2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT82), .ZN(new_n526));
  XNOR2_X1  g0326(.A(new_n525), .B(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n276), .A2(new_n218), .A3(G68), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n218), .B1(new_n391), .B2(new_n523), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n529), .B1(G87), .B2(new_n209), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n273), .B1(new_n527), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n430), .A2(new_n288), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n522), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n519), .A2(new_n520), .A3(new_n534), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n416), .B(G87), .C1(G1), .C2(new_n255), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n536), .A2(new_n532), .A3(new_n533), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  AND2_X1   g0338(.A1(new_n501), .A2(new_n506), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(G190), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n507), .A2(G200), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n538), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n535), .A2(KEYINPUT83), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(KEYINPUT83), .B1(new_n535), .B2(new_n542), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT6), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n524), .A2(new_n436), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n546), .B1(new_n547), .B2(new_n208), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n436), .A2(KEYINPUT6), .A3(G97), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(G20), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(new_n367), .B2(new_n256), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n436), .B1(new_n277), .B2(new_n278), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n273), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n289), .A2(G97), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n555), .B1(new_n480), .B2(G97), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n365), .A2(KEYINPUT4), .A3(G244), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT4), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n559), .B1(new_n392), .B2(new_n497), .ZN(new_n560));
  NAND2_X1  g0360(.A1(G33), .A2(G283), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n276), .A2(G250), .A3(G1698), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n558), .A2(new_n560), .A3(new_n561), .A4(new_n562), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n563), .A2(new_n315), .B1(G257), .B2(new_n455), .ZN(new_n564));
  INV_X1    g0364(.A(new_n454), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n557), .B1(G200), .B2(new_n566), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n567), .B1(new_n331), .B2(new_n566), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n566), .A2(new_n318), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n564), .A2(new_n382), .A3(new_n565), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n569), .A2(new_n570), .A3(new_n557), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n480), .A2(G116), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n288), .A2(new_n470), .ZN(new_n574));
  AOI21_X1  g0374(.A(G20), .B1(new_n255), .B2(G97), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n575), .A2(new_n561), .B1(G20), .B2(new_n470), .ZN(new_n576));
  AOI21_X1  g0376(.A(KEYINPUT20), .B1(new_n273), .B2(new_n576), .ZN(new_n577));
  AND3_X1   g0377(.A1(new_n273), .A2(KEYINPUT20), .A3(new_n576), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n573), .B(new_n574), .C1(new_n577), .C2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n276), .A2(G257), .A3(new_n311), .ZN(new_n581));
  INV_X1    g0381(.A(G303), .ZN(new_n582));
  INV_X1    g0382(.A(G264), .ZN(new_n583));
  OAI221_X1 g0383(.A(new_n581), .B1(new_n582), .B2(new_n276), .C1(new_n369), .C2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n315), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n454), .B1(new_n455), .B2(G270), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(G200), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n580), .B(new_n588), .C1(new_n331), .C2(new_n587), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT21), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n587), .A2(G169), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n590), .B1(new_n580), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n585), .A2(G179), .A3(new_n586), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n579), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n579), .A2(KEYINPUT21), .A3(G169), .A4(new_n587), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n589), .A2(new_n592), .A3(new_n595), .A4(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n572), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n449), .A2(new_n496), .A3(new_n545), .A4(new_n598), .ZN(new_n599));
  XOR2_X1   g0399(.A(new_n599), .B(KEYINPUT86), .Z(G372));
  OAI21_X1  g0400(.A(new_n420), .B1(new_n423), .B2(new_n443), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n601), .A2(new_n348), .A3(new_n352), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n324), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n603), .A2(new_n380), .B1(new_n363), .B2(new_n383), .ZN(new_n604));
  INV_X1    g0404(.A(new_n449), .ZN(new_n605));
  NOR3_X1   g0405(.A1(new_n543), .A2(new_n544), .A3(new_n571), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT26), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n596), .A2(new_n595), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n609), .A2(new_n486), .A3(new_n592), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  AND2_X1   g0411(.A1(new_n508), .A2(new_n513), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n534), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n542), .A2(new_n613), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n568), .A2(new_n614), .A3(new_n491), .A4(new_n571), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n571), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n617), .A2(new_n607), .A3(new_n614), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n613), .ZN(new_n619));
  NOR3_X1   g0419(.A1(new_n608), .A2(new_n616), .A3(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n604), .B1(new_n605), .B2(new_n620), .ZN(G369));
  NAND3_X1  g0421(.A1(new_n222), .A2(new_n218), .A3(G13), .ZN(new_n622));
  OR2_X1    g0422(.A1(new_n622), .A2(KEYINPUT27), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(KEYINPUT27), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n623), .A2(G213), .A3(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(G343), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n627), .B1(new_n609), .B2(new_n592), .ZN(new_n628));
  INV_X1    g0428(.A(new_n486), .ZN(new_n629));
  INV_X1    g0429(.A(new_n627), .ZN(new_n630));
  AOI22_X1  g0430(.A1(new_n496), .A2(new_n628), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n627), .B1(new_n479), .B2(new_n485), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n496), .A2(new_n632), .B1(new_n629), .B2(new_n627), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n609), .A2(new_n592), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n580), .A2(new_n630), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n636), .B1(new_n597), .B2(new_n635), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(G330), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n631), .B1(new_n633), .B2(new_n638), .ZN(new_n639));
  XNOR2_X1  g0439(.A(new_n639), .B(KEYINPUT87), .ZN(G399));
  NOR2_X1   g0440(.A1(new_n233), .A2(G41), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  NOR3_X1   g0442(.A1(new_n209), .A2(G87), .A3(G116), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n642), .A2(G1), .A3(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n644), .B1(new_n211), .B2(new_n642), .ZN(new_n645));
  XNOR2_X1  g0445(.A(new_n645), .B(KEYINPUT28), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n496), .A2(new_n545), .A3(new_n598), .A4(new_n630), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n563), .A2(new_n315), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n455), .A2(G257), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n539), .A2(new_n461), .A3(new_n456), .ZN(new_n651));
  NOR3_X1   g0451(.A1(new_n650), .A2(new_n651), .A3(new_n593), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT88), .ZN(new_n653));
  OAI21_X1  g0453(.A(KEYINPUT30), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT30), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n651), .A2(new_n593), .ZN(new_n656));
  OAI211_X1 g0456(.A(KEYINPUT88), .B(new_n655), .C1(new_n656), .C2(new_n650), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n539), .A2(G179), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n566), .A2(new_n462), .A3(new_n587), .A4(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n654), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  AND3_X1   g0460(.A1(new_n660), .A2(KEYINPUT31), .A3(new_n627), .ZN(new_n661));
  AOI21_X1  g0461(.A(KEYINPUT31), .B1(new_n660), .B2(new_n627), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n647), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(G330), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n616), .A2(new_n619), .ZN(new_n667));
  INV_X1    g0467(.A(new_n608), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n627), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  OR2_X1    g0469(.A1(new_n669), .A2(KEYINPUT29), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT89), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n671), .B1(new_n606), .B2(KEYINPUT26), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n617), .A2(KEYINPUT26), .A3(new_n614), .ZN(new_n673));
  INV_X1    g0473(.A(new_n544), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n535), .A2(KEYINPUT83), .A3(new_n542), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(new_n675), .A3(new_n617), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n676), .A2(KEYINPUT89), .A3(new_n607), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n672), .A2(new_n673), .A3(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n613), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT90), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n680), .B1(new_n611), .B2(new_n615), .ZN(new_n681));
  INV_X1    g0481(.A(new_n572), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n614), .A2(new_n491), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n682), .A2(new_n683), .A3(new_n610), .A4(KEYINPUT90), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n679), .B1(new_n681), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n678), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n686), .A2(KEYINPUT29), .A3(new_n630), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n666), .B1(new_n670), .B2(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n646), .B1(new_n688), .B2(G1), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n689), .B(KEYINPUT91), .ZN(G364));
  NOR2_X1   g0490(.A1(new_n232), .A2(G20), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n222), .B1(new_n691), .B2(G45), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n641), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n234), .A2(G116), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n233), .A2(new_n276), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n249), .B2(new_n451), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n697), .B1(new_n451), .B2(new_n212), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n233), .A2(new_n268), .ZN(new_n699));
  AOI211_X1 g0499(.A(new_n695), .B(new_n698), .C1(G355), .C2(new_n699), .ZN(new_n700));
  NOR3_X1   g0500(.A1(G13), .A2(G20), .A3(G33), .ZN(new_n701));
  XNOR2_X1  g0501(.A(new_n701), .B(KEYINPUT92), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n217), .B1(G20), .B2(new_n318), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n694), .B1(new_n700), .B2(new_n706), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n707), .A2(KEYINPUT93), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n218), .A2(new_n331), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n341), .A2(G179), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(G87), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n276), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  XOR2_X1   g0513(.A(new_n713), .B(KEYINPUT95), .Z(new_n714));
  NOR2_X1   g0514(.A1(new_n382), .A2(G200), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n709), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n218), .A2(G190), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(new_n710), .ZN(new_n718));
  OAI22_X1  g0518(.A1(new_n716), .A2(new_n201), .B1(new_n718), .B2(new_n436), .ZN(new_n719));
  NAND3_X1  g0519(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(G190), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n719), .B1(G68), .B2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT94), .ZN(new_n723));
  AND3_X1   g0523(.A1(new_n715), .A2(new_n717), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n723), .B1(new_n715), .B2(new_n717), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  OAI211_X1 g0526(.A(new_n714), .B(new_n722), .C1(new_n367), .C2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(G179), .A2(G200), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n717), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(new_n257), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n730), .B(KEYINPUT32), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n720), .A2(new_n331), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n218), .B1(new_n728), .B2(G190), .ZN(new_n734));
  OAI221_X1 g0534(.A(new_n731), .B1(new_n411), .B2(new_n733), .C1(new_n524), .C2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n716), .ZN(new_n736));
  XNOR2_X1  g0536(.A(KEYINPUT33), .B(G317), .ZN(new_n737));
  AOI22_X1  g0537(.A1(new_n736), .A2(G322), .B1(new_n721), .B2(new_n737), .ZN(new_n738));
  XOR2_X1   g0538(.A(new_n738), .B(KEYINPUT96), .Z(new_n739));
  INV_X1    g0539(.A(new_n726), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G311), .ZN(new_n741));
  INV_X1    g0541(.A(new_n718), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n276), .B1(new_n742), .B2(G283), .ZN(new_n743));
  INV_X1    g0543(.A(new_n711), .ZN(new_n744));
  INV_X1    g0544(.A(new_n729), .ZN(new_n745));
  AOI22_X1  g0545(.A1(G303), .A2(new_n744), .B1(new_n745), .B2(G329), .ZN(new_n746));
  INV_X1    g0546(.A(new_n734), .ZN(new_n747));
  AOI22_X1  g0547(.A1(new_n747), .A2(G294), .B1(G326), .B2(new_n732), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n741), .A2(new_n743), .A3(new_n746), .A4(new_n748), .ZN(new_n749));
  OAI22_X1  g0549(.A1(new_n727), .A2(new_n735), .B1(new_n739), .B2(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n708), .B1(new_n704), .B2(new_n750), .ZN(new_n751));
  OAI221_X1 g0551(.A(new_n751), .B1(KEYINPUT93), .B2(new_n707), .C1(new_n637), .C2(new_n702), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n637), .A2(G330), .ZN(new_n753));
  INV_X1    g0553(.A(new_n694), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n638), .A2(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n752), .B1(new_n753), .B2(new_n755), .ZN(G396));
  INV_X1    g0556(.A(new_n704), .ZN(new_n757));
  INV_X1    g0557(.A(new_n721), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n359), .ZN(new_n759));
  INV_X1    g0559(.A(G137), .ZN(new_n760));
  INV_X1    g0560(.A(G143), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n733), .A2(new_n760), .B1(new_n716), .B2(new_n761), .ZN(new_n762));
  AOI211_X1 g0562(.A(new_n759), .B(new_n762), .C1(G159), .C2(new_n740), .ZN(new_n763));
  AND2_X1   g0563(.A1(new_n763), .A2(KEYINPUT34), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n763), .A2(KEYINPUT34), .ZN(new_n765));
  INV_X1    g0565(.A(G132), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n276), .B1(new_n729), .B2(new_n766), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n767), .B(KEYINPUT98), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n742), .A2(G68), .ZN(new_n769));
  OAI221_X1 g0569(.A(new_n769), .B1(new_n411), .B2(new_n711), .C1(new_n201), .C2(new_n734), .ZN(new_n770));
  OR4_X1    g0570(.A1(new_n764), .A2(new_n765), .A3(new_n768), .A4(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n734), .A2(new_n524), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n733), .A2(new_n582), .ZN(new_n773));
  AOI211_X1 g0573(.A(new_n772), .B(new_n773), .C1(G283), .C2(new_n721), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n268), .B1(new_n711), .B2(new_n436), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT97), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n740), .A2(G116), .ZN(new_n777));
  INV_X1    g0577(.A(G294), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n716), .A2(new_n778), .B1(new_n718), .B2(new_n712), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n779), .B1(G311), .B2(new_n745), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n774), .A2(new_n776), .A3(new_n777), .A4(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n757), .B1(new_n771), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(G13), .A2(G33), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n704), .A2(new_n783), .ZN(new_n784));
  AOI211_X1 g0584(.A(new_n754), .B(new_n782), .C1(new_n367), .C2(new_n784), .ZN(new_n785));
  XOR2_X1   g0585(.A(new_n785), .B(KEYINPUT99), .Z(new_n786));
  INV_X1    g0586(.A(new_n783), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n433), .A2(new_n627), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n788), .B1(new_n445), .B2(new_n446), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(new_n443), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n444), .A2(new_n630), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n786), .B1(new_n787), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n669), .A2(new_n793), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(KEYINPUT100), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n669), .A2(new_n793), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(new_n666), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n754), .B1(new_n798), .B2(new_n666), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n794), .B1(new_n800), .B2(new_n801), .ZN(G384));
  OR2_X1    g0602(.A1(new_n550), .A2(KEYINPUT35), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n550), .A2(KEYINPUT35), .ZN(new_n804));
  NAND4_X1  g0604(.A1(new_n803), .A2(G116), .A3(new_n219), .A4(new_n804), .ZN(new_n805));
  XOR2_X1   g0605(.A(new_n805), .B(KEYINPUT36), .Z(new_n806));
  NAND4_X1  g0606(.A1(new_n206), .A2(G50), .A3(G77), .A4(new_n259), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n411), .A2(G68), .ZN(new_n808));
  AOI211_X1 g0608(.A(new_n222), .B(G13), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n407), .A2(new_n419), .A3(new_n630), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT39), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT38), .ZN(new_n814));
  INV_X1    g0614(.A(new_n625), .ZN(new_n815));
  INV_X1    g0615(.A(new_n295), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n261), .B1(new_n267), .B2(new_n270), .ZN(new_n817));
  AND2_X1   g0617(.A1(new_n817), .A2(new_n275), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n816), .B1(new_n818), .B2(new_n326), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n353), .A2(new_n815), .A3(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT37), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n287), .A2(new_n297), .B1(new_n320), .B2(new_n625), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n346), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT101), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n823), .B1(new_n351), .B2(new_n328), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n828), .A2(KEYINPUT101), .A3(new_n822), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n320), .A2(new_n625), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(new_n819), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n346), .A2(new_n831), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n827), .A2(new_n829), .B1(KEYINPUT37), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n814), .B1(new_n821), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n832), .A2(KEYINPUT37), .ZN(new_n835));
  AND4_X1   g0635(.A1(KEYINPUT101), .A2(new_n346), .A3(new_n822), .A4(new_n824), .ZN(new_n836));
  AOI21_X1  g0636(.A(KEYINPUT101), .B1(new_n828), .B2(new_n822), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n835), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n838), .A2(KEYINPUT38), .A3(new_n820), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n834), .A2(KEYINPUT102), .A3(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT102), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n841), .B(new_n814), .C1(new_n821), .C2(new_n833), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n813), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n353), .A2(new_n298), .A3(new_n815), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT103), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g0646(.A1(new_n353), .A2(KEYINPUT103), .A3(new_n298), .A4(new_n815), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n827), .A2(new_n829), .ZN(new_n848));
  OR2_X1    g0648(.A1(new_n828), .A2(new_n822), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n846), .A2(new_n847), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(new_n814), .ZN(new_n852));
  AOI21_X1  g0652(.A(KEYINPUT39), .B1(new_n852), .B2(new_n839), .ZN(new_n853));
  NOR3_X1   g0653(.A1(new_n843), .A2(new_n853), .A3(KEYINPUT104), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT104), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n839), .A2(KEYINPUT102), .ZN(new_n856));
  AOI21_X1  g0656(.A(KEYINPUT38), .B1(new_n838), .B2(new_n820), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n842), .ZN(new_n859));
  OAI21_X1  g0659(.A(KEYINPUT39), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n844), .A2(new_n845), .B1(new_n848), .B2(new_n849), .ZN(new_n861));
  AOI21_X1  g0661(.A(KEYINPUT38), .B1(new_n861), .B2(new_n847), .ZN(new_n862));
  AND3_X1   g0662(.A1(new_n838), .A2(KEYINPUT38), .A3(new_n820), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n813), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n855), .B1(new_n860), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n812), .B1(new_n854), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n795), .A2(new_n791), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n419), .A2(new_n627), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n420), .A2(new_n424), .A3(new_n868), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n419), .B(new_n627), .C1(new_n407), .C2(new_n423), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n867), .A2(new_n842), .A3(new_n840), .A4(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n625), .B1(new_n322), .B2(new_n323), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n866), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n449), .A2(new_n670), .A3(new_n687), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n604), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n876), .B(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n863), .B1(new_n851), .B2(new_n814), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n647), .A2(new_n663), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n792), .B1(new_n869), .B2(new_n870), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n881), .A2(new_n882), .A3(KEYINPUT40), .ZN(new_n883));
  OAI21_X1  g0683(.A(KEYINPUT105), .B1(new_n880), .B2(new_n883), .ZN(new_n884));
  AND3_X1   g0684(.A1(new_n881), .A2(new_n882), .A3(KEYINPUT40), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT105), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n885), .B(new_n886), .C1(new_n863), .C2(new_n862), .ZN(new_n887));
  AND2_X1   g0687(.A1(new_n881), .A2(new_n882), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n840), .A2(new_n888), .A3(new_n842), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT40), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n884), .A2(new_n887), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(new_n605), .B2(new_n664), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n891), .A2(new_n449), .A3(new_n881), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n893), .A2(G330), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n879), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n896), .B1(new_n222), .B2(new_n691), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n879), .A2(new_n895), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n810), .B1(new_n897), .B2(new_n898), .ZN(G367));
  AOI21_X1  g0699(.A(new_n706), .B1(new_n233), .B2(new_n521), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n245), .A2(new_n696), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n754), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n538), .A2(new_n630), .ZN(new_n903));
  MUX2_X1   g0703(.A(new_n614), .B(new_n679), .S(new_n903), .Z(new_n904));
  OAI221_X1 g0704(.A(new_n276), .B1(new_n716), .B2(new_n359), .C1(new_n257), .C2(new_n758), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n742), .A2(G77), .B1(new_n745), .B2(G137), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n201), .B2(new_n711), .ZN(new_n907));
  OAI22_X1  g0707(.A1(new_n733), .A2(new_n761), .B1(new_n734), .B2(new_n202), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n726), .A2(new_n411), .ZN(new_n909));
  OR4_X1    g0709(.A1(new_n905), .A2(new_n907), .A3(new_n908), .A4(new_n909), .ZN(new_n910));
  AOI22_X1  g0710(.A1(new_n747), .A2(G107), .B1(G294), .B2(new_n721), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n744), .A2(G116), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT46), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n911), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n740), .A2(G283), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n276), .B1(new_n742), .B2(G97), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n912), .A2(new_n913), .B1(new_n732), .B2(G311), .ZN(new_n917));
  XOR2_X1   g0717(.A(KEYINPUT108), .B(G317), .Z(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n745), .A2(new_n919), .B1(new_n736), .B2(G303), .ZN(new_n920));
  NAND4_X1  g0720(.A1(new_n915), .A2(new_n916), .A3(new_n917), .A4(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n910), .B1(new_n914), .B2(new_n921), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n922), .B(KEYINPUT110), .ZN(new_n923));
  XNOR2_X1  g0723(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n923), .B(new_n924), .ZN(new_n925));
  OAI221_X1 g0725(.A(new_n902), .B1(new_n702), .B2(new_n904), .C1(new_n925), .C2(new_n757), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n557), .A2(new_n627), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n682), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n617), .A2(new_n627), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n631), .A2(new_n930), .ZN(new_n931));
  XOR2_X1   g0731(.A(new_n931), .B(KEYINPUT45), .Z(new_n932));
  NOR2_X1   g0732(.A1(new_n631), .A2(new_n930), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT44), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n633), .A2(new_n638), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n935), .B(new_n936), .ZN(new_n937));
  MUX2_X1   g0737(.A(new_n633), .B(new_n496), .S(new_n628), .Z(new_n938));
  XOR2_X1   g0738(.A(new_n938), .B(new_n638), .Z(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n688), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n688), .B1(new_n937), .B2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n641), .B(KEYINPUT41), .Z(new_n943));
  OAI21_X1  g0743(.A(KEYINPUT107), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT107), .ZN(new_n945));
  INV_X1    g0745(.A(new_n943), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n941), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n693), .B1(new_n944), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n936), .A2(new_n930), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT106), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n904), .A2(KEYINPUT43), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n950), .B(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n930), .A2(new_n496), .A3(new_n628), .ZN(new_n953));
  OR2_X1    g0753(.A1(new_n953), .A2(KEYINPUT42), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n571), .B1(new_n928), .B2(new_n486), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n953), .A2(KEYINPUT42), .B1(new_n630), .B2(new_n955), .ZN(new_n956));
  AOI22_X1  g0756(.A1(new_n954), .A2(new_n956), .B1(KEYINPUT43), .B2(new_n904), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n952), .B(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n926), .B1(new_n948), .B2(new_n958), .ZN(G387));
  INV_X1    g0759(.A(new_n699), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n960), .A2(new_n643), .B1(G107), .B2(new_n234), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n242), .A2(new_n451), .ZN(new_n962));
  INV_X1    g0762(.A(new_n643), .ZN(new_n963));
  AOI211_X1 g0763(.A(G45), .B(new_n963), .C1(G68), .C2(G77), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n291), .A2(G50), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT50), .ZN(new_n966));
  AOI211_X1 g0766(.A(new_n233), .B(new_n276), .C1(new_n964), .C2(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n961), .B1(new_n962), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n744), .A2(G77), .ZN(new_n969));
  OAI221_X1 g0769(.A(new_n969), .B1(new_n411), .B2(new_n716), .C1(new_n359), .C2(new_n729), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n734), .A2(new_n430), .ZN(new_n971));
  AOI211_X1 g0771(.A(new_n268), .B(new_n971), .C1(G97), .C2(new_n742), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n972), .B1(new_n257), .B2(new_n733), .C1(new_n291), .C2(new_n758), .ZN(new_n973));
  AOI211_X1 g0773(.A(new_n970), .B(new_n973), .C1(G68), .C2(new_n740), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n919), .A2(new_n736), .B1(G311), .B2(new_n721), .ZN(new_n975));
  INV_X1    g0775(.A(G322), .ZN(new_n976));
  OAI221_X1 g0776(.A(new_n975), .B1(new_n976), .B2(new_n733), .C1(new_n582), .C2(new_n726), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT48), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n977), .A2(new_n978), .ZN(new_n980));
  AOI22_X1  g0780(.A1(new_n744), .A2(G294), .B1(new_n747), .B2(G283), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n979), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT49), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n276), .B1(new_n745), .B2(G326), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n470), .B2(new_n718), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n982), .A2(new_n983), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n974), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n694), .B1(new_n706), .B2(new_n968), .C1(new_n989), .C2(new_n757), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n990), .B1(new_n633), .B2(new_n703), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(new_n939), .B2(new_n693), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n940), .A2(new_n641), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n939), .A2(new_n688), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n992), .B1(new_n993), .B2(new_n994), .ZN(G393));
  OAI21_X1  g0795(.A(new_n705), .B1(new_n524), .B2(new_n234), .ZN(new_n996));
  AND2_X1   g0796(.A1(new_n252), .A2(new_n696), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n694), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n736), .A2(G311), .B1(G317), .B2(new_n732), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT52), .ZN(new_n1000));
  INV_X1    g0800(.A(G283), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n711), .A2(new_n1001), .B1(new_n729), .B2(new_n976), .ZN(new_n1002));
  AOI211_X1 g0802(.A(new_n276), .B(new_n1002), .C1(G107), .C2(new_n742), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n747), .A2(G116), .B1(G303), .B2(new_n721), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n1003), .B(new_n1004), .C1(new_n778), .C2(new_n726), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n711), .A2(new_n202), .B1(new_n729), .B2(new_n761), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n268), .B(new_n1006), .C1(G87), .C2(new_n742), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n734), .A2(new_n367), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(new_n721), .B2(G50), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n1007), .B(new_n1009), .C1(new_n291), .C2(new_n726), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n736), .A2(G159), .B1(G150), .B2(new_n732), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT51), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n1000), .A2(new_n1005), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n998), .B1(new_n1013), .B2(new_n704), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n930), .B2(new_n702), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n937), .B2(new_n692), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  OR2_X1    g0817(.A1(new_n937), .A2(new_n940), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n937), .A2(new_n940), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1018), .A2(new_n641), .A3(new_n1019), .ZN(new_n1020));
  AND2_X1   g0820(.A1(new_n1020), .A2(KEYINPUT111), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1020), .A2(KEYINPUT111), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1017), .B1(new_n1021), .B2(new_n1022), .ZN(G390));
  OAI21_X1  g0823(.A(KEYINPUT104), .B1(new_n843), .B2(new_n853), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n860), .A2(new_n855), .A3(new_n864), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n867), .A2(new_n871), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(new_n811), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1024), .A2(new_n1025), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n790), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n627), .B(new_n1029), .C1(new_n678), .C2(new_n685), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n791), .ZN(new_n1031));
  OAI21_X1  g0831(.A(KEYINPUT112), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n686), .A2(new_n630), .A3(new_n790), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT112), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1033), .A2(new_n1034), .A3(new_n791), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1032), .A2(new_n871), .A3(new_n1035), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n880), .A2(new_n812), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1028), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n871), .ZN(new_n1040));
  NOR4_X1   g0840(.A1(new_n664), .A2(new_n1040), .A3(new_n665), .A4(new_n792), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1041), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1028), .A2(new_n1038), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n449), .A2(new_n666), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n877), .A2(new_n604), .A3(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n871), .B1(new_n666), .B2(new_n793), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n867), .B1(new_n1047), .B2(new_n1041), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1047), .A2(new_n1041), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1046), .B1(new_n1048), .B2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1042), .A2(new_n1044), .A3(new_n1052), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1053), .A2(KEYINPUT113), .A3(new_n641), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1052), .ZN(new_n1055));
  AND3_X1   g0855(.A1(new_n1028), .A2(new_n1038), .A3(new_n1043), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1043), .B1(new_n1028), .B2(new_n1038), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1055), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1054), .A2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(KEYINPUT113), .B1(new_n1053), .B2(new_n641), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1042), .A2(new_n693), .A3(new_n1044), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT116), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1024), .A2(new_n1025), .A3(new_n783), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n769), .B1(new_n470), .B2(new_n716), .C1(new_n778), .C2(new_n729), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(G97), .B2(new_n740), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n733), .A2(new_n1001), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n1008), .B(new_n1066), .C1(G107), .C2(new_n721), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n268), .B1(new_n711), .B2(new_n712), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT115), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1065), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n744), .A2(G150), .ZN(new_n1071));
  INV_X1    g0871(.A(G128), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n1071), .A2(KEYINPUT53), .B1(new_n1072), .B2(new_n733), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n758), .A2(new_n760), .B1(new_n734), .B2(new_n257), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n276), .B1(new_n718), .B2(new_n411), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT114), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(KEYINPUT54), .B(G143), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n740), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(G125), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n716), .A2(new_n766), .B1(new_n729), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(KEYINPUT53), .B2(new_n1071), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n1075), .A2(new_n1077), .A3(new_n1080), .A4(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n757), .B1(new_n1070), .B2(new_n1084), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n754), .B(new_n1085), .C1(new_n291), .C2(new_n784), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1063), .A2(new_n1086), .ZN(new_n1087));
  AND3_X1   g0887(.A1(new_n1061), .A2(new_n1062), .A3(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1062), .B1(new_n1061), .B2(new_n1087), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n1059), .A2(new_n1060), .B1(new_n1088), .B2(new_n1089), .ZN(G378));
  INV_X1    g0890(.A(KEYINPUT119), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n889), .A2(new_n890), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n852), .A2(new_n839), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n886), .B1(new_n1093), .B2(new_n885), .ZN(new_n1094));
  NOR3_X1   g0894(.A1(new_n880), .A2(KEYINPUT105), .A3(new_n883), .ZN(new_n1095));
  OAI211_X1 g0895(.A(G330), .B(new_n1092), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n363), .A2(new_n815), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT55), .Z(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n385), .B(new_n1099), .ZN(new_n1100));
  XOR2_X1   g0900(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n385), .B(new_n1098), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1101), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  AND2_X1   g0905(.A1(new_n1102), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1096), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1102), .A2(new_n1105), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n891), .A2(G330), .A3(new_n1108), .ZN(new_n1109));
  AND4_X1   g0909(.A1(new_n866), .A2(new_n1107), .A3(new_n875), .A4(new_n1109), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n1109), .A2(new_n1107), .B1(new_n866), .B2(new_n875), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n693), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1106), .A2(new_n783), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(G128), .A2(new_n736), .B1(new_n744), .B2(new_n1079), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n766), .B2(new_n758), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n747), .A2(G150), .B1(G125), .B2(new_n732), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1116), .B(new_n1117), .C1(new_n760), .C2(new_n726), .ZN(new_n1118));
  OR2_X1    g0918(.A1(new_n1118), .A2(KEYINPUT59), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(KEYINPUT59), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n742), .A2(G159), .ZN(new_n1121));
  AOI211_X1 g0921(.A(G33), .B(G41), .C1(new_n745), .C2(G124), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .A4(new_n1122), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n718), .A2(new_n201), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n276), .A2(G41), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n1124), .B(new_n1126), .C1(G283), .C2(new_n745), .ZN(new_n1127));
  OAI221_X1 g0927(.A(new_n969), .B1(new_n202), .B2(new_n734), .C1(new_n436), .C2(new_n716), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(G116), .B2(new_n732), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n740), .A2(new_n521), .B1(G97), .B2(new_n721), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT117), .ZN(new_n1131));
  AND2_X1   g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1127), .B(new_n1129), .C1(new_n1132), .C2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT58), .ZN(new_n1135));
  OR2_X1    g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1126), .B(new_n411), .C1(G33), .C2(G41), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1123), .A2(new_n1136), .A3(new_n1137), .A4(new_n1138), .ZN(new_n1139));
  AND2_X1   g0939(.A1(new_n1139), .A2(new_n704), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n754), .B(new_n1140), .C1(new_n411), .C2(new_n784), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1113), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1091), .B1(new_n1112), .B2(new_n1142), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1096), .A2(new_n1106), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1108), .B1(new_n891), .B2(G330), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n811), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n1144), .A2(new_n1145), .B1(new_n1146), .B2(new_n874), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1107), .A2(new_n866), .A3(new_n875), .A4(new_n1109), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n692), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1142), .ZN(new_n1150));
  NOR3_X1   g0950(.A1(new_n1149), .A2(KEYINPUT119), .A3(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1143), .A2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1051), .A2(new_n1048), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1046), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(KEYINPUT57), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1156));
  OAI21_X1  g0956(.A(KEYINPUT120), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1046), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1053), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT120), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1159), .A2(new_n1160), .A3(KEYINPUT57), .A4(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1157), .A2(new_n1162), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n1053), .A2(new_n1158), .B1(new_n1148), .B2(new_n1147), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n641), .B1(new_n1164), .B2(KEYINPUT57), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1152), .B1(new_n1163), .B2(new_n1165), .ZN(G375));
  INV_X1    g0966(.A(new_n1154), .ZN(new_n1167));
  OAI21_X1  g0967(.A(KEYINPUT121), .B1(new_n1167), .B2(new_n692), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT121), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1154), .A2(new_n1169), .A3(new_n693), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1040), .A2(new_n783), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n754), .B1(new_n784), .B2(new_n202), .ZN(new_n1172));
  XOR2_X1   g0972(.A(new_n1172), .B(KEYINPUT122), .Z(new_n1173));
  AOI211_X1 g0973(.A(new_n268), .B(new_n1124), .C1(new_n721), .C2(new_n1079), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n740), .A2(G150), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n747), .A2(G50), .B1(G132), .B2(new_n732), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n711), .A2(new_n257), .B1(new_n729), .B2(new_n1072), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(G137), .B2(new_n736), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .A4(new_n1178), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n276), .B(new_n971), .C1(G77), .C2(new_n742), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n740), .A2(G107), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(G116), .A2(new_n721), .B1(new_n732), .B2(G294), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n711), .A2(new_n524), .B1(new_n729), .B2(new_n582), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(G283), .B2(new_n736), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1180), .A2(new_n1181), .A3(new_n1182), .A4(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n757), .B1(new_n1179), .B2(new_n1185), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1173), .A2(new_n1186), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n1168), .A2(new_n1170), .B1(new_n1171), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1167), .A2(new_n1046), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1189), .A2(new_n946), .A3(new_n1055), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1188), .A2(new_n1190), .ZN(G381));
  OR3_X1    g0991(.A1(G384), .A2(G393), .A3(G396), .ZN(new_n1192));
  NOR4_X1   g0992(.A1(G387), .A2(G390), .A3(G381), .A4(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(G375), .ZN(new_n1194));
  INV_X1    g0994(.A(G378), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .ZN(G407));
  NAND2_X1  g0996(.A1(new_n626), .A2(G213), .ZN(new_n1197));
  XOR2_X1   g0997(.A(new_n1197), .B(KEYINPUT123), .Z(new_n1198));
  NAND3_X1  g0998(.A1(new_n1194), .A2(new_n1195), .A3(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(G407), .A2(new_n1199), .A3(G213), .ZN(G409));
  INV_X1    g1000(.A(KEYINPUT60), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1189), .B1(new_n1201), .B2(new_n1052), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1167), .A2(KEYINPUT60), .A3(new_n1046), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1202), .A2(new_n641), .A3(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(new_n1188), .ZN(new_n1205));
  INV_X1    g1005(.A(G384), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1204), .A2(G384), .A3(new_n1188), .ZN(new_n1208));
  AND2_X1   g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(G2897), .B2(new_n1198), .ZN(new_n1210));
  AND3_X1   g1010(.A1(new_n626), .A2(G213), .A3(G2897), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1210), .B1(new_n1209), .B2(new_n1211), .ZN(new_n1212));
  OAI211_X1 g1012(.A(G378), .B(new_n1152), .C1(new_n1163), .C2(new_n1165), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1164), .A2(new_n946), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1214), .A2(new_n1112), .A3(new_n1142), .ZN(new_n1215));
  OR2_X1    g1015(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1060), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1217), .A2(new_n1058), .A3(new_n1054), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1215), .A2(new_n1216), .A3(new_n1218), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n1213), .A2(new_n1219), .B1(G213), .B2(new_n626), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1212), .A2(new_n1220), .ZN(new_n1221));
  OR2_X1    g1021(.A1(new_n948), .A2(new_n958), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1222), .A2(G390), .A3(new_n926), .ZN(new_n1223));
  INV_X1    g1023(.A(G390), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(G387), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1223), .A2(new_n1225), .ZN(new_n1226));
  XOR2_X1   g1026(.A(G393), .B(G396), .Z(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1226), .A2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1223), .A2(new_n1227), .A3(new_n1225), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  NOR3_X1   g1031(.A1(new_n1221), .A2(KEYINPUT61), .A3(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1198), .B1(new_n1213), .B2(new_n1219), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1233), .A2(KEYINPUT63), .A3(new_n1209), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1213), .A2(new_n1219), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1235), .A2(new_n1197), .A3(new_n1209), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT124), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1220), .A2(KEYINPUT124), .A3(new_n1209), .ZN(new_n1239));
  AOI21_X1  g1039(.A(KEYINPUT63), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT125), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  AOI211_X1 g1042(.A(KEYINPUT125), .B(KEYINPUT63), .C1(new_n1238), .C2(new_n1239), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1232), .B(new_n1234), .C1(new_n1242), .C2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT61), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1245), .B1(new_n1212), .B2(new_n1233), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1198), .ZN(new_n1247));
  AND3_X1   g1047(.A1(new_n1207), .A2(new_n1208), .A3(KEYINPUT62), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1235), .A2(new_n1247), .A3(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT127), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1233), .A2(KEYINPUT127), .A3(new_n1248), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(KEYINPUT62), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1253), .B1(new_n1254), .B2(KEYINPUT126), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT62), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1257));
  AOI21_X1  g1057(.A(KEYINPUT124), .B1(new_n1220), .B2(new_n1209), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1256), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT126), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1246), .B1(new_n1255), .B2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1231), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1244), .B1(new_n1262), .B2(new_n1263), .ZN(G405));
  NOR2_X1   g1064(.A1(new_n1194), .A2(G378), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1213), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1267), .B(new_n1209), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(new_n1268), .B(new_n1263), .ZN(G402));
endmodule


