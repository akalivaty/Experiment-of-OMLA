//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 1 0 0 1 1 1 1 1 1 0 1 0 1 0 1 0 0 1 0 0 0 1 0 1 0 1 0 0 0 1 1 1 1 1 1 1 1 1 1 1 0 1 1 1 1 1 0 1 1 0 1 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:55 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n784, new_n785, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028;
  INV_X1    g000(.A(KEYINPUT23), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(G128), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G119), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n187), .A2(G128), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G119), .ZN(new_n191));
  OAI211_X1 g005(.A(new_n189), .B(new_n190), .C1(new_n191), .C2(new_n188), .ZN(new_n192));
  XOR2_X1   g006(.A(KEYINPUT72), .B(G110), .Z(new_n193));
  INV_X1    g007(.A(G119), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(G128), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(KEYINPUT64), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT64), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G119), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n195), .B1(new_n199), .B2(G128), .ZN(new_n200));
  XOR2_X1   g014(.A(KEYINPUT24), .B(G110), .Z(new_n201));
  OAI22_X1  g015(.A1(new_n192), .A2(new_n193), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G140), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G125), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(KEYINPUT16), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G125), .ZN(new_n207));
  AND3_X1   g021(.A1(new_n207), .A2(KEYINPUT71), .A3(G140), .ZN(new_n208));
  XNOR2_X1  g022(.A(G125), .B(G140), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT71), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT16), .ZN(new_n212));
  OAI211_X1 g026(.A(G146), .B(new_n206), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G146), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n209), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n202), .A2(new_n213), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(KEYINPUT73), .ZN(new_n217));
  INV_X1    g031(.A(new_n215), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n207), .A2(G140), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n219), .A2(new_n204), .A3(new_n210), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n207), .A2(KEYINPUT71), .A3(G140), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n205), .B1(new_n222), .B2(KEYINPUT16), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n218), .B1(new_n223), .B2(G146), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT73), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n224), .A2(new_n225), .A3(new_n202), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n217), .A2(new_n226), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n212), .B1(new_n220), .B2(new_n221), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n214), .B1(new_n228), .B2(new_n205), .ZN(new_n229));
  AOI22_X1  g043(.A1(new_n229), .A2(new_n213), .B1(G110), .B2(new_n192), .ZN(new_n230));
  AND3_X1   g044(.A1(new_n200), .A2(KEYINPUT70), .A3(new_n201), .ZN(new_n231));
  AOI21_X1  g045(.A(KEYINPUT70), .B1(new_n200), .B2(new_n201), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n230), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G953), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n235), .A2(G221), .A3(G234), .ZN(new_n236));
  XNOR2_X1  g050(.A(new_n236), .B(KEYINPUT22), .ZN(new_n237));
  XNOR2_X1  g051(.A(new_n237), .B(G137), .ZN(new_n238));
  AND3_X1   g052(.A1(new_n227), .A2(new_n234), .A3(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n238), .B1(new_n227), .B2(new_n234), .ZN(new_n240));
  OAI21_X1  g054(.A(KEYINPUT75), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G217), .ZN(new_n242));
  INV_X1    g056(.A(G902), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n242), .B1(G234), .B2(new_n243), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n244), .A2(G902), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n225), .B1(new_n224), .B2(new_n202), .ZN(new_n246));
  AND4_X1   g060(.A1(new_n225), .A2(new_n202), .A3(new_n213), .A4(new_n215), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n234), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n238), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT75), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n227), .A2(new_n234), .A3(new_n238), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n250), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n241), .A2(new_n245), .A3(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT76), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n241), .A2(KEYINPUT76), .A3(new_n253), .A4(new_n245), .ZN(new_n257));
  AND2_X1   g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n250), .A2(new_n243), .A3(new_n252), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT74), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT25), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  AND2_X1   g076(.A1(new_n259), .A2(new_n261), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n250), .A2(KEYINPUT25), .A3(new_n243), .A4(new_n252), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(KEYINPUT74), .ZN(new_n265));
  OAI211_X1 g079(.A(new_n262), .B(new_n244), .C1(new_n263), .C2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n258), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT11), .ZN(new_n268));
  INV_X1    g082(.A(G134), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n268), .B1(new_n269), .B2(G137), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(G137), .ZN(new_n271));
  INV_X1    g085(.A(G137), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n272), .A2(KEYINPUT11), .A3(G134), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n270), .A2(new_n271), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(G131), .ZN(new_n275));
  INV_X1    g089(.A(G131), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n270), .A2(new_n273), .A3(new_n276), .A4(new_n271), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  XNOR2_X1  g093(.A(G143), .B(G146), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n280), .A2(KEYINPUT0), .A3(G128), .ZN(new_n281));
  XNOR2_X1  g095(.A(KEYINPUT0), .B(G128), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n281), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n279), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G128), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n285), .A2(KEYINPUT1), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n214), .A2(G143), .ZN(new_n287));
  INV_X1    g101(.A(G143), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G146), .ZN(new_n289));
  AND3_X1   g103(.A1(new_n286), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n288), .B(G146), .C1(new_n285), .C2(KEYINPUT1), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n285), .A2(new_n214), .A3(G143), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n271), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n269), .A2(G137), .ZN(new_n296));
  OAI21_X1  g110(.A(G131), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n277), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n294), .A2(new_n298), .ZN(new_n299));
  NOR3_X1   g113(.A1(new_n284), .A2(KEYINPUT30), .A3(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT66), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT65), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n303), .B1(new_n290), .B2(new_n293), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n286), .A2(new_n287), .A3(new_n289), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n305), .A2(KEYINPUT65), .A3(new_n291), .A4(new_n292), .ZN(new_n306));
  AOI211_X1 g120(.A(new_n302), .B(new_n298), .C1(new_n304), .C2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n304), .A2(new_n306), .ZN(new_n308));
  INV_X1    g122(.A(new_n298), .ZN(new_n309));
  AOI21_X1  g123(.A(KEYINPUT66), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NOR3_X1   g124(.A1(new_n307), .A2(new_n310), .A3(new_n284), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT30), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n301), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n199), .A2(G116), .ZN(new_n314));
  INV_X1    g128(.A(G116), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G119), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  XOR2_X1   g131(.A(KEYINPUT2), .B(G113), .Z(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n314), .A2(new_n316), .A3(new_n318), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n313), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT31), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n307), .A2(new_n310), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n284), .A2(new_n322), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G237), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(KEYINPUT67), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT67), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G237), .ZN(new_n331));
  AOI21_X1  g145(.A(G953), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G210), .ZN(new_n333));
  XOR2_X1   g147(.A(KEYINPUT68), .B(KEYINPUT27), .Z(new_n334));
  XNOR2_X1  g148(.A(new_n333), .B(new_n334), .ZN(new_n335));
  XNOR2_X1  g149(.A(KEYINPUT26), .B(G101), .ZN(new_n336));
  XOR2_X1   g150(.A(new_n335), .B(new_n336), .Z(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n323), .A2(new_n324), .A3(new_n327), .A4(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n308), .A2(new_n309), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(new_n302), .ZN(new_n341));
  INV_X1    g155(.A(new_n283), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n278), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n308), .A2(KEYINPUT66), .A3(new_n309), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n341), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n300), .B1(new_n345), .B2(KEYINPUT30), .ZN(new_n346));
  AND2_X1   g160(.A1(new_n320), .A2(new_n321), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n327), .B(new_n338), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(KEYINPUT31), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT28), .ZN(new_n350));
  INV_X1    g164(.A(new_n299), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(new_n343), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(new_n322), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n350), .B1(new_n327), .B2(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(KEYINPUT28), .B1(new_n326), .B2(new_n340), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n337), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n339), .A2(new_n349), .A3(new_n356), .ZN(new_n357));
  NOR2_X1   g171(.A1(G472), .A2(G902), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n357), .A2(KEYINPUT32), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(KEYINPUT32), .B1(new_n357), .B2(new_n358), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT29), .ZN(new_n362));
  INV_X1    g176(.A(new_n355), .ZN(new_n363));
  AOI22_X1  g177(.A1(new_n325), .A2(new_n326), .B1(new_n352), .B2(new_n322), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n363), .B(new_n338), .C1(new_n364), .C2(new_n350), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n347), .A2(new_n343), .ZN(new_n366));
  NOR3_X1   g180(.A1(new_n366), .A2(new_n307), .A3(new_n310), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n367), .B1(new_n313), .B2(new_n322), .ZN(new_n368));
  OAI211_X1 g182(.A(new_n362), .B(new_n365), .C1(new_n368), .C2(new_n338), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(KEYINPUT69), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n327), .B1(new_n346), .B2(new_n347), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n337), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT69), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n372), .A2(new_n373), .A3(new_n362), .A4(new_n365), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n367), .B1(new_n322), .B2(new_n345), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n363), .B1(new_n375), .B2(new_n350), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n338), .A2(KEYINPUT29), .ZN(new_n377));
  OR2_X1    g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n370), .A2(new_n374), .A3(new_n243), .A4(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G472), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n267), .B1(new_n361), .B2(new_n380), .ZN(new_n381));
  XOR2_X1   g195(.A(KEYINPUT9), .B(G234), .Z(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  OAI21_X1  g197(.A(G221), .B1(new_n383), .B2(G902), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  XNOR2_X1  g199(.A(G110), .B(G140), .ZN(new_n386));
  AND2_X1   g200(.A1(new_n235), .A2(G227), .ZN(new_n387));
  XOR2_X1   g201(.A(new_n386), .B(new_n387), .Z(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n294), .ZN(new_n390));
  INV_X1    g204(.A(G101), .ZN(new_n391));
  INV_X1    g205(.A(G107), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G104), .ZN(new_n393));
  INV_X1    g207(.A(G104), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(G107), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n391), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT81), .ZN(new_n397));
  OR2_X1    g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n392), .A2(G104), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n394), .A2(G107), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT77), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n401), .A2(KEYINPUT3), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n399), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT3), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT77), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n404), .A2(KEYINPUT77), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n405), .B1(new_n406), .B2(new_n393), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n403), .A2(new_n391), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n396), .A2(new_n397), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n390), .A2(new_n398), .A3(new_n408), .A4(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT10), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n398), .A2(new_n408), .A3(new_n409), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n415), .A2(KEYINPUT10), .A3(new_n308), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n391), .B1(new_n403), .B2(new_n407), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n408), .B1(new_n418), .B2(KEYINPUT78), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n401), .A2(KEYINPUT3), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n402), .B1(new_n400), .B2(new_n420), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n404), .A2(new_n392), .A3(KEYINPUT77), .A4(G104), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n395), .ZN(new_n423));
  OAI211_X1 g237(.A(KEYINPUT78), .B(G101), .C1(new_n421), .C2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT4), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n342), .B1(new_n419), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT4), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n427), .B(G101), .C1(new_n421), .C2(new_n423), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT79), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n403), .A2(new_n407), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n431), .A2(KEYINPUT79), .A3(new_n427), .A4(G101), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(KEYINPUT80), .B1(new_n426), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(G101), .B1(new_n421), .B2(new_n423), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT78), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n437), .A2(KEYINPUT4), .A3(new_n408), .A4(new_n424), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n430), .A2(new_n432), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT80), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n438), .A2(new_n439), .A3(new_n440), .A4(new_n342), .ZN(new_n441));
  AOI211_X1 g255(.A(new_n413), .B(new_n417), .C1(new_n434), .C2(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n389), .B1(new_n442), .B2(new_n279), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n434), .A2(new_n441), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n444), .A2(new_n412), .A3(new_n416), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n278), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n444), .A2(new_n279), .A3(new_n412), .A4(new_n416), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n414), .A2(new_n294), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n410), .ZN(new_n449));
  AOI21_X1  g263(.A(KEYINPUT12), .B1(new_n449), .B2(new_n278), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n449), .A2(KEYINPUT12), .A3(new_n278), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n447), .A2(new_n453), .ZN(new_n454));
  AOI22_X1  g268(.A1(new_n443), .A2(new_n446), .B1(new_n454), .B2(new_n389), .ZN(new_n455));
  OAI21_X1  g269(.A(G469), .B1(new_n455), .B2(G902), .ZN(new_n456));
  XNOR2_X1  g270(.A(KEYINPUT82), .B(G469), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n388), .B1(new_n446), .B2(new_n447), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT12), .ZN(new_n460));
  AOI211_X1 g274(.A(new_n460), .B(new_n279), .C1(new_n448), .C2(new_n410), .ZN(new_n461));
  OAI21_X1  g275(.A(KEYINPUT83), .B1(new_n450), .B2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT83), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n451), .A2(new_n463), .A3(new_n452), .ZN(new_n464));
  AND4_X1   g278(.A1(new_n447), .A2(new_n388), .A3(new_n462), .A4(new_n464), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n243), .B(new_n458), .C1(new_n459), .C2(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n385), .B1(new_n456), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(G475), .A2(G902), .ZN(new_n468));
  XNOR2_X1  g282(.A(G113), .B(G122), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n469), .B(new_n394), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT18), .ZN(new_n471));
  NOR3_X1   g285(.A1(new_n471), .A2(new_n276), .A3(KEYINPUT88), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n329), .A2(new_n331), .ZN(new_n473));
  AND4_X1   g287(.A1(G143), .A2(new_n473), .A3(G214), .A4(new_n235), .ZN(new_n474));
  AOI21_X1  g288(.A(G143), .B1(new_n332), .B2(G214), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n472), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n215), .B1(new_n222), .B2(new_n214), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n473), .A2(G214), .A3(new_n235), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(new_n288), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n332), .A2(G143), .A3(G214), .ZN(new_n480));
  INV_X1    g294(.A(new_n472), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n476), .A2(new_n477), .A3(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(G131), .B1(new_n474), .B2(new_n475), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT17), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n479), .A2(new_n276), .A3(new_n480), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  OAI211_X1 g301(.A(KEYINPUT17), .B(G131), .C1(new_n474), .C2(new_n475), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n488), .A2(new_n213), .A3(new_n229), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n470), .B(new_n483), .C1(new_n487), .C2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n220), .A2(KEYINPUT19), .A3(new_n221), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT19), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n209), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n492), .A2(new_n214), .A3(new_n494), .ZN(new_n495));
  AOI22_X1  g309(.A1(new_n484), .A2(new_n486), .B1(KEYINPUT89), .B2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT89), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n492), .A2(new_n497), .A3(new_n214), .A4(new_n494), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n213), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n470), .B1(new_n500), .B2(new_n483), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n468), .B1(new_n491), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT90), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT20), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n506), .A2(new_n213), .A3(new_n229), .A4(new_n488), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n470), .B1(new_n507), .B2(new_n483), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n243), .B1(new_n491), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(G475), .ZN(new_n510));
  OAI211_X1 g324(.A(KEYINPUT90), .B(new_n468), .C1(new_n491), .C2(new_n501), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(KEYINPUT20), .ZN(new_n512));
  AND2_X1   g326(.A1(new_n476), .A2(new_n482), .ZN(new_n513));
  AOI22_X1  g327(.A1(new_n499), .A2(new_n496), .B1(new_n513), .B2(new_n477), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n490), .B1(new_n514), .B2(new_n470), .ZN(new_n515));
  AOI21_X1  g329(.A(KEYINPUT90), .B1(new_n515), .B2(new_n468), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n505), .B(new_n510), .C1(new_n512), .C2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(KEYINPUT91), .ZN(new_n518));
  OAI21_X1  g332(.A(KEYINPUT93), .B1(new_n285), .B2(G143), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT93), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n520), .A2(new_n288), .A3(G128), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n285), .A2(G143), .ZN(new_n523));
  AND3_X1   g337(.A1(new_n522), .A2(new_n269), .A3(new_n523), .ZN(new_n524));
  XNOR2_X1  g338(.A(KEYINPUT94), .B(KEYINPUT13), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT95), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OR2_X1    g342(.A1(new_n522), .A2(new_n525), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n522), .A2(KEYINPUT95), .A3(new_n525), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n528), .A2(new_n529), .A3(new_n523), .A4(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n524), .B1(new_n531), .B2(G134), .ZN(new_n532));
  XNOR2_X1  g346(.A(G116), .B(G122), .ZN(new_n533));
  XNOR2_X1  g347(.A(KEYINPUT92), .B(G107), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n533), .B(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  OR2_X1    g350(.A1(new_n315), .A2(G122), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n392), .B1(new_n537), .B2(KEYINPUT14), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n538), .B(new_n533), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n269), .B1(new_n522), .B2(new_n523), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n539), .B1(new_n524), .B2(new_n540), .ZN(new_n541));
  NOR3_X1   g355(.A1(new_n383), .A2(new_n242), .A3(G953), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n536), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n542), .B1(new_n536), .B2(new_n541), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n243), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(G478), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n547), .A2(KEYINPUT15), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n536), .A2(new_n541), .ZN(new_n550));
  INV_X1    g364(.A(new_n542), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n543), .ZN(new_n553));
  INV_X1    g367(.A(new_n548), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n553), .A2(new_n243), .A3(new_n554), .ZN(new_n555));
  AND2_X1   g369(.A1(new_n549), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n502), .A2(new_n503), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n557), .A2(KEYINPUT20), .A3(new_n511), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT91), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n558), .A2(new_n559), .A3(new_n505), .A4(new_n510), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n518), .A2(new_n556), .A3(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(G952), .ZN(new_n562));
  AOI211_X1 g376(.A(G953), .B(new_n562), .C1(G234), .C2(G237), .ZN(new_n563));
  XNOR2_X1  g377(.A(KEYINPUT21), .B(G898), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n564), .B(KEYINPUT96), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  AOI211_X1 g380(.A(new_n243), .B(new_n235), .C1(G234), .C2(G237), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n563), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(G214), .B1(G237), .B2(G902), .ZN(new_n570));
  AOI22_X1  g384(.A1(new_n430), .A2(new_n432), .B1(new_n320), .B2(new_n321), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n438), .ZN(new_n572));
  OAI211_X1 g386(.A(KEYINPUT5), .B(new_n316), .C1(new_n191), .C2(new_n315), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT5), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n199), .A2(new_n574), .A3(G116), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n573), .A2(G113), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n321), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n577), .A2(new_n414), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n572), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT85), .ZN(new_n581));
  XNOR2_X1  g395(.A(G110), .B(G122), .ZN(new_n582));
  XOR2_X1   g396(.A(new_n582), .B(KEYINPUT84), .Z(new_n583));
  NAND3_X1  g397(.A1(new_n580), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n578), .B1(new_n438), .B2(new_n571), .ZN(new_n585));
  INV_X1    g399(.A(new_n583), .ZN(new_n586));
  OAI21_X1  g400(.A(KEYINPUT85), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT6), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n588), .B1(new_n585), .B2(new_n582), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n584), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(KEYINPUT86), .B(KEYINPUT6), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n580), .A2(new_n583), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n294), .A2(new_n207), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n593), .B1(new_n342), .B2(new_n207), .ZN(new_n594));
  INV_X1    g408(.A(G224), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n595), .A2(G953), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(KEYINPUT87), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n594), .B(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n590), .A2(new_n592), .A3(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(G210), .B1(G237), .B2(G902), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n577), .B(new_n414), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n582), .B(KEYINPUT8), .ZN(new_n602));
  AOI22_X1  g416(.A1(new_n585), .A2(new_n582), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(KEYINPUT7), .B1(new_n595), .B2(G953), .ZN(new_n604));
  XOR2_X1   g418(.A(new_n594), .B(new_n604), .Z(new_n605));
  AOI21_X1  g419(.A(G902), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  AND3_X1   g420(.A1(new_n599), .A2(new_n600), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n600), .B1(new_n599), .B2(new_n606), .ZN(new_n608));
  OAI211_X1 g422(.A(new_n569), .B(new_n570), .C1(new_n607), .C2(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n561), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n381), .A2(new_n467), .A3(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(G101), .ZN(G3));
  INV_X1    g426(.A(new_n266), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n256), .A2(new_n257), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n356), .B1(new_n348), .B2(KEYINPUT31), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n324), .B1(new_n368), .B2(new_n338), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n243), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  AOI22_X1  g432(.A1(new_n618), .A2(G472), .B1(new_n358), .B2(new_n357), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n467), .A2(new_n615), .A3(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n518), .A2(new_n560), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT33), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n553), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n552), .A2(KEYINPUT33), .A3(new_n543), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n624), .A2(G478), .A3(new_n243), .A4(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n546), .A2(new_n547), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n622), .A2(new_n628), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n629), .A2(KEYINPUT97), .A3(new_n609), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT97), .ZN(new_n631));
  INV_X1    g445(.A(new_n609), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n626), .A2(new_n627), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n633), .B1(new_n518), .B2(new_n560), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n631), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n621), .B1(new_n630), .B2(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(new_n394), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(KEYINPUT98), .ZN(new_n638));
  XOR2_X1   g452(.A(new_n638), .B(KEYINPUT34), .Z(G6));
  NAND2_X1  g453(.A1(new_n549), .A2(new_n555), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n640), .A2(new_n558), .A3(new_n505), .A4(new_n510), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n609), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n621), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT35), .B(G107), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G9));
  NOR2_X1   g459(.A1(new_n249), .A2(KEYINPUT36), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n248), .B(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n245), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n266), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n610), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n467), .A2(new_n619), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT37), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G110), .ZN(G12));
  INV_X1    g468(.A(KEYINPUT99), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n517), .A2(new_n556), .ZN(new_n656));
  INV_X1    g470(.A(G900), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n567), .A2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n563), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n655), .B1(new_n656), .B2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n660), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n641), .A2(KEYINPUT99), .A3(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n361), .A2(new_n380), .ZN(new_n665));
  INV_X1    g479(.A(new_n570), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n599), .A2(new_n606), .ZN(new_n667));
  INV_X1    g481(.A(new_n600), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n599), .A2(new_n600), .A3(new_n606), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n666), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  AND2_X1   g485(.A1(new_n671), .A2(new_n649), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n664), .A2(new_n665), .A3(new_n467), .A4(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G128), .ZN(G30));
  NAND2_X1  g488(.A1(new_n456), .A2(new_n466), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n384), .ZN(new_n676));
  XOR2_X1   g490(.A(new_n660), .B(KEYINPUT39), .Z(new_n677));
  NOR2_X1   g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT40), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n358), .B1(new_n616), .B2(new_n617), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT32), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n357), .A2(KEYINPUT32), .A3(new_n358), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n368), .A2(new_n337), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n375), .A2(new_n337), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(new_n243), .ZN(new_n686));
  OAI21_X1  g500(.A(G472), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n682), .A2(new_n683), .A3(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT101), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n682), .A2(KEYINPUT101), .A3(new_n683), .A4(new_n687), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n648), .ZN(new_n693));
  INV_X1    g507(.A(new_n244), .ZN(new_n694));
  AND2_X1   g508(.A1(new_n264), .A2(KEYINPUT74), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n259), .A2(new_n261), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n694), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n693), .B1(new_n697), .B2(new_n262), .ZN(new_n698));
  AND4_X1   g512(.A1(new_n640), .A2(new_n622), .A3(new_n570), .A4(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(KEYINPUT102), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n607), .A2(new_n608), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT100), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n669), .A2(new_n670), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(KEYINPUT100), .ZN(new_n705));
  AND3_X1   g519(.A1(new_n703), .A2(new_n705), .A3(KEYINPUT38), .ZN(new_n706));
  AOI21_X1  g520(.A(KEYINPUT38), .B1(new_n703), .B2(new_n705), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n679), .A2(new_n692), .A3(new_n700), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G143), .ZN(G45));
  AOI211_X1 g524(.A(new_n662), .B(new_n633), .C1(new_n518), .C2(new_n560), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n711), .A2(new_n665), .A3(new_n467), .A4(new_n672), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G146), .ZN(G48));
  INV_X1    g527(.A(new_n447), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n417), .B1(new_n434), .B2(new_n441), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n279), .B1(new_n715), .B2(new_n412), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n389), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n447), .A2(new_n388), .A3(new_n462), .A4(new_n464), .ZN(new_n718));
  AOI211_X1 g532(.A(G902), .B(new_n457), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(G469), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n243), .B1(new_n459), .B2(new_n465), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT103), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n720), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(G902), .B1(new_n717), .B2(new_n718), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(KEYINPUT103), .ZN(new_n725));
  AOI211_X1 g539(.A(new_n385), .B(new_n719), .C1(new_n723), .C2(new_n725), .ZN(new_n726));
  OAI211_X1 g540(.A(new_n381), .B(new_n726), .C1(new_n630), .C2(new_n635), .ZN(new_n727));
  XNOR2_X1  g541(.A(KEYINPUT41), .B(G113), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(G15));
  NAND3_X1  g543(.A1(new_n726), .A2(new_n381), .A3(new_n642), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G116), .ZN(G18));
  AOI21_X1  g545(.A(new_n561), .B1(new_n361), .B2(new_n380), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n726), .A2(new_n732), .A3(new_n569), .A4(new_n672), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G119), .ZN(G21));
  OAI21_X1  g548(.A(G469), .B1(new_n724), .B2(KEYINPUT103), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n721), .A2(new_n722), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n384), .B(new_n466), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(new_n348), .ZN(new_n738));
  AOI22_X1  g552(.A1(new_n324), .A2(new_n738), .B1(new_n376), .B2(new_n337), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n349), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n358), .ZN(new_n741));
  INV_X1    g555(.A(G472), .ZN(new_n742));
  AOI211_X1 g556(.A(KEYINPUT104), .B(new_n742), .C1(new_n357), .C2(new_n243), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT104), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n744), .B1(new_n618), .B2(G472), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n741), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g560(.A(KEYINPUT105), .B1(new_n613), .B2(new_n614), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT105), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n258), .A2(new_n748), .A3(new_n266), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  NOR4_X1   g564(.A1(new_n737), .A2(new_n746), .A3(new_n750), .A4(new_n568), .ZN(new_n751));
  INV_X1    g565(.A(new_n622), .ZN(new_n752));
  NOR4_X1   g566(.A1(new_n752), .A2(new_n556), .A3(new_n666), .A4(new_n701), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G122), .ZN(G24));
  AOI211_X1 g569(.A(G472), .B(G902), .C1(new_n739), .C2(new_n349), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n618), .A2(G472), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(KEYINPUT104), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n618), .A2(new_n744), .A3(G472), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n756), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n726), .A2(new_n672), .A3(new_n711), .A4(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(KEYINPUT106), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G125), .ZN(G27));
  INV_X1    g577(.A(KEYINPUT107), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n379), .A2(G472), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n682), .A2(new_n683), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n615), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n607), .A2(new_n608), .A3(new_n666), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n467), .A2(new_n634), .A3(new_n660), .A4(new_n768), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n764), .B1(new_n767), .B2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT42), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n675), .A2(new_n768), .A3(new_n384), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n381), .A2(new_n772), .A3(KEYINPUT107), .A4(new_n711), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n770), .A2(new_n771), .A3(new_n773), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n747), .A2(new_n749), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n665), .ZN(new_n776));
  OR3_X1    g590(.A1(new_n776), .A2(new_n771), .A3(new_n769), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(KEYINPUT108), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT108), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n774), .A2(new_n777), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G131), .ZN(G33));
  AND3_X1   g597(.A1(new_n381), .A2(new_n772), .A3(new_n664), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(KEYINPUT109), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(new_n269), .ZN(G36));
  INV_X1    g600(.A(KEYINPUT45), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n447), .A2(new_n388), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n788), .A2(new_n716), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n388), .B1(new_n447), .B2(new_n453), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n787), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n446), .A2(new_n447), .A3(new_n388), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n454), .A2(new_n389), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n792), .A2(new_n793), .A3(KEYINPUT45), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n791), .A2(G469), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(G469), .A2(G902), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT46), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(KEYINPUT110), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n795), .A2(KEYINPUT46), .A3(new_n796), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT110), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n797), .A2(new_n802), .A3(new_n798), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n800), .A2(new_n466), .A3(new_n801), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(new_n384), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n677), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n518), .A2(new_n560), .A3(new_n628), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT43), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n518), .A2(new_n560), .A3(new_n628), .A4(KEYINPUT43), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n619), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(new_n649), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT44), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n806), .A2(new_n807), .A3(new_n815), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n768), .B1(new_n813), .B2(new_n814), .ZN(new_n817));
  OR2_X1    g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(G137), .ZN(G39));
  INV_X1    g633(.A(KEYINPUT111), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n820), .A2(KEYINPUT47), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n805), .A2(new_n822), .ZN(new_n823));
  NOR4_X1   g637(.A1(new_n665), .A2(new_n629), .A3(new_n615), .A4(new_n662), .ZN(new_n824));
  XNOR2_X1  g638(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n804), .A2(new_n384), .A3(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n823), .A2(new_n768), .A3(new_n824), .A4(new_n827), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(G140), .ZN(G42));
  NAND2_X1  g643(.A1(new_n701), .A2(new_n570), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n737), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n659), .B1(new_n810), .B2(new_n811), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n776), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  XOR2_X1   g649(.A(new_n835), .B(KEYINPUT48), .Z(new_n836));
  NOR3_X1   g650(.A1(new_n737), .A2(new_n267), .A3(new_n830), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n659), .B1(new_n690), .B2(new_n691), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n837), .A2(new_n838), .A3(new_n634), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n746), .A2(new_n750), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n840), .A2(new_n832), .A3(new_n671), .A4(new_n726), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n839), .A2(new_n841), .A3(G952), .A4(new_n235), .ZN(new_n842));
  XOR2_X1   g656(.A(new_n842), .B(KEYINPUT116), .Z(new_n843));
  NAND3_X1  g657(.A1(new_n840), .A2(new_n768), .A3(new_n832), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(KEYINPUT115), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n823), .A2(new_n827), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n719), .B1(new_n723), .B2(new_n725), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(new_n385), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n845), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  AND4_X1   g663(.A1(new_n649), .A2(new_n831), .A3(new_n760), .A4(new_n832), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n837), .A2(new_n838), .A3(new_n752), .A4(new_n633), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT50), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n840), .A2(new_n832), .A3(new_n666), .A4(new_n726), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n853), .B1(new_n854), .B2(new_n708), .ZN(new_n855));
  INV_X1    g669(.A(new_n855), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n854), .A2(new_n708), .A3(new_n853), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n851), .B(new_n852), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(KEYINPUT51), .B1(new_n849), .B2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n852), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n840), .A2(new_n726), .A3(new_n832), .ZN(new_n861));
  INV_X1    g675(.A(new_n708), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n861), .A2(KEYINPUT50), .A3(new_n862), .A4(new_n666), .ZN(new_n863));
  AOI211_X1 g677(.A(new_n850), .B(new_n860), .C1(new_n863), .C2(new_n855), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n804), .A2(new_n384), .A3(new_n826), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n821), .B1(new_n804), .B2(new_n384), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n848), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  XOR2_X1   g681(.A(new_n844), .B(KEYINPUT115), .Z(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT51), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n864), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  AOI211_X1 g685(.A(new_n836), .B(new_n843), .C1(new_n859), .C2(new_n871), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n640), .B(KEYINPUT113), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n830), .A2(new_n873), .A3(new_n517), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n874), .A2(new_n665), .A3(new_n467), .A4(new_n660), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n772), .A2(new_n760), .A3(new_n711), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n784), .B1(new_n877), .B2(new_n649), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT112), .ZN(new_n879));
  AND4_X1   g693(.A1(new_n665), .A2(new_n610), .A3(new_n615), .A4(new_n467), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n632), .A2(new_n634), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n620), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n879), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  OAI211_X1 g697(.A(new_n611), .B(KEYINPUT112), .C1(new_n881), .C2(new_n620), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n727), .A2(new_n730), .A3(new_n733), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n632), .A2(new_n752), .A3(new_n873), .ZN(new_n887));
  OAI22_X1  g701(.A1(new_n650), .A2(new_n651), .B1(new_n887), .B2(new_n620), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n888), .B1(new_n751), .B2(new_n753), .ZN(new_n889));
  AND4_X1   g703(.A1(new_n878), .A2(new_n885), .A3(new_n886), .A4(new_n889), .ZN(new_n890));
  AOI221_X4 g704(.A(new_n385), .B1(new_n669), .B2(new_n670), .C1(new_n456), .C2(new_n466), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n699), .A2(new_n891), .A3(new_n660), .A4(new_n688), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n761), .A2(new_n892), .A3(new_n673), .A4(new_n712), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(KEYINPUT52), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n676), .B1(new_n361), .B2(new_n380), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n895), .B(new_n672), .C1(new_n664), .C2(new_n711), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT52), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n896), .A2(new_n897), .A3(new_n761), .A4(new_n892), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n894), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(KEYINPUT114), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT114), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n894), .A2(new_n898), .A3(new_n901), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n890), .A2(new_n782), .A3(new_n900), .A4(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(KEYINPUT53), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT53), .ZN(new_n905));
  INV_X1    g719(.A(new_n899), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n890), .A2(new_n782), .A3(new_n905), .A4(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n904), .A2(KEYINPUT54), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n890), .A2(new_n782), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n900), .A2(new_n902), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n905), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT54), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n905), .B1(new_n774), .B2(new_n777), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n890), .A2(new_n906), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n911), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n872), .A2(new_n908), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n562), .A2(new_n235), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NOR4_X1   g732(.A1(new_n708), .A2(new_n692), .A3(new_n750), .A4(new_n808), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n847), .B(KEYINPUT49), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n919), .A2(new_n384), .A3(new_n570), .A4(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(KEYINPUT117), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT117), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n918), .A2(new_n924), .A3(new_n921), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n923), .A2(new_n925), .ZN(G75));
  AND2_X1   g740(.A1(new_n903), .A2(new_n905), .ZN(new_n927));
  AND3_X1   g741(.A1(new_n890), .A2(new_n906), .A3(new_n913), .ZN(new_n928));
  OAI211_X1 g742(.A(G210), .B(G902), .C1(new_n927), .C2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT56), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n590), .A2(new_n592), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(new_n598), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT55), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n933), .B1(KEYINPUT118), .B2(KEYINPUT56), .ZN(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n929), .A2(new_n930), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n935), .B1(new_n929), .B2(new_n930), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n235), .A2(G952), .ZN(new_n938));
  NOR3_X1   g752(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(G51));
  NAND2_X1  g753(.A1(new_n717), .A2(new_n718), .ZN(new_n940));
  OAI21_X1  g754(.A(KEYINPUT54), .B1(new_n927), .B2(new_n928), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n941), .A2(new_n915), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n796), .B(KEYINPUT57), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n940), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n928), .B1(new_n905), .B2(new_n903), .ZN(new_n945));
  OR3_X1    g759(.A1(new_n945), .A2(new_n243), .A3(new_n795), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n938), .B1(new_n944), .B2(new_n946), .ZN(G54));
  NOR2_X1   g761(.A1(new_n945), .A2(new_n243), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n948), .A2(KEYINPUT58), .A3(G475), .ZN(new_n949));
  INV_X1    g763(.A(new_n515), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(new_n938), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n948), .A2(KEYINPUT58), .A3(G475), .A4(new_n515), .ZN(new_n953));
  AND3_X1   g767(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(G60));
  NAND2_X1  g768(.A1(G478), .A2(G902), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT59), .Z(new_n956));
  AOI21_X1  g770(.A(new_n956), .B1(new_n908), .B2(new_n915), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n624), .A2(new_n625), .ZN(new_n958));
  INV_X1    g772(.A(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n952), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n942), .A2(new_n956), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n960), .B1(new_n961), .B2(new_n959), .ZN(G63));
  NAND2_X1  g776(.A1(new_n241), .A2(new_n253), .ZN(new_n963));
  NAND2_X1  g777(.A1(G217), .A2(G902), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT119), .Z(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT60), .Z(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n963), .B1(new_n945), .B2(new_n967), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n647), .B(new_n966), .C1(new_n927), .C2(new_n928), .ZN(new_n969));
  OR2_X1    g783(.A1(KEYINPUT120), .A2(KEYINPUT61), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n968), .A2(new_n969), .A3(new_n952), .A4(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(KEYINPUT120), .A2(KEYINPUT61), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n971), .B(new_n972), .ZN(G66));
  OAI21_X1  g787(.A(G953), .B1(new_n566), .B2(new_n595), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n885), .A2(new_n886), .A3(new_n889), .ZN(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n974), .B1(new_n976), .B2(G953), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n931), .B1(G898), .B2(new_n235), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(KEYINPUT121), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n977), .B(new_n979), .ZN(G69));
  NAND2_X1  g794(.A1(new_n492), .A2(new_n494), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n313), .B(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  AND2_X1   g797(.A1(new_n896), .A2(new_n761), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n984), .B1(new_n816), .B2(new_n817), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(KEYINPUT124), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT124), .ZN(new_n987));
  OAI211_X1 g801(.A(new_n987), .B(new_n984), .C1(new_n816), .C2(new_n817), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n784), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n806), .A2(new_n807), .A3(new_n753), .A4(new_n834), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n782), .A2(new_n828), .A3(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(G953), .B1(new_n989), .B2(new_n992), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n235), .A2(G900), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n994), .B(KEYINPUT123), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n983), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n818), .A2(new_n828), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n752), .A2(new_n873), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n998), .A2(new_n629), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n999), .A2(new_n678), .A3(new_n381), .A4(new_n768), .ZN(new_n1000));
  AND3_X1   g814(.A1(new_n709), .A2(KEYINPUT62), .A3(new_n984), .ZN(new_n1001));
  AOI21_X1  g815(.A(KEYINPUT62), .B1(new_n709), .B2(new_n984), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n1000), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n235), .B1(new_n997), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1004), .A2(new_n982), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n996), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n235), .B1(G227), .B2(G900), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n1007), .B(KEYINPUT122), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1006), .B(new_n1008), .ZN(G72));
  NAND3_X1  g823(.A1(new_n989), .A2(new_n976), .A3(new_n992), .ZN(new_n1010));
  NAND2_X1  g824(.A1(G472), .A2(G902), .ZN(new_n1011));
  XOR2_X1   g825(.A(new_n1011), .B(KEYINPUT63), .Z(new_n1012));
  XOR2_X1   g826(.A(new_n1012), .B(KEYINPUT125), .Z(new_n1013));
  INV_X1    g827(.A(new_n1013), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1010), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g829(.A(KEYINPUT127), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n1010), .A2(KEYINPUT127), .A3(new_n1014), .ZN(new_n1018));
  NAND4_X1  g832(.A1(new_n1017), .A2(new_n368), .A3(new_n337), .A4(new_n1018), .ZN(new_n1019));
  NOR3_X1   g833(.A1(new_n997), .A2(new_n1003), .A3(new_n975), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n684), .B1(new_n1020), .B2(new_n1013), .ZN(new_n1021));
  INV_X1    g835(.A(KEYINPUT126), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  OAI211_X1 g837(.A(KEYINPUT126), .B(new_n684), .C1(new_n1020), .C2(new_n1013), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n372), .A2(new_n348), .ZN(new_n1026));
  NAND4_X1  g840(.A1(new_n904), .A2(new_n907), .A3(new_n1012), .A4(new_n1026), .ZN(new_n1027));
  AND2_X1   g841(.A1(new_n1027), .A2(new_n952), .ZN(new_n1028));
  AND3_X1   g842(.A1(new_n1019), .A2(new_n1025), .A3(new_n1028), .ZN(G57));
endmodule


