//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 1 0 0 1 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 0 1 1 1 0 1 1 0 1 1 1 1 0 1 0 1 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:57 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1263, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1316, new_n1317,
    new_n1318;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  XOR2_X1   g0009(.A(KEYINPUT64), .B(G238), .Z(new_n210));
  INV_X1    g0010(.A(G68), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G107), .A2(G264), .ZN(new_n216));
  NAND4_X1  g0016(.A1(new_n213), .A2(new_n214), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n209), .B1(new_n212), .B2(new_n217), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT65), .Z(new_n219));
  INV_X1    g0019(.A(KEYINPUT1), .ZN(new_n220));
  OR2_X1    g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n219), .A2(new_n220), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n209), .A2(G13), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT0), .Z(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n226), .A2(new_n207), .ZN(new_n227));
  OAI21_X1  g0027(.A(G50), .B1(G58), .B2(G68), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n225), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  AND3_X1   g0030(.A1(new_n221), .A2(new_n222), .A3(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT2), .B(G226), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT66), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n236), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G50), .B(G68), .Z(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(G13), .ZN(new_n249));
  NOR3_X1   g0049(.A1(new_n249), .A2(new_n207), .A3(G1), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(new_n211), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(KEYINPUT12), .ZN(new_n252));
  NOR2_X1   g0052(.A1(G20), .A2(G33), .ZN(new_n253));
  AOI22_X1  g0053(.A1(new_n253), .A2(G50), .B1(G20), .B2(new_n211), .ZN(new_n254));
  INV_X1    g0054(.A(G77), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n207), .A2(G33), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n254), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(new_n226), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n257), .A2(KEYINPUT11), .A3(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n250), .A2(new_n259), .ZN(new_n261));
  OR3_X1    g0061(.A1(new_n207), .A2(KEYINPUT67), .A3(G1), .ZN(new_n262));
  OAI21_X1  g0062(.A(KEYINPUT67), .B1(new_n207), .B2(G1), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n261), .A2(new_n264), .A3(G68), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n252), .A2(new_n260), .A3(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(KEYINPUT11), .B1(new_n257), .B2(new_n259), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n226), .B1(G33), .B2(G41), .ZN(new_n270));
  INV_X1    g0070(.A(G274), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n272));
  NOR3_X1   g0072(.A1(new_n270), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n272), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n270), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n273), .B1(G238), .B2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT3), .ZN(new_n277));
  INV_X1    g0077(.A(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G1698), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n281), .A2(G226), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(G33), .A2(G97), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n281), .A2(G1698), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n283), .B(new_n284), .C1(new_n285), .C2(new_n233), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT71), .ZN(new_n287));
  AND3_X1   g0087(.A1(new_n286), .A2(new_n287), .A3(new_n270), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n287), .B1(new_n286), .B2(new_n270), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n276), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(KEYINPUT13), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT13), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n292), .B(new_n276), .C1(new_n288), .C2(new_n289), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT14), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n294), .A2(new_n295), .A3(G169), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n291), .A2(G179), .A3(new_n293), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n295), .B1(new_n294), .B2(G169), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n269), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G190), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n268), .B1(new_n294), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G200), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n303), .B1(new_n291), .B2(new_n293), .ZN(new_n304));
  OR2_X1    g0104(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n300), .A2(new_n305), .ZN(new_n306));
  AND2_X1   g0106(.A1(KEYINPUT3), .A2(G33), .ZN(new_n307));
  NOR2_X1   g0107(.A1(KEYINPUT3), .A2(G33), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n309), .A2(G1698), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(G222), .ZN(new_n311));
  INV_X1    g0111(.A(G223), .ZN(new_n312));
  OAI221_X1 g0112(.A(new_n311), .B1(new_n255), .B2(new_n281), .C1(new_n312), .C2(new_n285), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(new_n270), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n273), .B1(G226), .B2(new_n275), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(G200), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n253), .A2(G150), .ZN(new_n318));
  XNOR2_X1  g0118(.A(KEYINPUT8), .B(G58), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n318), .B1(new_n319), .B2(new_n256), .ZN(new_n320));
  NOR2_X1   g0120(.A1(G58), .A2(G68), .ZN(new_n321));
  INV_X1    g0121(.A(G50), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n207), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n259), .B1(new_n320), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n261), .A2(G50), .A3(new_n264), .ZN(new_n325));
  INV_X1    g0125(.A(new_n250), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n324), .B(new_n325), .C1(G50), .C2(new_n326), .ZN(new_n327));
  XNOR2_X1  g0127(.A(new_n327), .B(KEYINPUT9), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n317), .B(new_n328), .C1(new_n301), .C2(new_n316), .ZN(new_n329));
  XNOR2_X1  g0129(.A(new_n329), .B(KEYINPUT10), .ZN(new_n330));
  AND2_X1   g0130(.A1(new_n314), .A2(new_n315), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n327), .B1(new_n331), .B2(G169), .ZN(new_n332));
  OR2_X1    g0132(.A1(new_n332), .A2(KEYINPUT68), .ZN(new_n333));
  INV_X1    g0133(.A(G179), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n332), .A2(KEYINPUT68), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n333), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n330), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n310), .A2(G232), .ZN(new_n339));
  OAI221_X1 g0139(.A(new_n339), .B1(new_n203), .B2(new_n281), .C1(new_n210), .C2(new_n285), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n270), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n273), .B1(G244), .B2(new_n275), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G169), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(KEYINPUT70), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n346), .B1(G179), .B2(new_n343), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n341), .A2(KEYINPUT70), .A3(new_n334), .A4(new_n342), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n261), .A2(G77), .A3(new_n264), .ZN(new_n349));
  XNOR2_X1  g0149(.A(KEYINPUT15), .B(G87), .ZN(new_n350));
  OAI22_X1  g0150(.A1(new_n350), .A2(new_n256), .B1(new_n207), .B2(new_n255), .ZN(new_n351));
  XNOR2_X1  g0151(.A(new_n319), .B(KEYINPUT69), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n351), .B1(new_n352), .B2(new_n253), .ZN(new_n353));
  INV_X1    g0153(.A(new_n259), .ZN(new_n354));
  OAI221_X1 g0154(.A(new_n349), .B1(G77), .B2(new_n326), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n348), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n347), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n355), .B1(new_n343), .B2(G200), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(new_n301), .B2(new_n343), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NOR3_X1   g0161(.A1(new_n306), .A2(new_n338), .A3(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n264), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n363), .A2(new_n319), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n364), .A2(new_n261), .B1(new_n250), .B2(new_n319), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT7), .ZN(new_n367));
  XNOR2_X1  g0167(.A(KEYINPUT72), .B(G33), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n279), .B1(new_n368), .B2(new_n277), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n367), .B1(new_n369), .B2(G20), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n278), .A2(KEYINPUT72), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT72), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(G33), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n308), .B1(new_n374), .B2(KEYINPUT3), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT73), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n367), .A2(G20), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n279), .B(new_n377), .C1(new_n368), .C2(new_n277), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(KEYINPUT73), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n370), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(G68), .ZN(new_n382));
  INV_X1    g0182(.A(G58), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n383), .A2(new_n211), .ZN(new_n384));
  OR2_X1    g0184(.A1(new_n384), .A2(new_n321), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n385), .A2(G20), .B1(G159), .B2(new_n253), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n382), .A2(KEYINPUT16), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n368), .A2(new_n277), .ZN(new_n388));
  NOR3_X1   g0188(.A1(new_n307), .A2(new_n367), .A3(G20), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n279), .A2(new_n207), .A3(new_n280), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n388), .A2(new_n389), .B1(new_n390), .B2(new_n367), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n386), .B1(new_n391), .B2(new_n211), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT16), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n387), .A2(new_n259), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(KEYINPUT74), .ZN(new_n396));
  INV_X1    g0196(.A(new_n386), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n397), .B1(new_n381), .B2(G68), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n354), .B1(new_n398), .B2(KEYINPUT16), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT74), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n399), .A2(new_n400), .A3(new_n394), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n366), .B1(new_n396), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT75), .ZN(new_n403));
  INV_X1    g0203(.A(G41), .ZN(new_n404));
  OAI211_X1 g0204(.A(G1), .B(G13), .C1(new_n278), .C2(new_n404), .ZN(new_n405));
  MUX2_X1   g0205(.A(G223), .B(G226), .S(G1698), .Z(new_n406));
  NAND2_X1  g0206(.A1(new_n369), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(G33), .A2(G87), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n405), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n273), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n275), .A2(G232), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n403), .B1(new_n409), .B2(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n273), .B1(G232), .B2(new_n275), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n369), .A2(new_n406), .B1(G33), .B2(G87), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n414), .B(KEYINPUT75), .C1(new_n405), .C2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n344), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT76), .ZN(new_n419));
  NOR3_X1   g0219(.A1(new_n409), .A2(new_n412), .A3(G179), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n418), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(G169), .B1(new_n413), .B2(new_n416), .ZN(new_n423));
  OAI21_X1  g0223(.A(KEYINPUT76), .B1(new_n423), .B2(new_n420), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(KEYINPUT18), .B1(new_n402), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n417), .A2(new_n303), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n414), .B1(new_n415), .B2(new_n405), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n427), .B1(G190), .B2(new_n428), .ZN(new_n429));
  AND4_X1   g0229(.A1(new_n400), .A2(new_n387), .A3(new_n259), .A4(new_n394), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n400), .B1(new_n399), .B2(new_n394), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n365), .B(new_n429), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT17), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n365), .B1(new_n430), .B2(new_n431), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT18), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n419), .B1(new_n418), .B2(new_n421), .ZN(new_n437));
  NOR3_X1   g0237(.A1(new_n423), .A2(KEYINPUT76), .A3(new_n420), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n435), .A2(new_n436), .A3(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n402), .A2(KEYINPUT17), .A3(new_n429), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n426), .A2(new_n434), .A3(new_n440), .A4(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  AND2_X1   g0243(.A1(new_n362), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(G116), .ZN(new_n446));
  AOI22_X1  g0246(.A1(new_n258), .A2(new_n226), .B1(G20), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(G33), .A2(G283), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n448), .B(new_n207), .C1(G33), .C2(new_n202), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n447), .A2(KEYINPUT20), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT80), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n447), .A2(new_n449), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT20), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT80), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n447), .A2(new_n455), .A3(new_n449), .A4(KEYINPUT20), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n451), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n326), .A2(G116), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n278), .A2(G1), .ZN(new_n459));
  NOR3_X1   g0259(.A1(new_n250), .A2(new_n259), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n458), .B1(new_n460), .B2(G116), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n270), .A2(new_n271), .ZN(new_n463));
  INV_X1    g0263(.A(G45), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n464), .A2(G1), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT77), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT5), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(G41), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n465), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n206), .B(G45), .C1(new_n404), .C2(KEYINPUT5), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(KEYINPUT77), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n404), .A2(KEYINPUT5), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n463), .A2(new_n469), .A3(new_n471), .A4(new_n472), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n472), .B1(new_n470), .B2(KEYINPUT77), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n466), .B1(new_n465), .B2(new_n468), .ZN(new_n475));
  OAI211_X1 g0275(.A(G270), .B(new_n405), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(G303), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n281), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g0278(.A1(G257), .A2(G1698), .ZN(new_n479));
  INV_X1    g0279(.A(G264), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n479), .B1(new_n480), .B2(G1698), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n478), .B1(new_n369), .B2(new_n481), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n473), .B(new_n476), .C1(new_n482), .C2(new_n405), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n462), .A2(new_n483), .A3(G169), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT21), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n480), .A2(G1698), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n487), .B1(G257), .B2(G1698), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n372), .A2(G33), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n278), .A2(KEYINPUT72), .ZN(new_n490));
  OAI21_X1  g0290(.A(KEYINPUT3), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n488), .B1(new_n491), .B2(new_n279), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n270), .B1(new_n492), .B2(new_n478), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n493), .A2(G190), .A3(new_n473), .A4(new_n476), .ZN(new_n494));
  AND2_X1   g0294(.A1(new_n457), .A2(new_n461), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n476), .A2(new_n473), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n277), .B1(new_n371), .B2(new_n373), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n481), .B1(new_n497), .B2(new_n308), .ZN(new_n498));
  INV_X1    g0298(.A(new_n478), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n405), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n494), .B(new_n495), .C1(new_n501), .C2(new_n303), .ZN(new_n502));
  NOR3_X1   g0302(.A1(new_n496), .A2(new_n500), .A3(new_n334), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n462), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n462), .A2(new_n483), .A3(KEYINPUT21), .A4(G169), .ZN(new_n505));
  AND4_X1   g0305(.A1(new_n486), .A2(new_n502), .A3(new_n504), .A4(new_n505), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n207), .B(G68), .C1(new_n497), .C2(new_n308), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT19), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n509), .B1(new_n256), .B2(new_n202), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(KEYINPUT78), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT78), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n512), .B(new_n509), .C1(new_n256), .C2(new_n202), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n207), .B1(new_n284), .B2(new_n509), .ZN(new_n514));
  INV_X1    g0314(.A(G87), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n515), .A2(new_n202), .A3(new_n203), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n511), .A2(new_n513), .A3(new_n517), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n259), .B1(new_n508), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n350), .A2(new_n250), .ZN(new_n520));
  INV_X1    g0320(.A(new_n350), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n460), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n519), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n465), .A2(new_n271), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n524), .B(new_n405), .C1(G250), .C2(new_n465), .ZN(new_n525));
  NOR2_X1   g0325(.A1(G238), .A2(G1698), .ZN(new_n526));
  INV_X1    g0326(.A(G244), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n526), .B1(new_n527), .B2(G1698), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n369), .A2(new_n528), .B1(G116), .B2(new_n374), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n525), .B1(new_n529), .B2(new_n405), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n344), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n528), .B1(new_n497), .B2(new_n308), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n374), .A2(G116), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n405), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n535), .A2(new_n334), .A3(new_n525), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n523), .A2(new_n531), .A3(new_n536), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n507), .A2(new_n513), .A3(new_n517), .A4(new_n511), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n538), .A2(new_n259), .B1(new_n250), .B2(new_n350), .ZN(new_n539));
  INV_X1    g0339(.A(new_n525), .ZN(new_n540));
  OAI21_X1  g0340(.A(G200), .B1(new_n534), .B2(new_n540), .ZN(new_n541));
  OAI211_X1 g0341(.A(G190), .B(new_n525), .C1(new_n529), .C2(new_n405), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n460), .A2(G87), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n539), .A2(new_n541), .A3(new_n542), .A4(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n537), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(KEYINPUT79), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n527), .A2(G1698), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n547), .B1(new_n497), .B2(new_n308), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT4), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AND2_X1   g0350(.A1(KEYINPUT4), .A2(G244), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n282), .B(new_n551), .C1(new_n307), .C2(new_n308), .ZN(new_n552));
  OAI211_X1 g0352(.A(G250), .B(G1698), .C1(new_n307), .C2(new_n308), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n552), .A2(new_n553), .A3(new_n448), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n405), .B1(new_n550), .B2(new_n555), .ZN(new_n556));
  OAI211_X1 g0356(.A(G257), .B(new_n405), .C1(new_n474), .C2(new_n475), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n473), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n344), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n389), .B1(KEYINPUT3), .B2(new_n374), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n390), .A2(new_n367), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n203), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(G97), .A2(G107), .ZN(new_n563));
  AOI21_X1  g0363(.A(KEYINPUT6), .B1(new_n204), .B2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT6), .ZN(new_n565));
  NOR3_X1   g0365(.A1(new_n565), .A2(new_n202), .A3(G107), .ZN(new_n566));
  OAI21_X1  g0366(.A(G20), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n253), .A2(G77), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n259), .B1(new_n562), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n460), .A2(G97), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n571), .B1(G97), .B2(new_n326), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n557), .A2(new_n473), .ZN(new_n575));
  AOI21_X1  g0375(.A(KEYINPUT4), .B1(new_n369), .B2(new_n547), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n270), .B1(new_n576), .B2(new_n554), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n575), .A2(new_n577), .A3(new_n334), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n559), .A2(new_n574), .A3(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(G200), .B1(new_n556), .B2(new_n558), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n575), .A2(new_n577), .A3(G190), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n568), .B(new_n567), .C1(new_n391), .C2(new_n203), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n572), .B1(new_n582), .B2(new_n259), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n580), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  AND2_X1   g0384(.A1(new_n579), .A2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT79), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n537), .A2(new_n544), .A3(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n506), .A2(new_n546), .A3(new_n585), .A4(new_n587), .ZN(new_n588));
  OAI211_X1 g0388(.A(G264), .B(new_n405), .C1(new_n474), .C2(new_n475), .ZN(new_n589));
  MUX2_X1   g0389(.A(G250), .B(G257), .S(G1698), .Z(new_n590));
  AOI22_X1  g0390(.A1(new_n369), .A2(new_n590), .B1(G294), .B2(new_n374), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n473), .B(new_n589), .C1(new_n591), .C2(new_n405), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n592), .A2(G179), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n593), .B1(new_n344), .B2(new_n592), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n207), .B(G87), .C1(new_n497), .C2(new_n308), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT81), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n595), .A2(new_n596), .A3(KEYINPUT22), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n596), .B1(new_n595), .B2(KEYINPUT22), .ZN(new_n598));
  NOR4_X1   g0398(.A1(new_n309), .A2(KEYINPUT22), .A3(G20), .A4(new_n515), .ZN(new_n599));
  NOR3_X1   g0399(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n374), .A2(new_n207), .A3(G116), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT23), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n602), .B1(G20), .B2(new_n203), .ZN(new_n603));
  NOR3_X1   g0403(.A1(new_n207), .A2(KEYINPUT23), .A3(G107), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AND3_X1   g0405(.A1(new_n601), .A2(KEYINPUT82), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(KEYINPUT82), .B1(new_n601), .B2(new_n605), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(KEYINPUT24), .B1(new_n600), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n595), .A2(KEYINPUT22), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(KEYINPUT81), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n595), .A2(new_n596), .A3(KEYINPUT22), .ZN(new_n612));
  INV_X1    g0412(.A(new_n599), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT24), .ZN(new_n615));
  INV_X1    g0415(.A(new_n608), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n354), .B1(new_n609), .B2(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(KEYINPUT25), .B1(new_n250), .B2(new_n203), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n250), .A2(KEYINPUT25), .A3(new_n203), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n620), .A2(new_n621), .B1(new_n460), .B2(G107), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n594), .B1(new_n618), .B2(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n599), .B1(new_n610), .B2(KEYINPUT81), .ZN(new_n625));
  AOI211_X1 g0425(.A(KEYINPUT24), .B(new_n608), .C1(new_n625), .C2(new_n612), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n615), .B1(new_n614), .B2(new_n616), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n259), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n592), .A2(new_n303), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n629), .B1(G190), .B2(new_n592), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n628), .A2(new_n622), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n624), .A2(new_n631), .ZN(new_n632));
  NOR3_X1   g0432(.A1(new_n445), .A2(new_n588), .A3(new_n632), .ZN(G372));
  INV_X1    g0433(.A(new_n337), .ZN(new_n634));
  INV_X1    g0434(.A(new_n299), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n635), .A2(new_n297), .A3(new_n296), .ZN(new_n636));
  INV_X1    g0436(.A(new_n358), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n269), .A2(new_n636), .B1(new_n305), .B2(new_n637), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n434), .B(new_n441), .C1(new_n638), .C2(KEYINPUT85), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n638), .A2(KEYINPUT85), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n426), .B(new_n440), .C1(new_n639), .C2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n634), .B1(new_n641), .B2(new_n330), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n525), .A2(KEYINPUT83), .ZN(new_n643));
  OR2_X1    g0443(.A1(new_n465), .A2(G250), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT83), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n644), .A2(new_n645), .A3(new_n405), .A4(new_n524), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n643), .B(new_n646), .C1(new_n529), .C2(new_n405), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n344), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n523), .A2(new_n648), .A3(new_n536), .ZN(new_n649));
  AND3_X1   g0449(.A1(new_n559), .A2(new_n578), .A3(new_n574), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n647), .A2(G200), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n651), .A2(new_n539), .A3(new_n542), .A4(new_n543), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n650), .A2(new_n649), .A3(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT26), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AND3_X1   g0455(.A1(new_n546), .A2(new_n650), .A3(new_n587), .ZN(new_n656));
  OAI211_X1 g0456(.A(new_n649), .B(new_n655), .C1(new_n656), .C2(new_n654), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT84), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n652), .A2(new_n649), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n631), .A2(new_n658), .A3(new_n585), .A4(new_n659), .ZN(new_n660));
  AND3_X1   g0460(.A1(new_n486), .A2(new_n504), .A3(new_n505), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n624), .A2(new_n661), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n631), .A2(new_n585), .A3(new_n659), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(KEYINPUT84), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n657), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n642), .B1(new_n445), .B2(new_n666), .ZN(G369));
  NAND2_X1  g0467(.A1(new_n628), .A2(new_n622), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n669));
  OR2_X1    g0469(.A1(new_n669), .A2(KEYINPUT27), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(KEYINPUT27), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(G213), .A3(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(G343), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n668), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(new_n631), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n624), .ZN(new_n677));
  INV_X1    g0477(.A(new_n674), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n668), .A2(new_n594), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g0480(.A(new_n680), .B(KEYINPUT86), .Z(new_n681));
  NAND2_X1  g0481(.A1(new_n462), .A2(new_n674), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n506), .A2(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n683), .B1(new_n661), .B2(new_n682), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n684), .A2(G330), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n681), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n661), .A2(new_n674), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n681), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n686), .A2(new_n688), .A3(new_n679), .ZN(G399));
  OR2_X1    g0489(.A1(new_n516), .A2(G116), .ZN(new_n690));
  XOR2_X1   g0490(.A(new_n690), .B(KEYINPUT87), .Z(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n223), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(G41), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n692), .A2(G1), .A3(new_n695), .ZN(new_n696));
  OAI22_X1  g0496(.A1(new_n696), .A2(KEYINPUT88), .B1(new_n228), .B2(new_n695), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n697), .B1(KEYINPUT88), .B2(new_n696), .ZN(new_n698));
  XOR2_X1   g0498(.A(new_n698), .B(KEYINPUT28), .Z(new_n699));
  XNOR2_X1  g0499(.A(new_n585), .B(KEYINPUT91), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n700), .A2(new_n662), .A3(new_n631), .A4(new_n659), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n649), .B1(new_n653), .B2(new_n654), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n702), .B1(new_n654), .B2(new_n656), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n674), .B1(new_n701), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(KEYINPUT29), .ZN(new_n705));
  OR2_X1    g0505(.A1(new_n705), .A2(KEYINPUT92), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n665), .A2(new_n662), .A3(new_n660), .ZN(new_n707));
  INV_X1    g0507(.A(new_n657), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(new_n678), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT29), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n705), .A2(KEYINPUT92), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n706), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n590), .B1(new_n497), .B2(new_n308), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n374), .A2(G294), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(new_n270), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n535), .A2(new_n718), .A3(new_n525), .A4(new_n589), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n493), .A2(G179), .A3(new_n473), .A4(new_n476), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n556), .A2(new_n558), .ZN(new_n722));
  AOI21_X1  g0522(.A(KEYINPUT30), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n589), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n405), .B1(new_n715), .B2(new_n716), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n534), .A2(new_n540), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n501), .A2(new_n726), .A3(G179), .A4(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n575), .A2(new_n577), .A3(KEYINPUT30), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n592), .A2(new_n647), .A3(new_n334), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n483), .B1(new_n556), .B2(new_n558), .ZN(new_n731));
  OAI22_X1  g0531(.A1(new_n728), .A2(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI211_X1 g0532(.A(KEYINPUT31), .B(new_n674), .C1(new_n723), .C2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n589), .B1(new_n591), .B2(new_n405), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(new_n530), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n736), .A2(new_n722), .A3(new_n503), .A4(KEYINPUT30), .ZN(new_n737));
  AND2_X1   g0537(.A1(new_n643), .A2(new_n646), .ZN(new_n738));
  AOI21_X1  g0538(.A(G179), .B1(new_n738), .B2(new_n535), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n554), .B1(new_n549), .B2(new_n548), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n473), .B(new_n557), .C1(new_n740), .C2(new_n405), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n739), .A2(new_n483), .A3(new_n741), .A4(new_n592), .ZN(new_n742));
  NOR3_X1   g0542(.A1(new_n719), .A2(new_n741), .A3(new_n720), .ZN(new_n743));
  OAI211_X1 g0543(.A(new_n737), .B(new_n742), .C1(new_n743), .C2(KEYINPUT30), .ZN(new_n744));
  AOI21_X1  g0544(.A(KEYINPUT31), .B1(new_n744), .B2(new_n674), .ZN(new_n745));
  OAI21_X1  g0545(.A(KEYINPUT89), .B1(new_n734), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n674), .B1(new_n723), .B2(new_n732), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT31), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT89), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n749), .A2(new_n750), .A3(new_n733), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n746), .A2(new_n751), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n632), .A2(new_n588), .A3(new_n674), .ZN(new_n753));
  OAI21_X1  g0553(.A(G330), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(KEYINPUT90), .ZN(new_n755));
  AND4_X1   g0555(.A1(new_n506), .A2(new_n546), .A3(new_n587), .A4(new_n585), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n756), .A2(new_n624), .A3(new_n631), .A4(new_n678), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n757), .A2(new_n746), .A3(new_n751), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT90), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n758), .A2(new_n759), .A3(G330), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n755), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n714), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n699), .B1(new_n764), .B2(G1), .ZN(G364));
  NOR2_X1   g0565(.A1(new_n249), .A2(G20), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n206), .B1(new_n766), .B2(G45), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n694), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G13), .A2(G33), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(G20), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  OR2_X1    g0574(.A1(new_n684), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n207), .A2(new_n301), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n776), .A2(new_n334), .A3(G200), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n281), .B1(new_n777), .B2(new_n515), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n207), .A2(G190), .ZN(new_n779));
  NOR2_X1   g0579(.A1(G179), .A2(G200), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G159), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  XOR2_X1   g0583(.A(new_n783), .B(KEYINPUT32), .Z(new_n784));
  AOI21_X1  g0584(.A(new_n207), .B1(new_n780), .B2(G190), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n778), .B(new_n784), .C1(G97), .C2(new_n786), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n207), .A2(new_n334), .A3(new_n303), .ZN(new_n788));
  OR2_X1    g0588(.A1(new_n788), .A2(KEYINPUT94), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(KEYINPUT94), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n789), .A2(G190), .A3(new_n790), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n789), .A2(new_n301), .A3(new_n790), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n787), .B1(new_n322), .B2(new_n791), .C1(new_n211), .C2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n334), .A2(G200), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n776), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n794), .A2(new_n779), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI22_X1  g0598(.A1(G58), .A2(new_n796), .B1(new_n798), .B2(G77), .ZN(new_n799));
  OR2_X1    g0599(.A1(new_n799), .A2(KEYINPUT93), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(KEYINPUT93), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n779), .A2(new_n334), .A3(G200), .ZN(new_n802));
  XOR2_X1   g0602(.A(new_n802), .B(KEYINPUT95), .Z(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(G107), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n800), .A2(new_n801), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n803), .A2(G283), .ZN(new_n806));
  INV_X1    g0606(.A(G322), .ZN(new_n807));
  INV_X1    g0607(.A(G311), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n795), .A2(new_n807), .B1(new_n797), .B2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n777), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n809), .B1(G303), .B2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(G294), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n785), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n781), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n281), .B(new_n813), .C1(G329), .C2(new_n814), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n806), .A2(new_n811), .A3(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(G326), .ZN(new_n817));
  XOR2_X1   g0617(.A(KEYINPUT33), .B(G317), .Z(new_n818));
  OAI22_X1  g0618(.A1(new_n817), .A2(new_n791), .B1(new_n792), .B2(new_n818), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n793), .A2(new_n805), .B1(new_n816), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n226), .B1(G20), .B2(new_n344), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n773), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n693), .A2(new_n309), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n823), .A2(G355), .B1(new_n446), .B2(new_n693), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n693), .A2(new_n369), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(G45), .B2(new_n228), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n247), .A2(new_n464), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n824), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n820), .A2(new_n821), .B1(new_n822), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n770), .B1(new_n775), .B2(new_n829), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n684), .B(G330), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n830), .B1(new_n770), .B2(new_n831), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n832), .B(KEYINPUT96), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(G396));
  NOR2_X1   g0634(.A1(new_n821), .A2(new_n771), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n769), .B1(new_n836), .B2(G77), .ZN(new_n837));
  AOI22_X1  g0637(.A1(G143), .A2(new_n796), .B1(new_n798), .B2(G159), .ZN(new_n838));
  INV_X1    g0638(.A(G150), .ZN(new_n839));
  INV_X1    g0639(.A(G137), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n838), .B1(new_n792), .B2(new_n839), .C1(new_n840), .C2(new_n791), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT34), .ZN(new_n842));
  OR2_X1    g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n841), .A2(new_n842), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n803), .A2(G68), .ZN(new_n845));
  INV_X1    g0645(.A(G132), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n777), .A2(new_n322), .B1(new_n781), .B2(new_n846), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n375), .B(new_n847), .C1(G58), .C2(new_n786), .ZN(new_n848));
  NAND4_X1  g0648(.A1(new_n843), .A2(new_n844), .A3(new_n845), .A4(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n803), .A2(G87), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n850), .B1(new_n808), .B2(new_n781), .ZN(new_n851));
  XNOR2_X1  g0651(.A(new_n851), .B(KEYINPUT98), .ZN(new_n852));
  INV_X1    g0652(.A(new_n792), .ZN(new_n853));
  INV_X1    g0653(.A(new_n791), .ZN(new_n854));
  AOI22_X1  g0654(.A1(G283), .A2(new_n853), .B1(new_n854), .B2(G303), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n281), .B1(new_n810), .B2(G107), .ZN(new_n856));
  OR2_X1    g0656(.A1(new_n856), .A2(KEYINPUT97), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(KEYINPUT97), .ZN(new_n858));
  OAI22_X1  g0658(.A1(new_n795), .A2(new_n812), .B1(new_n797), .B2(new_n446), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n859), .B1(G97), .B2(new_n786), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n855), .A2(new_n857), .A3(new_n858), .A4(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n849), .B1(new_n852), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n837), .B1(new_n862), .B2(new_n821), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n355), .A2(new_n674), .ZN(new_n864));
  INV_X1    g0664(.A(new_n343), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n345), .A2(KEYINPUT70), .B1(new_n865), .B2(new_n334), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n360), .B(new_n864), .C1(new_n866), .C2(new_n356), .ZN(new_n867));
  INV_X1    g0667(.A(new_n864), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n347), .A2(new_n357), .A3(new_n868), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n863), .B1(new_n871), .B2(new_n772), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n710), .A2(new_n870), .ZN(new_n873));
  INV_X1    g0673(.A(new_n361), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n678), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n873), .B1(new_n666), .B2(new_n875), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n876), .A2(new_n762), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(KEYINPUT99), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n878), .B(new_n770), .C1(new_n762), .C2(new_n876), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n877), .A2(KEYINPUT99), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n872), .B1(new_n879), .B2(new_n880), .ZN(G384));
  NOR2_X1   g0681(.A1(new_n766), .A2(new_n206), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT39), .ZN(new_n883));
  OR2_X1    g0683(.A1(new_n398), .A2(KEYINPUT16), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n366), .B1(new_n884), .B2(new_n399), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n885), .A2(new_n672), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n426), .A2(new_n440), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n434), .A2(new_n441), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n886), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n435), .A2(new_n439), .ZN(new_n890));
  INV_X1    g0690(.A(new_n672), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n435), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT37), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n890), .A2(new_n892), .A3(new_n893), .A4(new_n432), .ZN(new_n894));
  INV_X1    g0694(.A(new_n432), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n885), .B1(new_n425), .B2(new_n672), .ZN(new_n896));
  OAI21_X1  g0696(.A(KEYINPUT37), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  AND3_X1   g0698(.A1(new_n889), .A2(KEYINPUT38), .A3(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n432), .B1(new_n425), .B2(new_n402), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n402), .A2(new_n672), .ZN(new_n901));
  OAI21_X1  g0701(.A(KEYINPUT37), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n894), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n442), .A2(new_n901), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT38), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n883), .B1(new_n899), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n889), .A2(new_n898), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT38), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n889), .A2(KEYINPUT38), .A3(new_n898), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n909), .A2(KEYINPUT39), .A3(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n636), .A2(new_n269), .A3(new_n678), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n906), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n909), .A2(new_n910), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n637), .A2(new_n678), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n875), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n917), .B1(new_n709), .B2(new_n918), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n300), .B(new_n305), .C1(new_n268), .C2(new_n678), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n302), .A2(new_n304), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n269), .B(new_n674), .C1(new_n636), .C2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n919), .A2(new_n924), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n915), .A2(new_n925), .B1(new_n887), .B2(new_n672), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n914), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g0727(.A1(new_n706), .A2(new_n444), .A3(new_n712), .A4(new_n713), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n642), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n927), .B(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n870), .B1(new_n920), .B2(new_n922), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n749), .B1(new_n734), .B2(KEYINPUT101), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT101), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n747), .A2(new_n933), .A3(new_n748), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n757), .A2(new_n932), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n931), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n903), .A2(new_n904), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n908), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n936), .B1(new_n938), .B2(new_n910), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT40), .ZN(new_n940));
  AOI21_X1  g0740(.A(KEYINPUT38), .B1(new_n889), .B2(new_n898), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n899), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n931), .A2(new_n940), .A3(new_n935), .ZN(new_n943));
  OAI22_X1  g0743(.A1(new_n939), .A2(new_n940), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n944), .A2(new_n444), .A3(new_n935), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n894), .A2(new_n902), .B1(new_n442), .B2(new_n901), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n910), .B1(new_n946), .B2(KEYINPUT38), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n931), .A2(new_n935), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n940), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n943), .B1(new_n909), .B2(new_n910), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n444), .A2(new_n935), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n945), .A2(new_n953), .A3(G330), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n882), .B1(new_n930), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n930), .B2(new_n954), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n564), .A2(new_n566), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n958), .A2(KEYINPUT35), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(KEYINPUT35), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n959), .A2(G116), .A3(new_n227), .A4(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT36), .ZN(new_n962));
  NOR3_X1   g0762(.A1(new_n384), .A2(new_n228), .A3(new_n255), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n963), .A2(KEYINPUT100), .B1(new_n322), .B2(G68), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(KEYINPUT100), .B2(new_n963), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n965), .A2(G1), .A3(new_n249), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n956), .A2(new_n962), .A3(new_n966), .ZN(G367));
  OAI21_X1  g0767(.A(new_n700), .B1(new_n583), .B2(new_n678), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n968), .A2(new_n624), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n674), .B1(new_n969), .B2(new_n579), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n650), .A2(new_n674), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n681), .A2(new_n687), .A3(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT42), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n973), .A2(new_n974), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n970), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT102), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n539), .A2(new_n543), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n674), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n659), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n649), .B2(new_n980), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n982), .B(KEYINPUT43), .Z(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  OR3_X1    g0784(.A1(new_n977), .A2(new_n978), .A3(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n978), .B1(new_n977), .B2(new_n984), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n977), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n985), .A2(new_n986), .A3(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n972), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n686), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n989), .B(new_n991), .ZN(new_n992));
  XNOR2_X1  g0792(.A(KEYINPUT103), .B(KEYINPUT41), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n694), .B(new_n993), .Z(new_n994));
  NAND3_X1  g0794(.A1(new_n688), .A2(new_n679), .A3(new_n972), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT45), .Z(new_n996));
  AOI21_X1  g0796(.A(new_n972), .B1(new_n688), .B2(new_n679), .ZN(new_n997));
  OR2_X1    g0797(.A1(KEYINPUT104), .A2(KEYINPUT44), .ZN(new_n998));
  AND2_X1   g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(KEYINPUT104), .A2(KEYINPUT44), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n997), .B2(new_n998), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n996), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n686), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n996), .B(new_n686), .C1(new_n999), .C2(new_n1001), .ZN(new_n1005));
  OAI21_X1  g0805(.A(KEYINPUT105), .B1(new_n681), .B2(new_n687), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(new_n688), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT106), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n685), .A2(new_n1008), .ZN(new_n1009));
  AND2_X1   g0809(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1004), .A2(new_n764), .A3(new_n1005), .A4(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n994), .B1(new_n1013), .B2(new_n764), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n992), .B1(new_n1014), .B2(new_n768), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n825), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n240), .A2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n822), .B1(new_n223), .B2(new_n350), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n769), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n777), .A2(new_n383), .B1(new_n781), .B2(new_n840), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n802), .A2(new_n255), .B1(new_n797), .B2(new_n322), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n281), .B1(new_n795), .B2(new_n839), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n785), .A2(new_n211), .ZN(new_n1023));
  NOR4_X1   g0823(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(G143), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1024), .B1(new_n1025), .B2(new_n791), .C1(new_n782), .C2(new_n792), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n375), .B1(new_n203), .B2(new_n785), .ZN(new_n1027));
  INV_X1    g0827(.A(G317), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n802), .A2(new_n202), .B1(new_n781), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(G283), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n795), .A2(new_n477), .B1(new_n797), .B2(new_n1030), .ZN(new_n1031));
  NOR3_X1   g0831(.A1(new_n1027), .A2(new_n1029), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT46), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n777), .B2(new_n446), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n810), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1034), .B(new_n1035), .C1(new_n792), .C2(new_n812), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n1032), .B1(new_n808), .B2(new_n791), .C1(new_n1036), .C2(KEYINPUT107), .ZN(new_n1037));
  AND2_X1   g0837(.A1(new_n1036), .A2(KEYINPUT107), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1026), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT47), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1019), .B1(new_n1040), .B2(new_n821), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n774), .B2(new_n982), .ZN(new_n1042));
  AND2_X1   g0842(.A1(new_n1015), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(G387));
  NOR2_X1   g0844(.A1(new_n681), .A2(new_n774), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n692), .B(new_n464), .C1(new_n211), .C2(new_n255), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n352), .A2(new_n322), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT50), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n825), .B1(new_n464), .B2(new_n236), .C1(new_n1046), .C2(new_n1048), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n691), .A2(new_n823), .B1(new_n203), .B2(new_n693), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1049), .A2(KEYINPUT108), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n822), .ZN(new_n1052));
  AOI21_X1  g0852(.A(KEYINPUT108), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n769), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n802), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n1055), .A2(G116), .B1(new_n814), .B2(G326), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n777), .A2(new_n812), .B1(new_n785), .B2(new_n1030), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(G317), .A2(new_n796), .B1(new_n798), .B2(G303), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1058), .B1(new_n792), .B2(new_n808), .C1(new_n807), .C2(new_n791), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT110), .Z(new_n1060));
  AOI21_X1  g0860(.A(new_n1057), .B1(new_n1060), .B2(KEYINPUT48), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT111), .Z(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(KEYINPUT48), .B2(new_n1060), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT49), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n375), .B(new_n1056), .C1(new_n1063), .C2(new_n1064), .ZN(new_n1065));
  AND2_X1   g0865(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n803), .A2(G97), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n777), .A2(new_n255), .B1(new_n795), .B2(new_n322), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(KEYINPUT109), .B(G150), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n797), .A2(new_n211), .B1(new_n781), .B2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n785), .A2(new_n350), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n375), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1067), .A2(new_n1071), .A3(new_n1073), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n782), .A2(new_n791), .B1(new_n792), .B2(new_n319), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n1065), .A2(new_n1066), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT112), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n1045), .B(new_n1054), .C1(new_n1077), .C2(new_n821), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(new_n1012), .B2(new_n768), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1012), .A2(new_n764), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n694), .B(KEYINPUT113), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n763), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1080), .B(new_n1081), .C1(new_n1082), .C2(KEYINPUT114), .ZN(new_n1083));
  AND2_X1   g0883(.A1(new_n1082), .A2(KEYINPUT114), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1079), .B1(new_n1083), .B2(new_n1084), .ZN(G393));
  NAND2_X1  g0885(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n990), .A2(new_n773), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n822), .B1(new_n202), .B2(new_n223), .C1(new_n1016), .C2(new_n244), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n769), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n791), .A2(new_n1028), .B1(new_n808), .B2(new_n795), .ZN(new_n1091));
  XOR2_X1   g0891(.A(new_n1091), .B(KEYINPUT52), .Z(new_n1092));
  OAI22_X1  g0892(.A1(new_n777), .A2(new_n1030), .B1(new_n797), .B2(new_n812), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n281), .B(new_n1093), .C1(G322), .C2(new_n814), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n853), .A2(G303), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n786), .A2(G116), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n1094), .A2(new_n804), .A3(new_n1095), .A4(new_n1096), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n791), .A2(new_n839), .B1(new_n782), .B2(new_n795), .ZN(new_n1098));
  XOR2_X1   g0898(.A(new_n1098), .B(KEYINPUT51), .Z(new_n1099));
  NAND2_X1  g0899(.A1(new_n853), .A2(G50), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n777), .A2(new_n211), .B1(new_n781), .B2(new_n1025), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n785), .A2(new_n255), .ZN(new_n1102));
  NOR3_X1   g0902(.A1(new_n1101), .A2(new_n375), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n352), .A2(new_n798), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n1100), .A2(new_n850), .A3(new_n1103), .A4(new_n1104), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n1092), .A2(new_n1097), .B1(new_n1099), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1090), .B1(new_n1106), .B2(new_n821), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n1087), .A2(new_n768), .B1(new_n1088), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1086), .A2(new_n1080), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1109), .A2(new_n1013), .A3(new_n1081), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1108), .A2(new_n1110), .ZN(G390));
  OAI21_X1  g0911(.A(new_n916), .B1(new_n666), .B2(new_n875), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n913), .B1(new_n1112), .B2(new_n923), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(KEYINPUT39), .B1(new_n938), .B2(new_n910), .ZN(new_n1115));
  NOR3_X1   g0915(.A1(new_n899), .A2(new_n941), .A3(new_n883), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1114), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  AND3_X1   g0917(.A1(new_n758), .A2(new_n759), .A3(G330), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n759), .B1(new_n758), .B2(G330), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n931), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(KEYINPUT115), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT115), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1122), .B(new_n931), .C1(new_n1118), .C2(new_n1119), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n674), .B(new_n870), .C1(new_n703), .C2(new_n701), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n923), .B1(new_n1125), .B2(new_n917), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1126), .A2(new_n947), .A3(new_n912), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1117), .A2(new_n1124), .A3(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n935), .A2(G330), .ZN(new_n1129));
  NOR3_X1   g0929(.A1(new_n924), .A2(new_n1129), .A3(new_n870), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1113), .B1(new_n906), .B2(new_n911), .ZN(new_n1131));
  AND3_X1   g0931(.A1(new_n1126), .A2(new_n947), .A3(new_n912), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1130), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  AND2_X1   g0933(.A1(new_n1128), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT117), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n772), .B1(new_n906), .B2(new_n911), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n821), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(G128), .A2(new_n854), .B1(new_n853), .B2(G137), .ZN(new_n1138));
  INV_X1    g0938(.A(G125), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n795), .A2(new_n846), .B1(new_n781), .B2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(G50), .B2(new_n1055), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n777), .A2(new_n1069), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT53), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(KEYINPUT54), .B(G143), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n281), .B1(new_n797), .B2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n1142), .A2(new_n1143), .B1(G159), .B2(new_n786), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1138), .A2(new_n1141), .A3(new_n1147), .A4(new_n1148), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(G107), .A2(new_n853), .B1(new_n854), .B2(G283), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n797), .A2(new_n202), .B1(new_n781), .B2(new_n812), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(G116), .B2(new_n796), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n281), .B(new_n1102), .C1(G87), .C2(new_n810), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1150), .A2(new_n845), .A3(new_n1152), .A4(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1137), .B1(new_n1149), .B2(new_n1154), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n770), .B(new_n1155), .C1(new_n319), .C2(new_n835), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1156), .B(KEYINPUT116), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1135), .B1(new_n1136), .B2(new_n1157), .ZN(new_n1158));
  OR3_X1    g0958(.A1(new_n1136), .A2(new_n1135), .A3(new_n1157), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n1134), .A2(new_n768), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n935), .A2(G330), .A3(new_n871), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n917), .B(new_n1125), .C1(new_n1161), .C2(new_n924), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1122), .B1(new_n761), .B2(new_n931), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1123), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1162), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n923), .B1(new_n761), .B2(new_n871), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1112), .B1(new_n1166), .B2(new_n1130), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n444), .A2(G330), .A3(new_n935), .ZN(new_n1169));
  AND3_X1   g0969(.A1(new_n928), .A2(new_n642), .A3(new_n1169), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n1168), .A2(new_n1170), .B1(new_n1128), .B2(new_n1133), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1168), .A2(new_n1128), .A3(new_n1133), .A4(new_n1170), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(new_n1081), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1160), .B1(new_n1171), .B2(new_n1173), .ZN(G378));
  NAND2_X1  g0974(.A1(new_n327), .A2(new_n891), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1175), .B(KEYINPUT118), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n338), .B(new_n1176), .ZN(new_n1177));
  XOR2_X1   g0977(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1178));
  XOR2_X1   g0978(.A(new_n1177), .B(new_n1178), .Z(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(G330), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1180), .B1(new_n951), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n927), .ZN(new_n1183));
  OAI211_X1 g0983(.A(G330), .B(new_n1179), .C1(new_n949), .C2(new_n950), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1179), .B1(new_n944), .B2(G330), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1184), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT119), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n927), .A2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n914), .A2(new_n926), .A3(KEYINPUT119), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1185), .B1(new_n1188), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1172), .A2(new_n1170), .ZN(new_n1194));
  AOI21_X1  g0994(.A(KEYINPUT57), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT120), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1190), .B(new_n1191), .C1(new_n1186), .C2(new_n1187), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n1198), .A2(new_n1185), .B1(new_n1172), .B2(new_n1170), .ZN(new_n1199));
  OAI21_X1  g0999(.A(KEYINPUT120), .B1(new_n1199), .B2(KEYINPUT57), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1081), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT57), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(new_n1172), .B2(new_n1170), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n927), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(new_n1185), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1201), .B1(new_n1203), .B2(new_n1205), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1197), .A2(new_n1200), .A3(new_n1206), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n369), .A2(G41), .ZN(new_n1208));
  AOI211_X1 g1008(.A(G50), .B(new_n1208), .C1(new_n278), .C2(new_n404), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n796), .A2(G107), .B1(new_n798), .B2(new_n521), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1210), .B1(new_n1030), .B2(new_n781), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n777), .A2(new_n255), .B1(new_n802), .B2(new_n383), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(new_n1211), .A2(new_n1023), .A3(new_n1212), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(G97), .A2(new_n853), .B1(new_n854), .B2(G116), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1213), .A2(new_n1214), .A3(new_n1208), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT58), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1209), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n785), .A2(new_n839), .ZN(new_n1218));
  INV_X1    g1018(.A(G128), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n777), .A2(new_n1145), .B1(new_n795), .B2(new_n1219), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n1218), .B(new_n1220), .C1(G137), .C2(new_n798), .ZN(new_n1221));
  OAI221_X1 g1021(.A(new_n1221), .B1(new_n1139), .B2(new_n791), .C1(new_n846), .C2(new_n792), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1222), .B(KEYINPUT59), .ZN(new_n1223));
  AOI211_X1 g1023(.A(G33), .B(G41), .C1(new_n1055), .C2(G159), .ZN(new_n1224));
  INV_X1    g1024(.A(G124), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1224), .B1(new_n1225), .B2(new_n781), .ZN(new_n1226));
  OAI221_X1 g1026(.A(new_n1217), .B1(new_n1216), .B2(new_n1215), .C1(new_n1223), .C2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(new_n821), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n1228), .B(new_n769), .C1(G50), .C2(new_n836), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(new_n1180), .B2(new_n771), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(new_n1193), .B2(new_n768), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1207), .A2(new_n1231), .ZN(G375));
  OR2_X1    g1032(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n994), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1233), .A2(new_n1234), .A3(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n924), .A2(new_n771), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n769), .B1(new_n836), .B2(G68), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n803), .A2(G77), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n795), .A2(new_n1030), .B1(new_n797), .B2(new_n203), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(G303), .B2(new_n814), .ZN(new_n1241));
  AOI211_X1 g1041(.A(new_n281), .B(new_n1072), .C1(G97), .C2(new_n810), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1239), .A2(new_n1241), .A3(new_n1242), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n446), .A2(new_n792), .B1(new_n791), .B2(new_n812), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n777), .A2(new_n782), .B1(new_n781), .B2(new_n1219), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(G137), .B2(new_n796), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n786), .A2(G50), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(G58), .A2(new_n1055), .B1(new_n798), .B2(G150), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1246), .A2(new_n369), .A3(new_n1247), .A4(new_n1248), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n846), .A2(new_n791), .B1(new_n792), .B2(new_n1145), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n1243), .A2(new_n1244), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1238), .B1(new_n1251), .B2(new_n821), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n1168), .A2(new_n768), .B1(new_n1237), .B2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1236), .A2(new_n1253), .ZN(G381));
  OR2_X1    g1054(.A1(G381), .A2(G384), .ZN(new_n1255));
  NOR4_X1   g1055(.A1(G390), .A2(G396), .A3(G393), .A4(new_n1255), .ZN(new_n1256));
  XNOR2_X1  g1056(.A(G378), .B(KEYINPUT121), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1256), .A2(new_n1043), .A3(new_n1258), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1259), .A2(G375), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT122), .ZN(new_n1261));
  XNOR2_X1  g1061(.A(new_n1260), .B(new_n1261), .ZN(G407));
  NAND2_X1  g1062(.A1(new_n1258), .A2(new_n673), .ZN(new_n1263));
  OAI211_X1 g1063(.A(G407), .B(G213), .C1(G375), .C2(new_n1263), .ZN(G409));
  AOI21_X1  g1064(.A(new_n767), .B1(new_n1204), .B2(new_n1185), .ZN(new_n1265));
  OAI21_X1  g1065(.A(KEYINPUT124), .B1(new_n1265), .B2(new_n1230), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1199), .A2(new_n1234), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  NOR3_X1   g1068(.A1(new_n1265), .A2(KEYINPUT124), .A3(new_n1230), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1257), .A2(new_n1270), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1206), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1272));
  NOR3_X1   g1072(.A1(new_n1199), .A2(KEYINPUT120), .A3(KEYINPUT57), .ZN(new_n1273));
  OAI211_X1 g1073(.A(G378), .B(new_n1231), .C1(new_n1272), .C2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(KEYINPUT123), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT123), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1207), .A2(new_n1276), .A3(G378), .A4(new_n1231), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1271), .B1(new_n1275), .B2(new_n1277), .ZN(new_n1278));
  AND2_X1   g1078(.A1(new_n673), .A2(G213), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT60), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1233), .A2(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1281), .A2(new_n1081), .A3(new_n1235), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1233), .A2(new_n1280), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1253), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  XNOR2_X1  g1084(.A(new_n1284), .B(G384), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  NOR3_X1   g1086(.A1(new_n1278), .A2(new_n1279), .A3(new_n1286), .ZN(new_n1287));
  OR2_X1    g1087(.A1(new_n1287), .A2(KEYINPUT63), .ZN(new_n1288));
  AND3_X1   g1088(.A1(new_n1015), .A2(G390), .A3(new_n1042), .ZN(new_n1289));
  AOI21_X1  g1089(.A(G390), .B1(new_n1015), .B2(new_n1042), .ZN(new_n1290));
  OAI21_X1  g1090(.A(KEYINPUT125), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  XNOR2_X1  g1091(.A(G393), .B(new_n833), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1291), .A2(new_n1293), .ZN(new_n1294));
  OAI211_X1 g1094(.A(KEYINPUT125), .B(new_n1292), .C1(new_n1289), .C2(new_n1290), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT61), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1275), .A2(new_n1277), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1271), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1279), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1279), .A2(G2897), .ZN(new_n1301));
  XNOR2_X1  g1101(.A(new_n1285), .B(new_n1301), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1297), .B1(new_n1300), .B2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1287), .A2(KEYINPUT63), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1288), .A2(new_n1296), .A3(new_n1304), .A4(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT62), .ZN(new_n1307));
  NOR4_X1   g1107(.A1(new_n1278), .A2(new_n1307), .A3(new_n1286), .A4(new_n1279), .ZN(new_n1308));
  XNOR2_X1  g1108(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1309), .B1(new_n1300), .B2(new_n1285), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT127), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1308), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  OAI21_X1  g1112(.A(KEYINPUT127), .B1(new_n1287), .B2(new_n1309), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1303), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1306), .B1(new_n1314), .B2(new_n1296), .ZN(G405));
  NAND2_X1  g1115(.A1(new_n1258), .A2(G375), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1298), .A2(new_n1316), .ZN(new_n1317));
  XNOR2_X1  g1117(.A(new_n1317), .B(new_n1286), .ZN(new_n1318));
  XNOR2_X1  g1118(.A(new_n1296), .B(new_n1318), .ZN(G402));
endmodule


