

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591;

  XNOR2_X1 U325 ( .A(n384), .B(KEYINPUT31), .ZN(n385) );
  XNOR2_X1 U326 ( .A(n386), .B(n385), .ZN(n389) );
  XNOR2_X1 U327 ( .A(n412), .B(n396), .ZN(n397) );
  XNOR2_X1 U328 ( .A(n398), .B(n397), .ZN(n586) );
  XNOR2_X1 U329 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U330 ( .A(n452), .B(n451), .ZN(G1351GAT) );
  XOR2_X1 U331 ( .A(KEYINPUT0), .B(G134GAT), .Z(n294) );
  XNOR2_X1 U332 ( .A(KEYINPUT78), .B(G127GAT), .ZN(n293) );
  XNOR2_X1 U333 ( .A(n294), .B(n293), .ZN(n295) );
  XNOR2_X1 U334 ( .A(G113GAT), .B(n295), .ZN(n434) );
  XOR2_X1 U335 ( .A(KEYINPUT89), .B(KEYINPUT1), .Z(n297) );
  XNOR2_X1 U336 ( .A(KEYINPUT88), .B(KEYINPUT5), .ZN(n296) );
  XNOR2_X1 U337 ( .A(n297), .B(n296), .ZN(n312) );
  XOR2_X1 U338 ( .A(G155GAT), .B(G148GAT), .Z(n299) );
  XNOR2_X1 U339 ( .A(G29GAT), .B(G120GAT), .ZN(n298) );
  XNOR2_X1 U340 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U341 ( .A(G57GAT), .B(KEYINPUT6), .Z(n301) );
  XNOR2_X1 U342 ( .A(G1GAT), .B(KEYINPUT4), .ZN(n300) );
  XNOR2_X1 U343 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U344 ( .A(n303), .B(n302), .Z(n310) );
  XOR2_X1 U345 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n305) );
  XNOR2_X1 U346 ( .A(G141GAT), .B(KEYINPUT85), .ZN(n304) );
  XNOR2_X1 U347 ( .A(n305), .B(n304), .ZN(n418) );
  XOR2_X1 U348 ( .A(G85GAT), .B(G162GAT), .Z(n307) );
  NAND2_X1 U349 ( .A1(G225GAT), .A2(G233GAT), .ZN(n306) );
  XNOR2_X1 U350 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U351 ( .A(n418), .B(n308), .ZN(n309) );
  XNOR2_X1 U352 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U353 ( .A(n312), .B(n311), .Z(n313) );
  XOR2_X1 U354 ( .A(n434), .B(n313), .Z(n543) );
  XOR2_X1 U355 ( .A(G211GAT), .B(KEYINPUT84), .Z(n315) );
  XNOR2_X1 U356 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n314) );
  XNOR2_X1 U357 ( .A(n315), .B(n314), .ZN(n417) );
  XNOR2_X1 U358 ( .A(G176GAT), .B(G92GAT), .ZN(n321) );
  INV_X1 U359 ( .A(KEYINPUT73), .ZN(n316) );
  NAND2_X1 U360 ( .A1(G64GAT), .A2(n316), .ZN(n319) );
  INV_X1 U361 ( .A(G64GAT), .ZN(n317) );
  NAND2_X1 U362 ( .A1(n317), .A2(KEYINPUT73), .ZN(n318) );
  NAND2_X1 U363 ( .A1(n319), .A2(n318), .ZN(n320) );
  XNOR2_X1 U364 ( .A(n321), .B(n320), .ZN(n383) );
  XNOR2_X1 U365 ( .A(n417), .B(n383), .ZN(n326) );
  XNOR2_X1 U366 ( .A(G36GAT), .B(G190GAT), .ZN(n322) );
  XNOR2_X1 U367 ( .A(n322), .B(G218GAT), .ZN(n377) );
  XOR2_X1 U368 ( .A(n377), .B(KEYINPUT90), .Z(n324) );
  NAND2_X1 U369 ( .A1(G226GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U370 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U371 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U372 ( .A(n327), .B(KEYINPUT91), .Z(n329) );
  XOR2_X1 U373 ( .A(G169GAT), .B(G8GAT), .Z(n334) );
  XNOR2_X1 U374 ( .A(n334), .B(G204GAT), .ZN(n328) );
  XNOR2_X1 U375 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U376 ( .A(KEYINPUT18), .B(KEYINPUT19), .Z(n331) );
  XNOR2_X1 U377 ( .A(KEYINPUT81), .B(G183GAT), .ZN(n330) );
  XNOR2_X1 U378 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U379 ( .A(KEYINPUT17), .B(n332), .ZN(n444) );
  XOR2_X1 U380 ( .A(n333), .B(n444), .Z(n533) );
  INV_X1 U381 ( .A(n533), .ZN(n515) );
  XOR2_X1 U382 ( .A(G141GAT), .B(G113GAT), .Z(n336) );
  XNOR2_X1 U383 ( .A(G15GAT), .B(G1GAT), .ZN(n352) );
  XOR2_X1 U384 ( .A(n334), .B(n352), .Z(n335) );
  XNOR2_X1 U385 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U386 ( .A(n337), .B(G36GAT), .Z(n342) );
  XOR2_X1 U387 ( .A(KEYINPUT68), .B(KEYINPUT29), .Z(n339) );
  XNOR2_X1 U388 ( .A(G197GAT), .B(G22GAT), .ZN(n338) );
  XNOR2_X1 U389 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U390 ( .A(n340), .B(G50GAT), .ZN(n341) );
  XNOR2_X1 U391 ( .A(n342), .B(n341), .ZN(n346) );
  XOR2_X1 U392 ( .A(KEYINPUT30), .B(KEYINPUT65), .Z(n344) );
  NAND2_X1 U393 ( .A1(G229GAT), .A2(G233GAT), .ZN(n343) );
  XNOR2_X1 U394 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U395 ( .A(n346), .B(n345), .Z(n351) );
  XOR2_X1 U396 ( .A(KEYINPUT7), .B(KEYINPUT67), .Z(n348) );
  XNOR2_X1 U397 ( .A(G43GAT), .B(G29GAT), .ZN(n347) );
  XNOR2_X1 U398 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U399 ( .A(KEYINPUT8), .B(n349), .ZN(n380) );
  XOR2_X1 U400 ( .A(n380), .B(KEYINPUT66), .Z(n350) );
  XOR2_X1 U401 ( .A(n351), .B(n350), .Z(n508) );
  INV_X1 U402 ( .A(n508), .ZN(n581) );
  XNOR2_X1 U403 ( .A(G183GAT), .B(G71GAT), .ZN(n353) );
  XNOR2_X1 U404 ( .A(n353), .B(n352), .ZN(n366) );
  XOR2_X1 U405 ( .A(G57GAT), .B(KEYINPUT13), .Z(n395) );
  XOR2_X1 U406 ( .A(n395), .B(KEYINPUT14), .Z(n355) );
  NAND2_X1 U407 ( .A1(G231GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U408 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U409 ( .A(KEYINPUT15), .B(KEYINPUT76), .Z(n357) );
  XNOR2_X1 U410 ( .A(G64GAT), .B(KEYINPUT12), .ZN(n356) );
  XNOR2_X1 U411 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U412 ( .A(n359), .B(n358), .Z(n364) );
  XOR2_X1 U413 ( .A(G22GAT), .B(G155GAT), .Z(n413) );
  XOR2_X1 U414 ( .A(G211GAT), .B(G78GAT), .Z(n361) );
  XNOR2_X1 U415 ( .A(G8GAT), .B(G127GAT), .ZN(n360) );
  XNOR2_X1 U416 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U417 ( .A(n413), .B(n362), .ZN(n363) );
  XNOR2_X1 U418 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U419 ( .A(n366), .B(n365), .Z(n590) );
  INV_X1 U420 ( .A(n590), .ZN(n490) );
  XOR2_X1 U421 ( .A(G50GAT), .B(G162GAT), .Z(n414) );
  XOR2_X1 U422 ( .A(KEYINPUT75), .B(KEYINPUT74), .Z(n368) );
  XNOR2_X1 U423 ( .A(KEYINPUT11), .B(KEYINPUT9), .ZN(n367) );
  XNOR2_X1 U424 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U425 ( .A(n414), .B(n369), .Z(n371) );
  NAND2_X1 U426 ( .A1(G232GAT), .A2(G233GAT), .ZN(n370) );
  XNOR2_X1 U427 ( .A(n371), .B(n370), .ZN(n375) );
  XOR2_X1 U428 ( .A(KEYINPUT10), .B(G92GAT), .Z(n373) );
  XNOR2_X1 U429 ( .A(G134GAT), .B(G106GAT), .ZN(n372) );
  XNOR2_X1 U430 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U431 ( .A(n375), .B(n374), .Z(n379) );
  XNOR2_X1 U432 ( .A(G99GAT), .B(G85GAT), .ZN(n376) );
  XNOR2_X1 U433 ( .A(n376), .B(KEYINPUT71), .ZN(n387) );
  XNOR2_X1 U434 ( .A(n377), .B(n387), .ZN(n378) );
  XNOR2_X1 U435 ( .A(n379), .B(n378), .ZN(n381) );
  XNOR2_X1 U436 ( .A(n381), .B(n380), .ZN(n461) );
  INV_X1 U437 ( .A(n461), .ZN(n569) );
  XOR2_X1 U438 ( .A(n569), .B(KEYINPUT36), .Z(n489) );
  NOR2_X1 U439 ( .A1(n490), .A2(n489), .ZN(n382) );
  XNOR2_X1 U440 ( .A(KEYINPUT45), .B(n382), .ZN(n399) );
  XOR2_X1 U441 ( .A(G120GAT), .B(G71GAT), .Z(n430) );
  XNOR2_X1 U442 ( .A(n383), .B(n430), .ZN(n386) );
  AND2_X1 U443 ( .A1(G230GAT), .A2(G233GAT), .ZN(n384) );
  XOR2_X1 U444 ( .A(n387), .B(KEYINPUT32), .Z(n388) );
  XNOR2_X1 U445 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U446 ( .A(n390), .B(KEYINPUT72), .ZN(n398) );
  XOR2_X1 U447 ( .A(KEYINPUT70), .B(KEYINPUT69), .Z(n392) );
  XNOR2_X1 U448 ( .A(G78GAT), .B(G148GAT), .ZN(n391) );
  XNOR2_X1 U449 ( .A(n392), .B(n391), .ZN(n394) );
  XOR2_X1 U450 ( .A(G106GAT), .B(G204GAT), .Z(n393) );
  XOR2_X1 U451 ( .A(n394), .B(n393), .Z(n412) );
  XOR2_X1 U452 ( .A(n395), .B(KEYINPUT33), .Z(n396) );
  INV_X1 U453 ( .A(n586), .ZN(n460) );
  NAND2_X1 U454 ( .A1(n399), .A2(n460), .ZN(n400) );
  NOR2_X1 U455 ( .A1(n581), .A2(n400), .ZN(n401) );
  XOR2_X1 U456 ( .A(KEYINPUT115), .B(n401), .Z(n408) );
  INV_X1 U457 ( .A(KEYINPUT41), .ZN(n402) );
  XNOR2_X1 U458 ( .A(n402), .B(n586), .ZN(n573) );
  NAND2_X1 U459 ( .A1(n581), .A2(n573), .ZN(n403) );
  XNOR2_X1 U460 ( .A(n403), .B(KEYINPUT46), .ZN(n404) );
  NAND2_X1 U461 ( .A1(n404), .A2(n490), .ZN(n405) );
  NOR2_X1 U462 ( .A1(n569), .A2(n405), .ZN(n406) );
  XOR2_X1 U463 ( .A(KEYINPUT47), .B(n406), .Z(n407) );
  NOR2_X1 U464 ( .A1(n408), .A2(n407), .ZN(n409) );
  XNOR2_X1 U465 ( .A(KEYINPUT48), .B(n409), .ZN(n542) );
  NOR2_X1 U466 ( .A1(n515), .A2(n542), .ZN(n410) );
  XNOR2_X1 U467 ( .A(n410), .B(KEYINPUT54), .ZN(n411) );
  AND2_X1 U468 ( .A1(n543), .A2(n411), .ZN(n455) );
  INV_X1 U469 ( .A(n412), .ZN(n428) );
  XOR2_X1 U470 ( .A(KEYINPUT87), .B(G218GAT), .Z(n416) );
  XNOR2_X1 U471 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U472 ( .A(n416), .B(n415), .ZN(n424) );
  XNOR2_X1 U473 ( .A(n418), .B(n417), .ZN(n422) );
  XOR2_X1 U474 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n420) );
  XNOR2_X1 U475 ( .A(KEYINPUT86), .B(KEYINPUT24), .ZN(n419) );
  XNOR2_X1 U476 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U477 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U478 ( .A(n424), .B(n423), .Z(n426) );
  NAND2_X1 U479 ( .A1(G228GAT), .A2(G233GAT), .ZN(n425) );
  XNOR2_X1 U480 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U481 ( .A(n428), .B(n427), .Z(n470) );
  NAND2_X1 U482 ( .A1(n455), .A2(n470), .ZN(n429) );
  XNOR2_X1 U483 ( .A(n429), .B(KEYINPUT55), .ZN(n447) );
  XOR2_X1 U484 ( .A(G99GAT), .B(G190GAT), .Z(n432) );
  XNOR2_X1 U485 ( .A(n430), .B(KEYINPUT82), .ZN(n431) );
  XNOR2_X1 U486 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U487 ( .A(n434), .B(n433), .ZN(n436) );
  NAND2_X1 U488 ( .A1(G227GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U489 ( .A(n436), .B(n435), .ZN(n440) );
  XOR2_X1 U490 ( .A(G176GAT), .B(G15GAT), .Z(n438) );
  XNOR2_X1 U491 ( .A(G169GAT), .B(G43GAT), .ZN(n437) );
  XNOR2_X1 U492 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U493 ( .A(n440), .B(n439), .Z(n446) );
  XOR2_X1 U494 ( .A(KEYINPUT83), .B(KEYINPUT80), .Z(n442) );
  XNOR2_X1 U495 ( .A(KEYINPUT20), .B(KEYINPUT79), .ZN(n441) );
  XNOR2_X1 U496 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U497 ( .A(n444), .B(n443), .Z(n445) );
  XOR2_X1 U498 ( .A(n446), .B(n445), .Z(n546) );
  INV_X1 U499 ( .A(n546), .ZN(n535) );
  NAND2_X1 U500 ( .A1(n447), .A2(n535), .ZN(n448) );
  XNOR2_X2 U501 ( .A(KEYINPUT123), .B(n448), .ZN(n578) );
  NAND2_X1 U502 ( .A1(n578), .A2(n569), .ZN(n452) );
  XOR2_X1 U503 ( .A(KEYINPUT126), .B(KEYINPUT58), .Z(n450) );
  INV_X1 U504 ( .A(G190GAT), .ZN(n449) );
  NOR2_X1 U505 ( .A1(n535), .A2(n470), .ZN(n454) );
  XNOR2_X1 U506 ( .A(KEYINPUT26), .B(KEYINPUT93), .ZN(n453) );
  XNOR2_X1 U507 ( .A(n454), .B(n453), .ZN(n468) );
  INV_X1 U508 ( .A(n455), .ZN(n456) );
  NOR2_X1 U509 ( .A1(n468), .A2(n456), .ZN(n589) );
  INV_X1 U510 ( .A(n589), .ZN(n457) );
  NOR2_X1 U511 ( .A1(n489), .A2(n457), .ZN(n458) );
  XNOR2_X1 U512 ( .A(KEYINPUT62), .B(n458), .ZN(n459) );
  XOR2_X1 U513 ( .A(G218GAT), .B(n459), .Z(G1355GAT) );
  XOR2_X1 U514 ( .A(KEYINPUT34), .B(KEYINPUT94), .Z(n478) );
  NAND2_X1 U515 ( .A1(n581), .A2(n460), .ZN(n494) );
  XOR2_X1 U516 ( .A(KEYINPUT16), .B(KEYINPUT77), .Z(n463) );
  NAND2_X1 U517 ( .A1(n461), .A2(n590), .ZN(n462) );
  XNOR2_X1 U518 ( .A(n463), .B(n462), .ZN(n476) );
  XOR2_X1 U519 ( .A(n533), .B(KEYINPUT92), .Z(n464) );
  XNOR2_X1 U520 ( .A(n464), .B(KEYINPUT27), .ZN(n467) );
  XOR2_X1 U521 ( .A(KEYINPUT64), .B(KEYINPUT28), .Z(n465) );
  XOR2_X1 U522 ( .A(n470), .B(n465), .Z(n522) );
  INV_X1 U523 ( .A(n522), .ZN(n538) );
  NOR2_X1 U524 ( .A1(n467), .A2(n538), .ZN(n544) );
  NAND2_X1 U525 ( .A1(n546), .A2(n544), .ZN(n466) );
  INV_X1 U526 ( .A(n543), .ZN(n530) );
  NAND2_X1 U527 ( .A1(n466), .A2(n530), .ZN(n475) );
  NOR2_X1 U528 ( .A1(n468), .A2(n467), .ZN(n560) );
  NAND2_X1 U529 ( .A1(n535), .A2(n533), .ZN(n469) );
  NAND2_X1 U530 ( .A1(n470), .A2(n469), .ZN(n471) );
  XNOR2_X1 U531 ( .A(KEYINPUT25), .B(n471), .ZN(n472) );
  NOR2_X1 U532 ( .A1(n560), .A2(n472), .ZN(n473) );
  NAND2_X1 U533 ( .A1(n473), .A2(n543), .ZN(n474) );
  NAND2_X1 U534 ( .A1(n475), .A2(n474), .ZN(n488) );
  OR2_X1 U535 ( .A1(n476), .A2(n488), .ZN(n510) );
  NOR2_X1 U536 ( .A1(n494), .A2(n510), .ZN(n485) );
  NAND2_X1 U537 ( .A1(n485), .A2(n530), .ZN(n477) );
  XNOR2_X1 U538 ( .A(n478), .B(n477), .ZN(n479) );
  XOR2_X1 U539 ( .A(G1GAT), .B(n479), .Z(G1324GAT) );
  XOR2_X1 U540 ( .A(G8GAT), .B(KEYINPUT95), .Z(n481) );
  NAND2_X1 U541 ( .A1(n485), .A2(n533), .ZN(n480) );
  XNOR2_X1 U542 ( .A(n481), .B(n480), .ZN(G1325GAT) );
  XOR2_X1 U543 ( .A(KEYINPUT35), .B(KEYINPUT96), .Z(n483) );
  NAND2_X1 U544 ( .A1(n485), .A2(n535), .ZN(n482) );
  XNOR2_X1 U545 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U546 ( .A(G15GAT), .B(n484), .ZN(G1326GAT) );
  XOR2_X1 U547 ( .A(G22GAT), .B(KEYINPUT97), .Z(n487) );
  NAND2_X1 U548 ( .A1(n485), .A2(n538), .ZN(n486) );
  XNOR2_X1 U549 ( .A(n487), .B(n486), .ZN(G1327GAT) );
  XOR2_X1 U550 ( .A(KEYINPUT99), .B(KEYINPUT39), .Z(n497) );
  XOR2_X1 U551 ( .A(KEYINPUT98), .B(KEYINPUT37), .Z(n493) );
  NOR2_X1 U552 ( .A1(n489), .A2(n488), .ZN(n491) );
  NAND2_X1 U553 ( .A1(n491), .A2(n490), .ZN(n492) );
  XNOR2_X1 U554 ( .A(n493), .B(n492), .ZN(n527) );
  NOR2_X1 U555 ( .A1(n527), .A2(n494), .ZN(n495) );
  XNOR2_X1 U556 ( .A(n495), .B(KEYINPUT38), .ZN(n505) );
  NAND2_X1 U557 ( .A1(n530), .A2(n505), .ZN(n496) );
  XNOR2_X1 U558 ( .A(n497), .B(n496), .ZN(n498) );
  XOR2_X1 U559 ( .A(G29GAT), .B(n498), .Z(G1328GAT) );
  NAND2_X1 U560 ( .A1(n505), .A2(n533), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n499), .B(KEYINPUT100), .ZN(n500) );
  XNOR2_X1 U562 ( .A(G36GAT), .B(n500), .ZN(G1329GAT) );
  XNOR2_X1 U563 ( .A(G43GAT), .B(KEYINPUT101), .ZN(n504) );
  XOR2_X1 U564 ( .A(KEYINPUT40), .B(KEYINPUT102), .Z(n502) );
  NAND2_X1 U565 ( .A1(n535), .A2(n505), .ZN(n501) );
  XNOR2_X1 U566 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U567 ( .A(n504), .B(n503), .ZN(G1330GAT) );
  XOR2_X1 U568 ( .A(G50GAT), .B(KEYINPUT103), .Z(n507) );
  NAND2_X1 U569 ( .A1(n538), .A2(n505), .ZN(n506) );
  XNOR2_X1 U570 ( .A(n507), .B(n506), .ZN(G1331GAT) );
  NAND2_X1 U571 ( .A1(n573), .A2(n508), .ZN(n509) );
  XOR2_X1 U572 ( .A(KEYINPUT105), .B(n509), .Z(n528) );
  NOR2_X1 U573 ( .A1(n528), .A2(n510), .ZN(n511) );
  XOR2_X1 U574 ( .A(KEYINPUT106), .B(n511), .Z(n521) );
  NOR2_X1 U575 ( .A1(n521), .A2(n543), .ZN(n513) );
  XNOR2_X1 U576 ( .A(KEYINPUT104), .B(KEYINPUT42), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n513), .B(n512), .ZN(n514) );
  XOR2_X1 U578 ( .A(G57GAT), .B(n514), .Z(G1332GAT) );
  XNOR2_X1 U579 ( .A(G64GAT), .B(KEYINPUT107), .ZN(n517) );
  NOR2_X1 U580 ( .A1(n515), .A2(n521), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n517), .B(n516), .ZN(G1333GAT) );
  NOR2_X1 U582 ( .A1(n521), .A2(n546), .ZN(n519) );
  XNOR2_X1 U583 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n518) );
  XNOR2_X1 U584 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U585 ( .A(G71GAT), .B(n520), .ZN(G1334GAT) );
  NOR2_X1 U586 ( .A1(n522), .A2(n521), .ZN(n526) );
  XOR2_X1 U587 ( .A(KEYINPUT111), .B(KEYINPUT43), .Z(n524) );
  XNOR2_X1 U588 ( .A(G78GAT), .B(KEYINPUT110), .ZN(n523) );
  XNOR2_X1 U589 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U590 ( .A(n526), .B(n525), .ZN(G1335GAT) );
  XOR2_X1 U591 ( .A(G85GAT), .B(KEYINPUT113), .Z(n532) );
  NOR2_X1 U592 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U593 ( .A(n529), .B(KEYINPUT112), .ZN(n537) );
  NAND2_X1 U594 ( .A1(n530), .A2(n537), .ZN(n531) );
  XNOR2_X1 U595 ( .A(n532), .B(n531), .ZN(G1336GAT) );
  NAND2_X1 U596 ( .A1(n537), .A2(n533), .ZN(n534) );
  XNOR2_X1 U597 ( .A(n534), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U598 ( .A1(n537), .A2(n535), .ZN(n536) );
  XNOR2_X1 U599 ( .A(n536), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT114), .B(KEYINPUT44), .Z(n540) );
  NAND2_X1 U601 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U602 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U603 ( .A(G106GAT), .B(n541), .Z(G1339GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n548) );
  NOR2_X1 U605 ( .A1(n543), .A2(n542), .ZN(n561) );
  NAND2_X1 U606 ( .A1(n561), .A2(n544), .ZN(n545) );
  NOR2_X1 U607 ( .A1(n546), .A2(n545), .ZN(n555) );
  NAND2_X1 U608 ( .A1(n555), .A2(n581), .ZN(n547) );
  XNOR2_X1 U609 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U610 ( .A(G113GAT), .B(n549), .ZN(G1340GAT) );
  XOR2_X1 U611 ( .A(G120GAT), .B(KEYINPUT49), .Z(n551) );
  NAND2_X1 U612 ( .A1(n555), .A2(n573), .ZN(n550) );
  XNOR2_X1 U613 ( .A(n551), .B(n550), .ZN(G1341GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n553) );
  NAND2_X1 U615 ( .A1(n555), .A2(n590), .ZN(n552) );
  XNOR2_X1 U616 ( .A(n553), .B(n552), .ZN(n554) );
  XOR2_X1 U617 ( .A(G127GAT), .B(n554), .Z(G1342GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT120), .B(KEYINPUT51), .Z(n557) );
  NAND2_X1 U619 ( .A1(n555), .A2(n569), .ZN(n556) );
  XNOR2_X1 U620 ( .A(n557), .B(n556), .ZN(n559) );
  XOR2_X1 U621 ( .A(G134GAT), .B(KEYINPUT119), .Z(n558) );
  XNOR2_X1 U622 ( .A(n559), .B(n558), .ZN(G1343GAT) );
  NAND2_X1 U623 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U624 ( .A(KEYINPUT121), .B(n562), .ZN(n568) );
  NAND2_X1 U625 ( .A1(n581), .A2(n568), .ZN(n563) );
  XNOR2_X1 U626 ( .A(G141GAT), .B(n563), .ZN(G1344GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n565) );
  NAND2_X1 U628 ( .A1(n568), .A2(n573), .ZN(n564) );
  XNOR2_X1 U629 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U630 ( .A(G148GAT), .B(n566), .ZN(G1345GAT) );
  NAND2_X1 U631 ( .A1(n590), .A2(n568), .ZN(n567) );
  XNOR2_X1 U632 ( .A(n567), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U633 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U634 ( .A(n570), .B(KEYINPUT122), .ZN(n571) );
  XNOR2_X1 U635 ( .A(G162GAT), .B(n571), .ZN(G1347GAT) );
  NAND2_X1 U636 ( .A1(n578), .A2(n581), .ZN(n572) );
  XNOR2_X1 U637 ( .A(n572), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U638 ( .A1(n578), .A2(n573), .ZN(n575) );
  XOR2_X1 U639 ( .A(KEYINPUT124), .B(KEYINPUT57), .Z(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n577) );
  XNOR2_X1 U641 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1349GAT) );
  XOR2_X1 U643 ( .A(G183GAT), .B(KEYINPUT125), .Z(n580) );
  NAND2_X1 U644 ( .A1(n578), .A2(n590), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1350GAT) );
  XOR2_X1 U646 ( .A(G197GAT), .B(KEYINPUT59), .Z(n583) );
  NAND2_X1 U647 ( .A1(n589), .A2(n581), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(n585) );
  XOR2_X1 U649 ( .A(KEYINPUT60), .B(KEYINPUT127), .Z(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(G1352GAT) );
  XOR2_X1 U651 ( .A(G204GAT), .B(KEYINPUT61), .Z(n588) );
  NAND2_X1 U652 ( .A1(n589), .A2(n586), .ZN(n587) );
  XNOR2_X1 U653 ( .A(n588), .B(n587), .ZN(G1353GAT) );
  NAND2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U655 ( .A(n591), .B(G211GAT), .ZN(G1354GAT) );
endmodule

