//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 0 0 1 1 0 1 1 0 1 0 1 1 0 1 1 1 1 1 1 0 1 1 0 0 0 0 0 1 1 0 0 0 0 1 1 0 0 0 1 1 0 0 0 0 1 1 0 0 0 1 0 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n624, new_n625, new_n626, new_n628, new_n629, new_n630, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n655, new_n656, new_n657, new_n659, new_n660, new_n661, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n773, new_n775, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n856,
    new_n857, new_n858, new_n859, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n883, new_n884, new_n885, new_n886, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900;
  NOR2_X1   g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(G169gat), .A2(G176gat), .ZN(new_n203));
  AOI21_X1  g002(.A(new_n202), .B1(KEYINPUT23), .B2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G169gat), .ZN(new_n206));
  INV_X1    g005(.A(G176gat), .ZN(new_n207));
  AND2_X1   g006(.A1(new_n207), .A2(KEYINPUT66), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(KEYINPUT66), .ZN(new_n209));
  OAI211_X1 g008(.A(KEYINPUT23), .B(new_n206), .C1(new_n208), .C2(new_n209), .ZN(new_n210));
  OAI21_X1  g009(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  NOR3_X1   g011(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  OAI22_X1  g014(.A1(new_n212), .A2(new_n213), .B1(new_n215), .B2(KEYINPUT24), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT24), .ZN(new_n217));
  OAI21_X1  g016(.A(KEYINPUT64), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT64), .ZN(new_n219));
  NAND4_X1  g018(.A1(new_n219), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n205), .B(new_n210), .C1(new_n216), .C2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT25), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT68), .ZN(new_n225));
  AND3_X1   g024(.A1(new_n214), .A2(new_n225), .A3(new_n217), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n217), .B1(new_n214), .B2(new_n225), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G183gat), .ZN(new_n229));
  INV_X1    g028(.A(G190gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n223), .B1(new_n228), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT67), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n202), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(KEYINPUT67), .B1(G169gat), .B2(G176gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n204), .B1(new_n236), .B2(KEYINPUT23), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n232), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n224), .A2(new_n238), .ZN(new_n239));
  OR2_X1    g038(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n241));
  AOI21_X1  g040(.A(G190gat), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(KEYINPUT28), .B1(new_n242), .B2(KEYINPUT69), .ZN(new_n243));
  INV_X1    g042(.A(new_n241), .ZN(new_n244));
  NOR2_X1   g043(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n230), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT69), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT28), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n246), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n215), .B1(new_n243), .B2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT26), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT70), .B1(new_n236), .B2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT70), .ZN(new_n253));
  AOI211_X1 g052(.A(new_n253), .B(KEYINPUT26), .C1(new_n234), .C2(new_n235), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n202), .B1(new_n251), .B2(new_n203), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n250), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n239), .A2(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(KEYINPUT72), .B(G120gat), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n260), .A2(KEYINPUT73), .A3(G113gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(KEYINPUT74), .B(G113gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(G120gat), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT73), .ZN(new_n264));
  INV_X1    g063(.A(G113gat), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n264), .B1(new_n259), .B2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n261), .A2(new_n263), .A3(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G127gat), .B(G134gat), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT1), .ZN(new_n269));
  AND2_X1   g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n268), .B(KEYINPUT71), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n265), .A2(G120gat), .ZN(new_n273));
  INV_X1    g072(.A(G120gat), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n274), .A2(G113gat), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n269), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n272), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n271), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n258), .B(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(G227gat), .A2(G233gat), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(KEYINPUT32), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT33), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  XOR2_X1   g084(.A(G15gat), .B(G43gat), .Z(new_n286));
  XNOR2_X1  g085(.A(G71gat), .B(G99gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n286), .B(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n283), .B1(new_n285), .B2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT34), .ZN(new_n291));
  OR3_X1    g090(.A1(new_n279), .A2(new_n291), .A3(new_n281), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n291), .B1(new_n279), .B2(new_n281), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT75), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT75), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n292), .A2(new_n296), .A3(new_n293), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n283), .A2(new_n285), .A3(new_n288), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n290), .A2(new_n295), .A3(new_n297), .A4(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n298), .ZN(new_n300));
  OAI211_X1 g099(.A(KEYINPUT75), .B(new_n294), .C1(new_n300), .C2(new_n289), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(KEYINPUT76), .A2(KEYINPUT36), .ZN(new_n303));
  OR2_X1    g102(.A1(KEYINPUT76), .A2(KEYINPUT36), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n299), .A2(new_n301), .A3(KEYINPUT76), .A4(KEYINPUT36), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G22gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(G228gat), .A2(G233gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(G155gat), .A2(G162gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n310), .B(KEYINPUT83), .ZN(new_n311));
  OR2_X1    g110(.A1(G155gat), .A2(G162gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(G141gat), .B(G148gat), .ZN(new_n313));
  AND2_X1   g112(.A1(KEYINPUT83), .A2(KEYINPUT2), .ZN(new_n314));
  OAI211_X1 g113(.A(new_n311), .B(new_n312), .C1(new_n313), .C2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(G141gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(G148gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(KEYINPUT84), .B(G148gat), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n317), .B1(new_n318), .B2(new_n316), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n310), .B1(new_n312), .B2(KEYINPUT2), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n315), .A2(new_n321), .ZN(new_n322));
  XOR2_X1   g121(.A(KEYINPUT77), .B(G204gat), .Z(new_n323));
  INV_X1    g122(.A(G197gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AND2_X1   g124(.A1(G211gat), .A2(G218gat), .ZN(new_n326));
  OR2_X1    g125(.A1(new_n326), .A2(KEYINPUT22), .ZN(new_n327));
  XNOR2_X1  g126(.A(KEYINPUT77), .B(G204gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(G197gat), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n325), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  XOR2_X1   g129(.A(G211gat), .B(G218gat), .Z(new_n331));
  NAND3_X1  g130(.A1(new_n330), .A2(KEYINPUT78), .A3(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n328), .B(new_n324), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n331), .A2(KEYINPUT78), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n333), .A2(new_n334), .A3(new_n327), .ZN(new_n335));
  AOI21_X1  g134(.A(KEYINPUT29), .B1(new_n332), .B2(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n322), .B1(new_n336), .B2(KEYINPUT3), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT90), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n309), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  AND3_X1   g138(.A1(new_n332), .A2(KEYINPUT79), .A3(new_n335), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT79), .B1(new_n332), .B2(new_n335), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AND2_X1   g141(.A1(new_n315), .A2(new_n321), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT3), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT29), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n342), .A2(new_n347), .ZN(new_n348));
  OAI211_X1 g147(.A(new_n339), .B(new_n348), .C1(new_n338), .C2(new_n337), .ZN(new_n349));
  INV_X1    g148(.A(new_n331), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n346), .B1(new_n330), .B2(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n331), .B1(new_n333), .B2(new_n327), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n344), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  AND3_X1   g152(.A1(new_n315), .A2(new_n321), .A3(KEYINPUT85), .ZN(new_n354));
  AOI21_X1  g153(.A(KEYINPUT85), .B1(new_n315), .B2(new_n321), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n348), .A2(new_n357), .ZN(new_n358));
  XOR2_X1   g157(.A(new_n309), .B(KEYINPUT89), .Z(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n308), .B1(new_n349), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n349), .A2(new_n360), .A3(new_n308), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n362), .A2(KEYINPUT91), .A3(new_n363), .ZN(new_n364));
  XNOR2_X1  g163(.A(KEYINPUT88), .B(KEYINPUT31), .ZN(new_n365));
  INV_X1    g164(.A(G50gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n365), .B(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(G78gat), .B(G106gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n367), .B(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  OR2_X1    g169(.A1(new_n364), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT91), .ZN(new_n372));
  INV_X1    g171(.A(new_n363), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n372), .B1(new_n373), .B2(new_n361), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n364), .A2(new_n374), .A3(new_n370), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n371), .A2(new_n375), .ZN(new_n376));
  NOR3_X1   g175(.A1(new_n242), .A2(KEYINPUT69), .A3(KEYINPUT28), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n248), .B1(new_n246), .B2(new_n247), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n214), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n235), .ZN(new_n380));
  NOR3_X1   g179(.A1(KEYINPUT67), .A2(G169gat), .A3(G176gat), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n251), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(new_n253), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n236), .A2(KEYINPUT70), .A3(new_n251), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n256), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n379), .A2(new_n385), .ZN(new_n386));
  AOI22_X1  g185(.A1(new_n223), .A2(new_n222), .B1(new_n232), .B2(new_n237), .ZN(new_n387));
  OAI21_X1  g186(.A(KEYINPUT80), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(G226gat), .A2(G233gat), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT80), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n239), .A2(new_n257), .A3(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n388), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n258), .A2(new_n346), .A3(new_n389), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n342), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT81), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n388), .A2(new_n392), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n400), .A2(new_n346), .A3(new_n389), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n239), .A2(new_n257), .A3(new_n390), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n401), .A2(new_n342), .A3(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n395), .A2(KEYINPUT81), .A3(new_n396), .ZN(new_n404));
  XNOR2_X1  g203(.A(G8gat), .B(G36gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n405), .B(G64gat), .ZN(new_n406));
  INV_X1    g205(.A(G92gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n406), .B(new_n407), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n399), .A2(new_n403), .A3(new_n404), .A4(new_n408), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n409), .A2(KEYINPUT30), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT30), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n399), .A2(new_n403), .A3(new_n404), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n408), .B(KEYINPUT82), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n411), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n410), .B1(new_n409), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT39), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n278), .A2(new_n322), .ZN(new_n417));
  AOI22_X1  g216(.A1(new_n267), .A2(new_n270), .B1(new_n276), .B2(new_n272), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n418), .A2(new_n343), .ZN(new_n419));
  NAND2_X1  g218(.A1(G225gat), .A2(G233gat), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  OR3_X1    g220(.A1(new_n417), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n416), .B1(new_n422), .B2(KEYINPUT92), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n322), .A2(KEYINPUT3), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n278), .A2(new_n345), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(KEYINPUT4), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n418), .B1(new_n355), .B2(new_n354), .ZN(new_n427));
  AOI22_X1  g226(.A1(new_n426), .A2(new_n427), .B1(KEYINPUT4), .B2(new_n417), .ZN(new_n428));
  OAI221_X1 g227(.A(new_n423), .B1(KEYINPUT92), .B2(new_n422), .C1(new_n420), .C2(new_n428), .ZN(new_n429));
  XOR2_X1   g228(.A(G1gat), .B(G29gat), .Z(new_n430));
  XNOR2_X1  g229(.A(G57gat), .B(G85gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n430), .B(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(KEYINPUT86), .B(KEYINPUT0), .ZN(new_n433));
  XOR2_X1   g232(.A(new_n432), .B(new_n433), .Z(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  OR3_X1    g234(.A1(new_n428), .A2(KEYINPUT39), .A3(new_n420), .ZN(new_n436));
  AND4_X1   g235(.A1(KEYINPUT40), .A2(new_n429), .A3(new_n435), .A4(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n421), .B1(new_n417), .B2(new_n419), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n417), .B1(KEYINPUT4), .B2(new_n425), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT4), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n420), .B1(new_n427), .B2(new_n440), .ZN(new_n441));
  OAI211_X1 g240(.A(KEYINPUT5), .B(new_n438), .C1(new_n439), .C2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n417), .A2(KEYINPUT4), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n421), .A2(KEYINPUT5), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n435), .B1(new_n442), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(KEYINPUT40), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n429), .A2(new_n436), .A3(new_n435), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n437), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n376), .B1(new_n415), .B2(new_n451), .ZN(new_n452));
  OR2_X1    g251(.A1(new_n412), .A2(KEYINPUT37), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n408), .B1(new_n412), .B2(KEYINPUT37), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n453), .B1(new_n454), .B2(KEYINPUT94), .ZN(new_n455));
  AND2_X1   g254(.A1(new_n454), .A2(KEYINPUT94), .ZN(new_n456));
  OAI21_X1  g255(.A(KEYINPUT38), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n442), .A2(new_n446), .A3(new_n435), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT6), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n460), .B(new_n447), .ZN(new_n461));
  INV_X1    g260(.A(new_n413), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n393), .A2(new_n342), .A3(new_n394), .ZN(new_n463));
  OR2_X1    g262(.A1(new_n463), .A2(KEYINPUT93), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(KEYINPUT93), .ZN(new_n465));
  AND2_X1   g264(.A1(new_n401), .A2(new_n402), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n464), .B(new_n465), .C1(new_n342), .C2(new_n466), .ZN(new_n467));
  AOI211_X1 g266(.A(KEYINPUT38), .B(new_n462), .C1(new_n467), .C2(KEYINPUT37), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n461), .B1(new_n468), .B2(new_n453), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n457), .A2(new_n469), .A3(new_n409), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n307), .B1(new_n452), .B2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT87), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n460), .B(new_n448), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n472), .B1(new_n415), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n412), .A2(new_n413), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n475), .A2(KEYINPUT30), .A3(new_n409), .ZN(new_n476));
  OR2_X1    g275(.A1(new_n409), .A2(KEYINPUT30), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n478), .A2(KEYINPUT87), .A3(new_n461), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n474), .A2(new_n479), .A3(new_n376), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n471), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n302), .A2(new_n371), .A3(new_n375), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT35), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n483), .A2(new_n484), .A3(new_n461), .A4(new_n478), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n482), .B1(new_n474), .B2(new_n479), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n485), .B1(new_n486), .B2(new_n484), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n481), .A2(new_n487), .ZN(new_n488));
  XNOR2_X1  g287(.A(G15gat), .B(G22gat), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT16), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n489), .B1(new_n490), .B2(G1gat), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n491), .B1(G1gat), .B2(new_n489), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n492), .B(G8gat), .ZN(new_n493));
  XOR2_X1   g292(.A(G43gat), .B(G50gat), .Z(new_n494));
  INV_X1    g293(.A(KEYINPUT15), .ZN(new_n495));
  OR2_X1    g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n494), .A2(new_n495), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT14), .ZN(new_n498));
  INV_X1    g297(.A(G29gat), .ZN(new_n499));
  INV_X1    g298(.A(G36gat), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n502));
  AOI22_X1  g301(.A1(new_n501), .A2(new_n502), .B1(G29gat), .B2(G36gat), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n496), .A2(new_n497), .A3(new_n503), .ZN(new_n504));
  OR3_X1    g303(.A1(new_n503), .A2(new_n495), .A3(new_n494), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT96), .B1(new_n493), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT17), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n504), .A2(KEYINPUT17), .A3(new_n505), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n507), .B1(new_n511), .B2(new_n493), .ZN(new_n512));
  INV_X1    g311(.A(new_n493), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n513), .A2(KEYINPUT96), .A3(new_n510), .A4(new_n509), .ZN(new_n514));
  AOI22_X1  g313(.A1(new_n512), .A2(new_n514), .B1(G229gat), .B2(G233gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(KEYINPUT18), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT97), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT97), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n515), .A2(new_n518), .A3(KEYINPUT18), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n515), .A2(KEYINPUT18), .ZN(new_n521));
  XOR2_X1   g320(.A(new_n493), .B(new_n506), .Z(new_n522));
  NAND2_X1  g321(.A1(G229gat), .A2(G233gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n523), .B(KEYINPUT13), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n521), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n520), .A2(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(G113gat), .B(G141gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(G169gat), .B(G197gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(KEYINPUT95), .B(KEYINPUT11), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  XOR2_X1   g331(.A(new_n532), .B(KEYINPUT12), .Z(new_n533));
  OAI21_X1  g332(.A(new_n533), .B1(new_n521), .B2(KEYINPUT98), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n527), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n534), .B1(new_n520), .B2(new_n526), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(G230gat), .A2(G233gat), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(G99gat), .A2(G106gat), .ZN(new_n541));
  INV_X1    g340(.A(G85gat), .ZN(new_n542));
  AOI22_X1  g341(.A1(KEYINPUT8), .A2(new_n541), .B1(new_n542), .B2(new_n407), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(KEYINPUT104), .ZN(new_n544));
  NAND2_X1  g343(.A1(G85gat), .A2(G92gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(KEYINPUT7), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  XOR2_X1   g346(.A(G99gat), .B(G106gat), .Z(new_n548));
  OR2_X1    g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(new_n548), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT99), .ZN(new_n552));
  XNOR2_X1  g351(.A(G57gat), .B(G64gat), .ZN(new_n553));
  AND2_X1   g352(.A1(G71gat), .A2(G78gat), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n554), .A2(KEYINPUT9), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n552), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g355(.A1(G71gat), .A2(G78gat), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  XOR2_X1   g357(.A(new_n556), .B(new_n558), .Z(new_n559));
  NAND2_X1  g358(.A1(new_n551), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT10), .ZN(new_n561));
  INV_X1    g360(.A(new_n559), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n562), .A2(new_n549), .A3(new_n550), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n560), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  OR2_X1    g363(.A1(new_n563), .A2(new_n561), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n540), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n539), .B1(new_n560), .B2(new_n563), .ZN(new_n567));
  OR2_X1    g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G120gat), .B(G148gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(new_n207), .ZN(new_n570));
  XOR2_X1   g369(.A(new_n570), .B(G204gat), .Z(new_n571));
  XNOR2_X1  g370(.A(new_n568), .B(new_n571), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n538), .A2(new_n572), .ZN(new_n573));
  AND2_X1   g372(.A1(new_n488), .A2(new_n573), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n562), .A2(KEYINPUT21), .ZN(new_n575));
  XOR2_X1   g374(.A(G183gat), .B(G211gat), .Z(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(G127gat), .B(G155gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(KEYINPUT20), .ZN(new_n579));
  XOR2_X1   g378(.A(new_n577), .B(new_n579), .Z(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n493), .B1(new_n562), .B2(KEYINPUT21), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT103), .ZN(new_n583));
  XOR2_X1   g382(.A(KEYINPUT100), .B(KEYINPUT101), .Z(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(KEYINPUT102), .B(KEYINPUT19), .ZN(new_n586));
  OR2_X1    g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(G231gat), .ZN(new_n588));
  INV_X1    g387(.A(G233gat), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n585), .A2(new_n586), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n587), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n591), .B1(new_n587), .B2(new_n592), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n581), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n595), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n597), .A2(new_n593), .A3(new_n580), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n549), .A2(new_n550), .A3(new_n506), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT41), .ZN(new_n602));
  NAND2_X1  g401(.A1(G232gat), .A2(G233gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n551), .B(KEYINPUT105), .ZN(new_n604));
  OAI221_X1 g403(.A(new_n601), .B1(new_n602), .B2(new_n603), .C1(new_n604), .C2(new_n511), .ZN(new_n605));
  XNOR2_X1  g404(.A(G134gat), .B(G162gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  XOR2_X1   g406(.A(G190gat), .B(G218gat), .Z(new_n608));
  NAND2_X1  g407(.A1(new_n603), .A2(new_n602), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n607), .B(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n574), .A2(new_n600), .A3(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(new_n473), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g414(.A1(new_n612), .A2(new_n478), .ZN(new_n616));
  INV_X1    g415(.A(G8gat), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n490), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n619), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n620));
  OR2_X1    g419(.A1(new_n620), .A2(KEYINPUT42), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(KEYINPUT42), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n621), .B(new_n622), .C1(new_n617), .C2(new_n616), .ZN(G1325gat));
  AOI21_X1  g422(.A(G15gat), .B1(new_n613), .B2(new_n302), .ZN(new_n624));
  INV_X1    g423(.A(new_n307), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n612), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n624), .B1(G15gat), .B2(new_n626), .ZN(G1326gat));
  INV_X1    g426(.A(new_n376), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n612), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g428(.A(KEYINPUT43), .B(G22gat), .Z(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(G1327gat));
  INV_X1    g430(.A(KEYINPUT106), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n480), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n474), .A2(new_n479), .A3(KEYINPUT106), .A4(new_n376), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AND3_X1   g434(.A1(new_n635), .A2(KEYINPUT107), .A3(new_n471), .ZN(new_n636));
  AOI21_X1  g435(.A(KEYINPUT107), .B1(new_n635), .B2(new_n471), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n487), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT44), .ZN(new_n639));
  INV_X1    g438(.A(new_n611), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT108), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n488), .A2(new_n640), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n642), .B1(new_n643), .B2(KEYINPUT44), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n638), .A2(new_n642), .A3(new_n639), .A4(new_n640), .ZN(new_n646));
  AND2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n599), .A2(new_n573), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g448(.A(G29gat), .B1(new_n649), .B2(new_n461), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n488), .A2(new_n640), .A3(new_n648), .ZN(new_n651));
  NOR3_X1   g450(.A1(new_n651), .A2(G29gat), .A3(new_n461), .ZN(new_n652));
  XOR2_X1   g451(.A(new_n652), .B(KEYINPUT45), .Z(new_n653));
  NAND2_X1  g452(.A1(new_n650), .A2(new_n653), .ZN(G1328gat));
  OAI21_X1  g453(.A(G36gat), .B1(new_n649), .B2(new_n478), .ZN(new_n655));
  NOR3_X1   g454(.A1(new_n651), .A2(G36gat), .A3(new_n478), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(KEYINPUT46), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n655), .A2(new_n657), .ZN(G1329gat));
  NAND2_X1  g457(.A1(new_n307), .A2(G43gat), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n651), .B1(new_n301), .B2(new_n299), .ZN(new_n660));
  OAI22_X1  g459(.A1(new_n649), .A2(new_n659), .B1(G43gat), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g461(.A(new_n366), .B1(new_n651), .B2(new_n628), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n376), .A2(G50gat), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n663), .B1(new_n649), .B2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT48), .ZN(G1331gat));
  NAND3_X1  g465(.A1(new_n596), .A2(new_n598), .A3(new_n611), .ZN(new_n667));
  INV_X1    g466(.A(new_n538), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n635), .A2(new_n471), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT107), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n635), .A2(KEYINPUT107), .A3(new_n471), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AOI211_X1 g472(.A(new_n667), .B(new_n668), .C1(new_n673), .C2(new_n487), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n674), .A2(new_n572), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(new_n473), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g476(.A1(new_n674), .A2(new_n572), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n415), .B(KEYINPUT109), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n682));
  AND2_X1   g481(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n681), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n684), .B1(new_n681), .B2(new_n682), .ZN(G1333gat));
  INV_X1    g484(.A(G71gat), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n302), .B(KEYINPUT110), .Z(new_n687));
  NAND3_X1  g486(.A1(new_n675), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(G71gat), .B1(new_n678), .B2(new_n625), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XOR2_X1   g489(.A(new_n690), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g490(.A1(new_n678), .A2(new_n628), .ZN(new_n692));
  XOR2_X1   g491(.A(KEYINPUT111), .B(G78gat), .Z(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT112), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n692), .B(new_n694), .ZN(G1335gat));
  NAND2_X1  g494(.A1(new_n599), .A2(new_n538), .ZN(new_n696));
  INV_X1    g495(.A(new_n572), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n647), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(G85gat), .B1(new_n699), .B2(new_n461), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n611), .B1(new_n673), .B2(new_n487), .ZN(new_n701));
  INV_X1    g500(.A(new_n696), .ZN(new_n702));
  AOI21_X1  g501(.A(KEYINPUT51), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  AND4_X1   g502(.A1(KEYINPUT51), .A2(new_n638), .A3(new_n640), .A4(new_n702), .ZN(new_n704));
  OR3_X1    g503(.A1(new_n703), .A2(new_n704), .A3(KEYINPUT113), .ZN(new_n705));
  OAI21_X1  g504(.A(KEYINPUT113), .B1(new_n703), .B2(new_n704), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n473), .A2(new_n542), .A3(new_n572), .ZN(new_n707));
  XOR2_X1   g506(.A(new_n707), .B(KEYINPUT114), .Z(new_n708));
  NAND3_X1  g507(.A1(new_n705), .A2(new_n706), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n700), .A2(new_n709), .ZN(G1336gat));
  OAI21_X1  g509(.A(G92gat), .B1(new_n699), .B2(new_n680), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT52), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n680), .A2(G92gat), .A3(new_n697), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n713), .B1(new_n703), .B2(new_n704), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n711), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n645), .A2(new_n415), .A3(new_n646), .A4(new_n698), .ZN(new_n716));
  AND3_X1   g515(.A1(new_n716), .A2(KEYINPUT115), .A3(G92gat), .ZN(new_n717));
  AOI21_X1  g516(.A(KEYINPUT115), .B1(new_n716), .B2(G92gat), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n703), .A2(new_n704), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n713), .B(KEYINPUT116), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n717), .A2(new_n718), .A3(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n715), .B1(new_n722), .B2(new_n712), .ZN(G1337gat));
  OAI21_X1  g522(.A(G99gat), .B1(new_n699), .B2(new_n625), .ZN(new_n724));
  INV_X1    g523(.A(G99gat), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n705), .A2(new_n725), .A3(new_n302), .A4(new_n706), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n724), .B1(new_n726), .B2(new_n697), .ZN(G1338gat));
  INV_X1    g526(.A(KEYINPUT53), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n645), .A2(new_n376), .A3(new_n646), .A4(new_n698), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(G106gat), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT117), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n628), .A2(G106gat), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n572), .B(new_n732), .C1(new_n703), .C2(new_n704), .ZN(new_n733));
  AND3_X1   g532(.A1(new_n730), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n731), .B1(new_n730), .B2(new_n733), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n728), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n730), .A2(new_n733), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(KEYINPUT117), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n730), .A2(new_n731), .A3(new_n733), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n738), .A2(KEYINPUT53), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n736), .A2(new_n740), .ZN(G1339gat));
  NAND2_X1  g540(.A1(new_n522), .A2(new_n524), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n512), .A2(new_n514), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n742), .B1(new_n743), .B2(new_n523), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n532), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n572), .B(new_n745), .C1(new_n533), .C2(new_n527), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n568), .A2(new_n571), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n564), .A2(new_n565), .A3(new_n540), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(KEYINPUT54), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n749), .A2(new_n566), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n564), .A2(new_n565), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT54), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n751), .A2(new_n752), .A3(new_n539), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n571), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n750), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n747), .B1(new_n755), .B2(KEYINPUT55), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n756), .B1(KEYINPUT55), .B2(new_n755), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n746), .B1(new_n757), .B2(new_n538), .ZN(new_n758));
  AND2_X1   g557(.A1(new_n758), .A2(new_n611), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n745), .B1(new_n527), .B2(new_n533), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n611), .A2(new_n757), .A3(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n599), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n600), .A2(new_n611), .A3(new_n697), .A4(new_n538), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(KEYINPUT118), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT118), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n762), .A2(new_n763), .A3(new_n766), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n768), .A2(new_n473), .A3(new_n628), .A4(new_n302), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n769), .A2(new_n679), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n668), .ZN(new_n771));
  MUX2_X1   g570(.A(new_n262), .B(G113gat), .S(new_n771), .Z(G1340gat));
  NAND2_X1  g571(.A1(new_n770), .A2(new_n572), .ZN(new_n773));
  MUX2_X1   g572(.A(new_n260), .B(G120gat), .S(new_n773), .Z(G1341gat));
  NAND2_X1  g573(.A1(new_n770), .A2(new_n600), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(G127gat), .ZN(G1342gat));
  INV_X1    g575(.A(new_n770), .ZN(new_n777));
  OAI21_X1  g576(.A(G134gat), .B1(new_n777), .B2(new_n611), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n611), .A2(new_n415), .ZN(new_n779));
  INV_X1    g578(.A(G134gat), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(KEYINPUT56), .B1(new_n769), .B2(new_n781), .ZN(new_n782));
  OR3_X1    g581(.A1(new_n769), .A2(KEYINPUT56), .A3(new_n781), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n778), .A2(new_n782), .A3(new_n783), .ZN(G1343gat));
  AND2_X1   g583(.A1(new_n768), .A2(new_n376), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n307), .A2(new_n461), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(new_n680), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n785), .A2(new_n316), .A3(new_n668), .A4(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT57), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n765), .A2(new_n790), .A3(new_n376), .A4(new_n767), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(new_n788), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT119), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n793), .B1(new_n750), .B2(new_n754), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT55), .ZN(new_n795));
  INV_X1    g594(.A(new_n571), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n796), .B1(new_n566), .B2(new_n752), .ZN(new_n797));
  OAI211_X1 g596(.A(new_n797), .B(KEYINPUT119), .C1(new_n566), .C2(new_n749), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n794), .A2(new_n795), .A3(new_n798), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n799), .B(new_n756), .C1(new_n536), .C2(new_n537), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT120), .ZN(new_n801));
  AND3_X1   g600(.A1(new_n800), .A2(new_n801), .A3(new_n746), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n801), .B1(new_n800), .B2(new_n746), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n802), .A2(new_n803), .A3(new_n640), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n599), .B1(new_n804), .B2(new_n761), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(new_n763), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n790), .B1(new_n806), .B2(new_n376), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n792), .A2(new_n538), .A3(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n789), .B1(new_n316), .B2(new_n808), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(KEYINPUT58), .ZN(G1344gat));
  NOR2_X1   g609(.A1(new_n792), .A2(new_n807), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n572), .ZN(new_n812));
  AOI21_X1  g611(.A(KEYINPUT59), .B1(new_n812), .B2(new_n318), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n785), .A2(new_n788), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n814), .A2(new_n318), .A3(new_n697), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n805), .A2(KEYINPUT121), .A3(new_n763), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT121), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n800), .A2(new_n746), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(KEYINPUT120), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n800), .A2(new_n801), .A3(new_n746), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n820), .A2(new_n611), .A3(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(new_n761), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n600), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n667), .A2(new_n572), .A3(new_n668), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n818), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n817), .A2(new_n826), .A3(new_n376), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n790), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(KEYINPUT122), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n768), .A2(KEYINPUT57), .A3(new_n376), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT122), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n827), .A2(new_n831), .A3(new_n790), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n829), .A2(new_n830), .A3(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n833), .A2(new_n572), .A3(new_n788), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n834), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n816), .A2(new_n835), .ZN(G1345gat));
  NOR2_X1   g635(.A1(new_n814), .A2(new_n599), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n837), .A2(G155gat), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n811), .A2(G155gat), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n838), .B1(new_n839), .B2(new_n600), .ZN(G1346gat));
  INV_X1    g639(.A(G162gat), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n785), .A2(new_n841), .A3(new_n779), .A4(new_n786), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n792), .A2(new_n611), .A3(new_n807), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n842), .B1(new_n843), .B2(new_n841), .ZN(G1347gat));
  AND4_X1   g643(.A1(new_n461), .A2(new_n765), .A3(new_n679), .A4(new_n767), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n483), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n847), .A2(new_n206), .A3(new_n668), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n765), .A2(new_n628), .A3(new_n687), .A4(new_n767), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n478), .A2(new_n473), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(G169gat), .B1(new_n853), .B2(new_n538), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n848), .A2(new_n854), .ZN(G1348gat));
  NOR4_X1   g654(.A1(new_n853), .A2(new_n697), .A3(new_n208), .A4(new_n209), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n207), .B1(new_n846), .B2(new_n697), .ZN(new_n857));
  OR2_X1    g656(.A1(new_n857), .A2(KEYINPUT123), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(KEYINPUT123), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n856), .B1(new_n858), .B2(new_n859), .ZN(G1349gat));
  INV_X1    g659(.A(KEYINPUT124), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n861), .B1(new_n852), .B2(new_n600), .ZN(new_n862));
  NOR4_X1   g661(.A1(new_n849), .A2(KEYINPUT124), .A3(new_n599), .A4(new_n851), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n862), .A2(new_n229), .A3(new_n863), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n244), .A2(new_n245), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n846), .A2(new_n599), .A3(new_n865), .ZN(new_n866));
  OR3_X1    g665(.A1(new_n864), .A2(KEYINPUT60), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(KEYINPUT60), .B1(new_n864), .B2(new_n866), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(G1350gat));
  AOI21_X1  g668(.A(new_n230), .B1(new_n852), .B2(new_n640), .ZN(new_n870));
  XOR2_X1   g669(.A(new_n870), .B(KEYINPUT61), .Z(new_n871));
  NAND3_X1  g670(.A1(new_n847), .A2(new_n230), .A3(new_n640), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(G1351gat));
  NOR2_X1   g672(.A1(new_n307), .A2(new_n628), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n845), .A2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(G197gat), .B1(new_n876), .B2(new_n668), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n307), .A2(new_n851), .ZN(new_n878));
  XOR2_X1   g677(.A(new_n878), .B(KEYINPUT125), .Z(new_n879));
  AND2_X1   g678(.A1(new_n833), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n538), .A2(new_n324), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n877), .B1(new_n880), .B2(new_n881), .ZN(G1352gat));
  NOR3_X1   g681(.A1(new_n875), .A2(G204gat), .A3(new_n697), .ZN(new_n883));
  XNOR2_X1  g682(.A(new_n883), .B(KEYINPUT62), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n833), .A2(new_n572), .A3(new_n879), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(G204gat), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n884), .A2(new_n886), .ZN(G1353gat));
  NAND3_X1  g686(.A1(new_n833), .A2(new_n600), .A3(new_n878), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT63), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(KEYINPUT126), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n888), .A2(G211gat), .A3(new_n890), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n889), .A2(KEYINPUT126), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OR3_X1    g692(.A1(new_n875), .A2(G211gat), .A3(new_n599), .ZN(new_n894));
  INV_X1    g693(.A(new_n892), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n888), .A2(G211gat), .A3(new_n895), .A4(new_n890), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n893), .A2(new_n894), .A3(new_n896), .ZN(G1354gat));
  AOI21_X1  g696(.A(G218gat), .B1(new_n876), .B2(new_n640), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n640), .A2(G218gat), .ZN(new_n899));
  XOR2_X1   g698(.A(new_n899), .B(KEYINPUT127), .Z(new_n900));
  AOI21_X1  g699(.A(new_n898), .B1(new_n880), .B2(new_n900), .ZN(G1355gat));
endmodule


