//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 1 1 1 1 0 1 1 0 1 0 0 1 1 0 1 0 1 1 0 1 0 1 1 0 0 1 0 0 1 0 1 1 0 0 0 1 1 0 1 0 1 0 0 1 1 1 1 0 0 1 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:35 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n734, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  NOR2_X1   g001(.A1(G237), .A2(G953), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G210), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(G101), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n190), .B(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT11), .ZN(new_n193));
  INV_X1    g007(.A(G134), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n193), .B1(new_n194), .B2(G137), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(G137), .ZN(new_n196));
  INV_X1    g010(.A(G137), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(KEYINPUT11), .A3(G134), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n195), .A2(new_n196), .A3(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n199), .A2(KEYINPUT64), .A3(G131), .ZN(new_n200));
  NAND2_X1  g014(.A1(KEYINPUT64), .A2(G131), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n195), .A2(new_n198), .A3(new_n201), .A4(new_n196), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G146), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G143), .ZN(new_n205));
  INV_X1    g019(.A(G143), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT0), .ZN(new_n209));
  INV_X1    g023(.A(G128), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(KEYINPUT0), .A2(G128), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n208), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  OAI211_X1 g027(.A(new_n205), .B(new_n207), .C1(new_n209), .C2(new_n210), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n203), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT2), .ZN(new_n217));
  INV_X1    g031(.A(G113), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(new_n218), .A3(KEYINPUT66), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT66), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n220), .B1(KEYINPUT2), .B2(G113), .ZN(new_n221));
  AOI22_X1  g035(.A1(new_n219), .A2(new_n221), .B1(KEYINPUT2), .B2(G113), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G116), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n224), .A2(G119), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT67), .ZN(new_n226));
  INV_X1    g040(.A(G119), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n226), .B1(new_n227), .B2(G116), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n224), .A2(KEYINPUT67), .A3(G119), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n225), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n230), .A2(KEYINPUT68), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT68), .ZN(new_n232));
  AOI211_X1 g046(.A(new_n232), .B(new_n225), .C1(new_n228), .C2(new_n229), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n223), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n222), .A2(new_n230), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n197), .A2(G134), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n194), .A2(G137), .ZN(new_n237));
  OAI21_X1  g051(.A(G131), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT65), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n210), .A2(KEYINPUT1), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n241), .A2(new_n205), .A3(new_n207), .ZN(new_n242));
  OAI211_X1 g056(.A(new_n206), .B(G146), .C1(new_n210), .C2(KEYINPUT1), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n210), .A2(new_n204), .A3(G143), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n242), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(G131), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n195), .A2(new_n198), .A3(new_n246), .A4(new_n196), .ZN(new_n247));
  OAI211_X1 g061(.A(KEYINPUT65), .B(G131), .C1(new_n236), .C2(new_n237), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n240), .A2(new_n245), .A3(new_n247), .A4(new_n248), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n216), .A2(new_n234), .A3(new_n235), .A4(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  AOI22_X1  g065(.A1(new_n216), .A2(new_n249), .B1(new_n234), .B2(new_n235), .ZN(new_n252));
  OAI21_X1  g066(.A(KEYINPUT28), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT28), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n250), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n192), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n234), .A2(new_n235), .ZN(new_n257));
  AND4_X1   g071(.A1(new_n247), .A2(new_n240), .A3(new_n245), .A4(new_n248), .ZN(new_n258));
  AOI22_X1  g072(.A1(new_n200), .A2(new_n202), .B1(new_n213), .B2(new_n214), .ZN(new_n259));
  NOR3_X1   g073(.A1(new_n258), .A2(KEYINPUT30), .A3(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT30), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n261), .B1(new_n216), .B2(new_n249), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n257), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n263), .A2(new_n250), .A3(new_n192), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT31), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(KEYINPUT30), .B1(new_n258), .B2(new_n259), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n216), .A2(new_n261), .A3(new_n249), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n251), .B1(new_n269), .B2(new_n257), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n270), .A2(KEYINPUT31), .A3(new_n192), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n256), .B1(new_n266), .B2(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(G472), .A2(G902), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n187), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n192), .ZN(new_n276));
  INV_X1    g090(.A(new_n252), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n254), .B1(new_n277), .B2(new_n250), .ZN(new_n278));
  INV_X1    g092(.A(new_n255), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n276), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(KEYINPUT31), .B1(new_n270), .B2(new_n192), .ZN(new_n281));
  AND4_X1   g095(.A1(KEYINPUT31), .A2(new_n263), .A3(new_n250), .A4(new_n192), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n283), .A2(KEYINPUT32), .A3(new_n273), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n275), .A2(new_n284), .A3(KEYINPUT69), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n283), .A2(new_n273), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT69), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n286), .A2(new_n287), .A3(new_n187), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(G472), .ZN(new_n290));
  OR2_X1    g104(.A1(new_n255), .A2(KEYINPUT70), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n255), .A2(KEYINPUT70), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n278), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT29), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n276), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(G902), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n270), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n276), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n253), .A2(new_n255), .A3(new_n192), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n298), .A2(new_n294), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n290), .B1(new_n296), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n289), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(KEYINPUT23), .B1(new_n210), .B2(G119), .ZN(new_n304));
  OAI21_X1  g118(.A(KEYINPUT72), .B1(new_n227), .B2(G128), .ZN(new_n305));
  XNOR2_X1  g119(.A(new_n304), .B(new_n305), .ZN(new_n306));
  XOR2_X1   g120(.A(KEYINPUT73), .B(G110), .Z(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  XOR2_X1   g122(.A(G119), .B(G128), .Z(new_n309));
  XNOR2_X1  g123(.A(KEYINPUT24), .B(G110), .ZN(new_n310));
  AOI21_X1  g124(.A(KEYINPUT74), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(new_n310), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT74), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n308), .B1(new_n311), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT75), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n308), .B(KEYINPUT75), .C1(new_n311), .C2(new_n314), .ZN(new_n318));
  OR2_X1    g132(.A1(G125), .A2(G140), .ZN(new_n319));
  NAND2_X1  g133(.A1(G125), .A2(G140), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(new_n204), .ZN(new_n322));
  AND2_X1   g136(.A1(G125), .A2(G140), .ZN(new_n323));
  NOR2_X1   g137(.A1(G125), .A2(G140), .ZN(new_n324));
  OAI21_X1  g138(.A(KEYINPUT16), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G125), .ZN(new_n326));
  OR3_X1    g140(.A1(new_n326), .A2(KEYINPUT16), .A3(G140), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n325), .A2(new_n327), .A3(G146), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n328), .B(KEYINPUT76), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n317), .A2(new_n318), .A3(new_n322), .A4(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(G110), .ZN(new_n331));
  OR2_X1    g145(.A1(new_n306), .A2(new_n331), .ZN(new_n332));
  OR2_X1    g146(.A1(new_n309), .A2(new_n310), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT71), .ZN(new_n334));
  OR2_X1    g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n325), .A2(new_n327), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n204), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n328), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n333), .A2(new_n334), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n332), .A2(new_n335), .A3(new_n338), .A4(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n330), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(KEYINPUT22), .B(G137), .ZN(new_n342));
  INV_X1    g156(.A(G221), .ZN(new_n343));
  INV_X1    g157(.A(G234), .ZN(new_n344));
  NOR3_X1   g158(.A1(new_n343), .A2(new_n344), .A3(G953), .ZN(new_n345));
  XOR2_X1   g159(.A(new_n342), .B(new_n345), .Z(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n341), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n330), .A2(new_n340), .A3(new_n346), .ZN(new_n349));
  INV_X1    g163(.A(G217), .ZN(new_n350));
  INV_X1    g164(.A(G902), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n350), .B1(G234), .B2(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n352), .A2(G902), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n348), .A2(new_n349), .A3(new_n353), .ZN(new_n354));
  XOR2_X1   g168(.A(new_n354), .B(KEYINPUT77), .Z(new_n355));
  NAND3_X1  g169(.A1(new_n348), .A2(new_n351), .A3(new_n349), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(KEYINPUT25), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT25), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n348), .A2(new_n358), .A3(new_n351), .A4(new_n349), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n357), .A2(new_n352), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n355), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n303), .A2(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(G214), .B1(G237), .B2(G902), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G107), .ZN(new_n366));
  OAI21_X1  g180(.A(KEYINPUT78), .B1(new_n366), .B2(G104), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT78), .ZN(new_n368));
  INV_X1    g182(.A(G104), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(new_n369), .A3(G107), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  XNOR2_X1  g185(.A(KEYINPUT79), .B(G101), .ZN(new_n372));
  OAI21_X1  g186(.A(KEYINPUT3), .B1(new_n369), .B2(G107), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT3), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n374), .A2(new_n366), .A3(G104), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n371), .A2(new_n372), .A3(new_n373), .A4(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT80), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n373), .A2(new_n375), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n380), .A2(KEYINPUT80), .A3(new_n372), .A4(new_n371), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n371), .ZN(new_n383));
  OAI21_X1  g197(.A(G101), .B1(new_n383), .B2(new_n379), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n382), .A2(KEYINPUT4), .A3(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n384), .A2(KEYINPUT4), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n385), .A2(new_n387), .A3(new_n257), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n228), .A2(new_n229), .ZN(new_n389));
  INV_X1    g203(.A(new_n225), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n232), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n230), .A2(KEYINPUT68), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n392), .A2(KEYINPUT5), .A3(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT5), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n218), .B1(new_n225), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G101), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n366), .A2(G104), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n369), .A2(G107), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n398), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n401), .B1(new_n378), .B2(new_n381), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n397), .A2(new_n235), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n388), .A2(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(G110), .B(G122), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n388), .A2(new_n405), .A3(new_n403), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n407), .A2(KEYINPUT6), .A3(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT6), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n404), .A2(new_n410), .A3(new_n406), .ZN(new_n411));
  INV_X1    g225(.A(new_n245), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n326), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n213), .A2(new_n214), .A3(G125), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(G953), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(G224), .ZN(new_n417));
  XOR2_X1   g231(.A(new_n415), .B(new_n417), .Z(new_n418));
  NAND3_X1  g232(.A1(new_n409), .A2(new_n411), .A3(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n401), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n382), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n421), .A2(new_n235), .A3(new_n397), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n396), .B1(new_n391), .B2(new_n395), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(new_n235), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n402), .A2(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n405), .B(KEYINPUT8), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n422), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n413), .A2(KEYINPUT83), .ZN(new_n428));
  OR3_X1    g242(.A1(new_n245), .A2(KEYINPUT83), .A3(G125), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n428), .A2(new_n414), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n417), .A2(KEYINPUT7), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n416), .A2(KEYINPUT84), .A3(G224), .ZN(new_n432));
  AND3_X1   g246(.A1(new_n413), .A2(new_n414), .A3(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT7), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT84), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n434), .B1(new_n417), .B2(new_n435), .ZN(new_n436));
  AOI22_X1  g250(.A1(new_n430), .A2(new_n431), .B1(new_n433), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n427), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT85), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n427), .A2(new_n437), .A3(KEYINPUT85), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n440), .A2(new_n441), .A3(new_n408), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n419), .A2(new_n351), .A3(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(G210), .B1(G237), .B2(G902), .ZN(new_n444));
  XOR2_X1   g258(.A(new_n444), .B(KEYINPUT86), .Z(new_n445));
  NAND2_X1  g259(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n419), .A2(new_n442), .A3(new_n351), .A4(new_n444), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n365), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT4), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n449), .B1(new_n378), .B2(new_n381), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n386), .B1(new_n450), .B2(new_n384), .ZN(new_n451));
  AOI211_X1 g265(.A(new_n401), .B(new_n412), .C1(new_n378), .C2(new_n381), .ZN(new_n452));
  AOI22_X1  g266(.A1(new_n451), .A2(new_n215), .B1(new_n452), .B2(KEYINPUT10), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n382), .A2(new_n245), .A3(new_n420), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT81), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT10), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n402), .A2(KEYINPUT81), .A3(new_n245), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n203), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n453), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(G110), .B(G140), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n416), .A2(G227), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n462), .B(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n421), .A2(new_n412), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n456), .A2(new_n458), .A3(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT12), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n467), .B1(new_n460), .B2(KEYINPUT82), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n466), .A2(new_n203), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n468), .B1(new_n466), .B2(new_n203), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n461), .B(new_n464), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n464), .ZN(new_n472));
  AND3_X1   g286(.A1(new_n453), .A2(new_n459), .A3(new_n460), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n460), .B1(new_n453), .B2(new_n459), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(G469), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n476), .A2(new_n477), .A3(new_n351), .ZN(new_n478));
  NAND2_X1  g292(.A1(G469), .A2(G902), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n461), .B1(new_n469), .B2(new_n470), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n472), .ZN(new_n481));
  INV_X1    g295(.A(new_n474), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n482), .A2(new_n461), .A3(new_n464), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n481), .A2(new_n483), .A3(G469), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n478), .A2(new_n479), .A3(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT91), .ZN(new_n486));
  XNOR2_X1  g300(.A(G113), .B(G122), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n487), .B(G104), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n319), .A2(KEYINPUT19), .A3(new_n320), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT19), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n491), .B1(new_n323), .B2(new_n324), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(KEYINPUT89), .B1(new_n493), .B2(G146), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT89), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n490), .A2(new_n492), .A3(new_n495), .A4(new_n204), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(G237), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n498), .A2(new_n416), .A3(G214), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n206), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n188), .A2(G143), .A3(G214), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n500), .A2(new_n246), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n246), .B1(new_n500), .B2(new_n501), .ZN(new_n504));
  OAI21_X1  g318(.A(KEYINPUT88), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n501), .ZN(new_n506));
  AOI21_X1  g320(.A(G143), .B1(new_n188), .B2(G214), .ZN(new_n507));
  OAI21_X1  g321(.A(G131), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT88), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n508), .A2(new_n509), .A3(new_n502), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n329), .A2(new_n497), .A3(new_n505), .A4(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n321), .B(new_n204), .ZN(new_n512));
  NAND2_X1  g326(.A1(KEYINPUT87), .A2(KEYINPUT18), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n500), .B(new_n501), .C1(new_n246), .C2(new_n513), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n512), .B(new_n514), .C1(new_n513), .C2(new_n508), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n489), .B1(new_n511), .B2(new_n515), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n488), .B(KEYINPUT90), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT17), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n508), .A2(new_n518), .A3(new_n502), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n504), .A2(KEYINPUT17), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n519), .A2(new_n328), .A3(new_n337), .A4(new_n520), .ZN(new_n521));
  AND3_X1   g335(.A1(new_n517), .A2(new_n515), .A3(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n486), .B1(new_n516), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT20), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(G475), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n526), .B(new_n351), .C1(new_n516), .C2(new_n522), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n511), .A2(new_n515), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(new_n488), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n517), .A2(new_n515), .A3(new_n521), .ZN(new_n531));
  AOI21_X1  g345(.A(G475), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n532), .A2(new_n523), .A3(new_n524), .A4(new_n351), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n528), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n521), .A2(new_n515), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n488), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n531), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(new_n351), .ZN(new_n538));
  XOR2_X1   g352(.A(KEYINPUT92), .B(G475), .Z(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n534), .A2(new_n541), .ZN(new_n542));
  XOR2_X1   g356(.A(KEYINPUT9), .B(G234), .Z(new_n543));
  NAND3_X1  g357(.A1(new_n543), .A2(G217), .A3(new_n416), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT93), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n545), .B1(new_n224), .B2(G122), .ZN(new_n546));
  INV_X1    g360(.A(G122), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n547), .A2(KEYINPUT93), .A3(G116), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n224), .A2(G122), .ZN(new_n550));
  AND3_X1   g364(.A1(new_n549), .A2(G107), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(G107), .B1(new_n549), .B2(new_n550), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n206), .A2(G128), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT13), .ZN(new_n555));
  OAI21_X1  g369(.A(KEYINPUT94), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n554), .A2(new_n555), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n210), .A2(G143), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT94), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n559), .A2(new_n206), .A3(KEYINPUT13), .A4(G128), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n556), .A2(new_n557), .A3(new_n558), .A4(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(G134), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n558), .A2(new_n554), .A3(new_n194), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n563), .B(KEYINPUT95), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n553), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n558), .A2(new_n554), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(G134), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n563), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n549), .A2(KEYINPUT14), .A3(G107), .A4(new_n550), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n545), .A2(new_n224), .A3(KEYINPUT14), .A4(G122), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n570), .B1(new_n553), .B2(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n544), .B1(new_n565), .B2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n552), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n549), .A2(G107), .A3(new_n550), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n574), .A2(new_n575), .A3(new_n571), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n576), .A2(new_n568), .A3(new_n569), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n553), .A2(new_n562), .A3(new_n564), .ZN(new_n578));
  INV_X1    g392(.A(new_n544), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT96), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n573), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n577), .A2(new_n578), .A3(KEYINPUT96), .A4(new_n579), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n582), .A2(new_n351), .A3(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT15), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n584), .A2(new_n585), .A3(G478), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(G478), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n582), .A2(new_n351), .A3(new_n583), .A4(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(G952), .ZN(new_n590));
  AOI211_X1 g404(.A(G953), .B(new_n590), .C1(G234), .C2(G237), .ZN(new_n591));
  OAI211_X1 g405(.A(G902), .B(G953), .C1(new_n344), .C2(new_n498), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(KEYINPUT97), .ZN(new_n593));
  XOR2_X1   g407(.A(KEYINPUT21), .B(G898), .Z(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n591), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  NOR3_X1   g410(.A1(new_n542), .A2(new_n589), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n343), .B1(new_n543), .B2(new_n351), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n448), .A2(new_n485), .A3(new_n597), .A4(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n363), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(new_n372), .ZN(G3));
  INV_X1    g416(.A(new_n444), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n443), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n365), .B1(new_n604), .B2(new_n447), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT33), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n582), .A2(new_n606), .A3(new_n583), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n573), .A2(KEYINPUT33), .A3(new_n580), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n607), .A2(G478), .A3(new_n351), .A4(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(G478), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n584), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n542), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n596), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n605), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT98), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n605), .A2(new_n614), .A3(KEYINPUT98), .A4(new_n615), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n361), .A2(new_n598), .ZN(new_n621));
  OAI21_X1  g435(.A(G472), .B1(new_n272), .B2(G902), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n622), .A2(new_n286), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n621), .A2(new_n485), .A3(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n620), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT34), .B(G104), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G6));
  NAND2_X1  g442(.A1(new_n530), .A2(new_n531), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n629), .A2(new_n524), .A3(new_n526), .A4(new_n351), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n527), .A2(KEYINPUT20), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n538), .A2(KEYINPUT99), .A3(new_n540), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT99), .ZN(new_n634));
  AOI21_X1  g448(.A(G902), .B1(new_n536), .B2(new_n531), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n634), .B1(new_n635), .B2(new_n539), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n589), .A2(new_n615), .A3(new_n632), .A4(new_n637), .ZN(new_n638));
  OR2_X1    g452(.A1(new_n638), .A2(KEYINPUT100), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(KEYINPUT100), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n639), .A2(new_n605), .A3(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT101), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT100), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n638), .B(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n645), .A2(KEYINPUT101), .A3(new_n605), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n625), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT35), .B(G107), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G9));
  NOR2_X1   g464(.A1(new_n347), .A2(KEYINPUT36), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n341), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n353), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n360), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n654), .A2(new_n286), .A3(new_n622), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT102), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n623), .A2(KEYINPUT102), .A3(new_n654), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n659), .A2(new_n600), .ZN(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT37), .B(G110), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G12));
  NAND2_X1  g476(.A1(new_n485), .A2(new_n599), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n301), .B1(new_n285), .B2(new_n288), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(G900), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n593), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n667), .A2(new_n591), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n632), .A2(new_n637), .A3(new_n669), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n586), .A2(new_n588), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n665), .A2(new_n605), .A3(new_n654), .A4(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G128), .ZN(G30));
  XOR2_X1   g488(.A(new_n668), .B(KEYINPUT39), .Z(new_n675));
  NAND3_X1  g489(.A1(new_n485), .A2(new_n599), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(KEYINPUT40), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n542), .A2(new_n589), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n446), .A2(new_n447), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(KEYINPUT38), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT38), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n446), .A2(new_n681), .A3(new_n447), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n678), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT40), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n485), .A2(new_n684), .A3(new_n599), .A4(new_n675), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n297), .A2(new_n192), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n277), .A2(new_n250), .A3(new_n276), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n351), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n290), .B1(new_n686), .B2(new_n689), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n690), .B1(new_n285), .B2(new_n288), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n677), .A2(new_n683), .A3(new_n685), .A4(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n654), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n364), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(new_n206), .ZN(G45));
  NOR2_X1   g511(.A1(new_n613), .A2(new_n668), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n665), .A2(new_n605), .A3(new_n654), .A4(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G146), .ZN(G48));
  AOI21_X1  g514(.A(new_n477), .B1(new_n476), .B2(new_n351), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n702), .A2(new_n599), .A3(new_n478), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n703), .A2(new_n664), .A3(new_n361), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n620), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(KEYINPUT41), .B(G113), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G15));
  NOR2_X1   g521(.A1(new_n641), .A2(new_n642), .ZN(new_n708));
  AOI21_X1  g522(.A(KEYINPUT101), .B1(new_n645), .B2(new_n605), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n704), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G116), .ZN(G18));
  AND2_X1   g525(.A1(new_n303), .A2(new_n597), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n604), .A2(new_n447), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n364), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n703), .A2(new_n714), .A3(new_n694), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G119), .ZN(G21));
  XNOR2_X1  g531(.A(new_n622), .B(KEYINPUT103), .ZN(new_n718));
  OR2_X1    g532(.A1(new_n293), .A2(new_n192), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n266), .A2(new_n271), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n274), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NOR4_X1   g535(.A1(new_n703), .A2(new_n718), .A3(new_n361), .A4(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n542), .A2(KEYINPUT104), .A3(new_n589), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT104), .ZN(new_n724));
  AOI22_X1  g538(.A1(new_n528), .A2(new_n533), .B1(new_n538), .B2(new_n540), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n724), .B1(new_n725), .B2(new_n671), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n713), .A2(new_n723), .A3(new_n726), .A4(new_n364), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n727), .A2(new_n596), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n722), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G122), .ZN(G24));
  NOR3_X1   g544(.A1(new_n718), .A2(new_n694), .A3(new_n721), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n703), .A2(new_n714), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n731), .A2(new_n732), .A3(new_n698), .ZN(new_n733));
  XNOR2_X1  g547(.A(KEYINPUT105), .B(G125), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n733), .B(new_n734), .ZN(G27));
  INV_X1    g549(.A(KEYINPUT42), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n361), .B1(new_n289), .B2(new_n302), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT106), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n485), .A2(new_n738), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n478), .A2(new_n484), .A3(KEYINPUT106), .A4(new_n479), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n446), .A2(new_n364), .A3(new_n447), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n741), .A2(new_n598), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n737), .A2(new_n739), .A3(new_n740), .A4(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(new_n698), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n736), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n302), .A2(new_n275), .A3(new_n284), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n362), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n747), .A2(new_n736), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n739), .A2(new_n740), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n748), .A2(new_n749), .A3(new_n698), .A4(new_n742), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n745), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G131), .ZN(G33));
  NAND3_X1  g566(.A1(new_n742), .A2(new_n739), .A3(new_n740), .ZN(new_n753));
  INV_X1    g567(.A(new_n672), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n753), .A2(new_n363), .A3(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(new_n194), .ZN(G36));
  XNOR2_X1  g570(.A(new_n725), .B(KEYINPUT108), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n757), .A2(KEYINPUT43), .A3(new_n612), .ZN(new_n758));
  AOI21_X1  g572(.A(KEYINPUT43), .B1(new_n725), .B2(new_n612), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT107), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  OR2_X1    g575(.A1(new_n759), .A2(new_n760), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n758), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n623), .B1(new_n763), .B2(KEYINPUT109), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT109), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n758), .A2(new_n761), .A3(new_n765), .A4(new_n762), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n764), .A2(new_n654), .A3(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT44), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT46), .ZN(new_n770));
  INV_X1    g584(.A(new_n468), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n402), .A2(KEYINPUT81), .A3(new_n245), .ZN(new_n772));
  AOI21_X1  g586(.A(KEYINPUT81), .B1(new_n402), .B2(new_n245), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n402), .A2(new_n245), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n772), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n771), .B1(new_n775), .B2(new_n460), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n466), .A2(new_n203), .A3(new_n468), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n464), .B1(new_n778), .B2(new_n461), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT45), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n473), .A2(new_n474), .A3(new_n472), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  AOI21_X1  g596(.A(KEYINPUT45), .B1(new_n481), .B2(new_n483), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n770), .B(G469), .C1(new_n784), .C2(G902), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n780), .B1(new_n779), .B2(new_n781), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n481), .A2(new_n483), .A3(KEYINPUT45), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n786), .A2(G469), .A3(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n788), .A2(KEYINPUT46), .A3(new_n479), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n785), .A2(new_n478), .A3(new_n789), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n790), .A2(new_n599), .A3(new_n675), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n741), .B(KEYINPUT110), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n764), .A2(KEYINPUT44), .A3(new_n654), .A4(new_n766), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n769), .A2(new_n791), .A3(new_n793), .A4(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G137), .ZN(G39));
  INV_X1    g610(.A(KEYINPUT47), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT111), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n790), .A2(new_n798), .A3(new_n599), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n798), .B1(new_n790), .B2(new_n599), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n797), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n788), .A2(KEYINPUT46), .A3(new_n479), .ZN(new_n802));
  AOI21_X1  g616(.A(KEYINPUT46), .B1(new_n788), .B2(new_n479), .ZN(new_n803));
  AOI211_X1 g617(.A(G469), .B(G902), .C1(new_n471), .C2(new_n475), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  OAI21_X1  g619(.A(KEYINPUT111), .B1(new_n805), .B2(new_n598), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n790), .A2(new_n798), .A3(new_n599), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n806), .A2(KEYINPUT47), .A3(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n741), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n664), .A2(new_n809), .A3(new_n361), .A4(new_n698), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(KEYINPUT112), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n801), .A2(new_n808), .A3(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(G140), .ZN(G42));
  INV_X1    g627(.A(KEYINPUT121), .ZN(new_n814));
  XOR2_X1   g628(.A(KEYINPUT117), .B(KEYINPUT51), .Z(new_n815));
  NOR3_X1   g629(.A1(new_n718), .A2(new_n361), .A3(new_n721), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n763), .A2(new_n591), .A3(new_n816), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n680), .A2(new_n682), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n701), .A2(new_n804), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n818), .A2(new_n599), .A3(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n817), .A2(new_n365), .A3(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT50), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n817), .A2(KEYINPUT50), .A3(new_n365), .A4(new_n820), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n799), .A2(new_n800), .A3(new_n797), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT47), .B1(new_n806), .B2(new_n807), .ZN(new_n828));
  OAI21_X1  g642(.A(KEYINPUT118), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n819), .A2(new_n598), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT118), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n801), .A2(new_n808), .A3(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n829), .A2(new_n830), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n817), .A2(new_n793), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n826), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n819), .A2(new_n591), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n837), .A2(new_n742), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n838), .A2(new_n763), .A3(new_n731), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n837), .A2(new_n362), .A3(new_n691), .A4(new_n742), .ZN(new_n840));
  OR2_X1    g654(.A1(new_n840), .A2(new_n612), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n839), .B1(new_n841), .B2(new_n542), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n815), .B1(new_n836), .B2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT51), .ZN(new_n845));
  OAI211_X1 g659(.A(KEYINPUT119), .B(new_n839), .C1(new_n841), .C2(new_n542), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT119), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n838), .A2(new_n763), .A3(new_n731), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n840), .A2(new_n542), .A3(new_n612), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n847), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n845), .B1(new_n846), .B2(new_n850), .ZN(new_n851));
  AOI22_X1  g665(.A1(new_n801), .A2(new_n808), .B1(new_n598), .B2(new_n819), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n851), .B(new_n825), .C1(new_n852), .C2(new_n834), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n817), .A2(new_n732), .ZN(new_n854));
  INV_X1    g668(.A(new_n747), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n838), .A2(new_n855), .A3(new_n763), .ZN(new_n856));
  XNOR2_X1  g670(.A(KEYINPUT120), .B(KEYINPUT48), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n856), .B(new_n857), .ZN(new_n858));
  OAI211_X1 g672(.A(G952), .B(new_n416), .C1(new_n840), .C2(new_n613), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n853), .A2(new_n854), .A3(new_n860), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n814), .B1(new_n844), .B2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT114), .ZN(new_n863));
  OR3_X1    g677(.A1(new_n670), .A2(new_n863), .A3(new_n589), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n863), .B1(new_n670), .B2(new_n589), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(new_n809), .ZN(new_n867));
  NOR4_X1   g681(.A1(new_n867), .A2(new_n664), .A3(new_n663), .A4(new_n694), .ZN(new_n868));
  AOI211_X1 g682(.A(new_n868), .B(new_n755), .C1(new_n745), .C2(new_n750), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n705), .A2(new_n710), .A3(new_n729), .A4(new_n716), .ZN(new_n870));
  INV_X1    g684(.A(new_n600), .ZN(new_n871));
  INV_X1    g685(.A(new_n659), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n871), .B1(new_n872), .B2(new_n737), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n613), .B1(new_n542), .B2(new_n671), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n874), .A2(new_n615), .A3(new_n448), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n624), .A2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n749), .A2(new_n731), .A3(new_n698), .A4(new_n742), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n873), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n870), .A2(new_n879), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n673), .A2(new_n699), .A3(new_n733), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT115), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n727), .A2(new_n691), .A3(new_n668), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n654), .A2(new_n598), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n883), .A2(new_n749), .A3(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n881), .A2(new_n882), .A3(KEYINPUT52), .A4(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n869), .A2(new_n880), .A3(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n885), .A2(new_n673), .A3(new_n699), .A4(new_n733), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT52), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n663), .A2(new_n664), .A3(new_n714), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n891), .B(new_n654), .C1(new_n672), .C2(new_n698), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n892), .A2(KEYINPUT52), .A3(new_n733), .A4(new_n885), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n890), .A2(KEYINPUT115), .A3(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(KEYINPUT53), .B1(new_n887), .B2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n755), .ZN(new_n896));
  INV_X1    g710(.A(new_n868), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n751), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  AOI22_X1  g712(.A1(new_n620), .A2(new_n704), .B1(new_n722), .B2(new_n728), .ZN(new_n899));
  AOI22_X1  g713(.A1(new_n647), .A2(new_n704), .B1(new_n715), .B2(new_n712), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n600), .B1(new_n363), .B2(new_n659), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n901), .A2(new_n876), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n899), .A2(new_n900), .A3(new_n902), .A4(new_n878), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n898), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n890), .A2(new_n893), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT53), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(KEYINPUT54), .B1(new_n895), .B2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT54), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n906), .B1(new_n887), .B2(new_n894), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n904), .A2(new_n905), .A3(KEYINPUT53), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(KEYINPUT116), .B1(new_n908), .B2(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n912), .A2(KEYINPUT116), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n853), .A2(new_n854), .A3(new_n860), .ZN(new_n916));
  AOI211_X1 g730(.A(new_n842), .B(new_n826), .C1(new_n833), .C2(new_n835), .ZN(new_n917));
  OAI211_X1 g731(.A(KEYINPUT121), .B(new_n916), .C1(new_n917), .C2(new_n815), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n862), .A2(new_n913), .A3(new_n915), .A4(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n590), .A2(new_n416), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n757), .A2(new_n612), .ZN(new_n922));
  OAI21_X1  g736(.A(KEYINPUT49), .B1(new_n701), .B2(new_n804), .ZN(new_n923));
  AND4_X1   g737(.A1(new_n364), .A2(new_n922), .A3(new_n621), .A4(new_n923), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n701), .A2(new_n804), .A3(KEYINPUT49), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT113), .Z(new_n926));
  NAND4_X1  g740(.A1(new_n924), .A2(new_n926), .A3(new_n691), .A4(new_n818), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n921), .A2(new_n927), .ZN(G75));
  NAND2_X1  g742(.A1(new_n590), .A2(G953), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT122), .Z(new_n930));
  NAND2_X1  g744(.A1(new_n895), .A2(new_n907), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n931), .A2(new_n351), .ZN(new_n932));
  AOI21_X1  g746(.A(KEYINPUT56), .B1(new_n932), .B2(G210), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n409), .A2(new_n411), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(new_n418), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT55), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n930), .B1(new_n933), .B2(new_n937), .ZN(new_n938));
  AOI211_X1 g752(.A(KEYINPUT56), .B(new_n936), .C1(new_n932), .C2(new_n445), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n938), .A2(new_n939), .ZN(G51));
  INV_X1    g754(.A(KEYINPUT123), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n931), .A2(new_n351), .A3(new_n788), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n479), .B(KEYINPUT57), .Z(new_n943));
  AND3_X1   g757(.A1(new_n895), .A2(KEYINPUT54), .A3(new_n907), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n943), .B1(new_n944), .B2(new_n908), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n942), .B1(new_n945), .B2(new_n476), .ZN(new_n946));
  INV_X1    g760(.A(new_n930), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n941), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n476), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n931), .A2(new_n909), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n895), .A2(KEYINPUT54), .A3(new_n907), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n949), .B1(new_n952), .B2(new_n943), .ZN(new_n953));
  OAI211_X1 g767(.A(KEYINPUT123), .B(new_n930), .C1(new_n953), .C2(new_n942), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n948), .A2(new_n954), .ZN(G54));
  NAND3_X1  g769(.A1(new_n932), .A2(KEYINPUT58), .A3(G475), .ZN(new_n956));
  OR2_X1    g770(.A1(new_n956), .A2(new_n629), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n629), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n947), .B1(new_n957), .B2(new_n958), .ZN(G60));
  NAND2_X1  g773(.A1(new_n607), .A2(new_n608), .ZN(new_n960));
  NAND2_X1  g774(.A1(G478), .A2(G902), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT59), .Z(new_n962));
  AOI211_X1 g776(.A(new_n960), .B(new_n962), .C1(new_n950), .C2(new_n951), .ZN(new_n963));
  INV_X1    g777(.A(new_n962), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT116), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n893), .A2(KEYINPUT115), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n966), .A2(new_n898), .A3(new_n903), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n890), .A2(KEYINPUT115), .A3(new_n893), .ZN(new_n968));
  AOI21_X1  g782(.A(KEYINPUT53), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n911), .ZN(new_n970));
  OAI21_X1  g784(.A(KEYINPUT54), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n965), .B1(new_n950), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n964), .B1(new_n972), .B2(new_n914), .ZN(new_n973));
  AOI211_X1 g787(.A(new_n947), .B(new_n963), .C1(new_n973), .C2(new_n960), .ZN(G63));
  AND2_X1   g788(.A1(new_n895), .A2(new_n907), .ZN(new_n975));
  NAND2_X1  g789(.A1(G217), .A2(G902), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT60), .Z(new_n977));
  NAND2_X1  g791(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n348), .A2(new_n349), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n975), .A2(new_n652), .A3(new_n977), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n980), .A2(new_n930), .A3(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT61), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n982), .B(new_n983), .ZN(G66));
  AOI21_X1  g798(.A(new_n416), .B1(new_n594), .B2(G224), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n899), .A2(new_n900), .A3(new_n902), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n985), .B1(new_n986), .B2(new_n416), .ZN(new_n987));
  INV_X1    g801(.A(G898), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n934), .B1(new_n988), .B2(G953), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n987), .B(new_n989), .ZN(G69));
  OAI211_X1 g804(.A(new_n881), .B(KEYINPUT62), .C1(new_n695), .C2(new_n693), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT62), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n892), .A2(new_n733), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n992), .B1(new_n993), .B2(new_n696), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n991), .A2(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(new_n676), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n996), .A2(new_n737), .A3(new_n809), .A4(new_n874), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n995), .A2(new_n795), .A3(new_n812), .A4(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n998), .A2(new_n416), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n269), .B(new_n493), .Z(new_n1000));
  INV_X1    g814(.A(new_n1000), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT124), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n999), .A2(KEYINPUT124), .A3(new_n1001), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n1004), .A2(KEYINPUT126), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g820(.A1(G227), .A2(G900), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n1006), .A2(G953), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g822(.A1(G900), .A2(G953), .ZN(new_n1009));
  INV_X1    g823(.A(new_n727), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n791), .A2(new_n1010), .A3(new_n855), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n795), .A2(new_n812), .A3(new_n1011), .ZN(new_n1012));
  AOI211_X1 g826(.A(KEYINPUT125), .B(new_n755), .C1(new_n745), .C2(new_n750), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT125), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1014), .B1(new_n751), .B2(new_n896), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n881), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  OR2_X1    g830(.A1(new_n1012), .A2(new_n1016), .ZN(new_n1017));
  OAI211_X1 g831(.A(new_n1000), .B(new_n1009), .C1(new_n1017), .C2(G953), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n1018), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1019));
  INV_X1    g833(.A(new_n1019), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1008), .A2(new_n1020), .ZN(new_n1021));
  NAND4_X1  g835(.A1(new_n1019), .A2(new_n1006), .A3(G953), .A4(new_n1007), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1021), .A2(new_n1022), .ZN(G72));
  NAND2_X1  g837(.A1(G472), .A2(G902), .ZN(new_n1024));
  XOR2_X1   g838(.A(new_n1024), .B(KEYINPUT63), .Z(new_n1025));
  NAND2_X1  g839(.A1(new_n298), .A2(new_n264), .ZN(new_n1026));
  OAI211_X1 g840(.A(new_n1025), .B(new_n1026), .C1(new_n969), .C2(new_n970), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n1025), .B1(new_n998), .B2(new_n986), .ZN(new_n1028));
  NAND3_X1  g842(.A1(new_n1028), .A2(new_n192), .A3(new_n297), .ZN(new_n1029));
  NOR3_X1   g843(.A1(new_n1012), .A2(new_n1016), .A3(new_n986), .ZN(new_n1030));
  INV_X1    g844(.A(new_n1025), .ZN(new_n1031));
  OAI211_X1 g845(.A(new_n276), .B(new_n270), .C1(new_n1030), .C2(new_n1031), .ZN(new_n1032));
  INV_X1    g846(.A(KEYINPUT127), .ZN(new_n1033));
  AND3_X1   g847(.A1(new_n1032), .A2(new_n1033), .A3(new_n930), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n1033), .B1(new_n1032), .B2(new_n930), .ZN(new_n1035));
  OAI211_X1 g849(.A(new_n1027), .B(new_n1029), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1036));
  INV_X1    g850(.A(new_n1036), .ZN(G57));
endmodule


