//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 1 1 1 0 0 1 1 0 0 1 0 1 0 1 1 0 0 1 1 1 0 0 1 1 1 1 1 1 0 1 0 0 1 1 1 1 0 1 0 1 0 1 0 0 1 1 0 0 0 0 1 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n623,
    new_n624, new_n625, new_n626, new_n628, new_n629, new_n630, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n786, new_n787, new_n789, new_n790, new_n791, new_n793, new_n794,
    new_n795, new_n796, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n839,
    new_n840, new_n842, new_n843, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n855, new_n856,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897;
  XNOR2_X1  g000(.A(G120gat), .B(G148gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G176gat), .B(G204gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(G85gat), .A2(G92gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(KEYINPUT7), .ZN(new_n206));
  INV_X1    g005(.A(G99gat), .ZN(new_n207));
  INV_X1    g006(.A(G106gat), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT8), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  OAI211_X1 g008(.A(new_n206), .B(new_n209), .C1(G85gat), .C2(G92gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(G99gat), .B(G106gat), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n210), .B(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(G57gat), .B(G64gat), .ZN(new_n213));
  AOI21_X1  g012(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(G71gat), .B(G78gat), .ZN(new_n216));
  OR2_X1    g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n215), .A2(new_n216), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n212), .B(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT10), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND4_X1  g021(.A1(new_n212), .A2(KEYINPUT10), .A3(new_n217), .A4(new_n218), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(G230gat), .A2(G233gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n220), .A2(new_n225), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n204), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n228), .A2(KEYINPUT96), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n230), .A2(new_n204), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n228), .A2(KEYINPUT96), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n231), .A2(new_n226), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n229), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT94), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT84), .B(KEYINPUT31), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n236), .B(G22gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n237), .B(G50gat), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(G197gat), .B(G204gat), .ZN(new_n240));
  AND2_X1   g039(.A1(G211gat), .A2(G218gat), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n240), .B1(KEYINPUT22), .B2(new_n241), .ZN(new_n242));
  NOR2_X1   g041(.A1(G211gat), .A2(G218gat), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n242), .A2(KEYINPUT85), .A3(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT29), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n242), .B(new_n244), .ZN(new_n247));
  OAI211_X1 g046(.A(new_n245), .B(new_n246), .C1(new_n247), .C2(KEYINPUT85), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(G155gat), .ZN(new_n251));
  INV_X1    g050(.A(G162gat), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT2), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n251), .B(new_n252), .C1(new_n253), .C2(KEYINPUT77), .ZN(new_n254));
  NAND2_X1  g053(.A1(G155gat), .A2(G162gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(G148gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(G141gat), .ZN(new_n258));
  INV_X1    g057(.A(G141gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(G148gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n255), .A2(KEYINPUT2), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT77), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n256), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT75), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n255), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(KEYINPUT75), .A2(G155gat), .A3(G162gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(G141gat), .B(G148gat), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n253), .B1(G155gat), .B2(G162gat), .ZN(new_n269));
  OAI211_X1 g068(.A(new_n266), .B(new_n267), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n251), .A2(new_n252), .A3(KEYINPUT76), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT76), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n272), .B1(G155gat), .B2(G162gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n264), .B1(new_n270), .B2(new_n274), .ZN(new_n275));
  AOI22_X1  g074(.A1(new_n250), .A2(new_n275), .B1(G228gat), .B2(G233gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n261), .A2(new_n262), .ZN(new_n277));
  AND2_X1   g076(.A1(new_n271), .A2(new_n273), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n277), .A2(new_n278), .A3(new_n266), .A4(new_n267), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n279), .A2(new_n249), .A3(new_n264), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n247), .B1(new_n246), .B2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT86), .ZN(new_n282));
  OR2_X1    g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n281), .A2(new_n282), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n276), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  AOI22_X1  g084(.A1(new_n258), .A2(new_n260), .B1(KEYINPUT2), .B2(new_n255), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n266), .A2(new_n267), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AOI22_X1  g087(.A1(new_n254), .A2(new_n255), .B1(new_n262), .B2(KEYINPUT77), .ZN(new_n289));
  AOI22_X1  g088(.A1(new_n288), .A2(new_n278), .B1(new_n261), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n247), .A2(new_n246), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n290), .B1(new_n291), .B2(new_n249), .ZN(new_n292));
  OAI211_X1 g091(.A(G228gat), .B(G233gat), .C1(new_n292), .C2(new_n281), .ZN(new_n293));
  XOR2_X1   g092(.A(G78gat), .B(G106gat), .Z(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n285), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n295), .B1(new_n285), .B2(new_n293), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n239), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n298), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n300), .A2(new_n238), .A3(new_n296), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  XOR2_X1   g101(.A(KEYINPUT80), .B(KEYINPUT0), .Z(new_n303));
  XNOR2_X1  g102(.A(G1gat), .B(G29gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(new_n303), .B(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G57gat), .B(G85gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n305), .B(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n264), .ZN(new_n309));
  NOR3_X1   g108(.A1(new_n286), .A2(new_n274), .A3(new_n287), .ZN(new_n310));
  OAI21_X1  g109(.A(KEYINPUT3), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(G120gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(G113gat), .ZN(new_n313));
  INV_X1    g112(.A(G113gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(G120gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT1), .ZN(new_n317));
  INV_X1    g116(.A(G134gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(G127gat), .ZN(new_n319));
  INV_X1    g118(.A(G127gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(G134gat), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n316), .A2(new_n317), .A3(new_n319), .A4(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n319), .A2(new_n321), .ZN(new_n323));
  XNOR2_X1  g122(.A(G113gat), .B(G120gat), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n323), .B1(new_n324), .B2(KEYINPUT1), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n311), .A2(new_n326), .A3(new_n280), .ZN(new_n327));
  NAND2_X1  g126(.A1(G225gat), .A2(G233gat), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  AND2_X1   g128(.A1(new_n322), .A2(new_n325), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n329), .B1(new_n290), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT4), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n327), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT78), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n334), .B1(new_n275), .B2(new_n326), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n330), .A2(KEYINPUT78), .A3(new_n264), .A4(new_n279), .ZN(new_n336));
  AOI21_X1  g135(.A(KEYINPUT4), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n333), .A2(new_n337), .ZN(new_n338));
  AOI22_X1  g137(.A1(new_n279), .A2(new_n264), .B1(new_n322), .B2(new_n325), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n339), .B1(new_n335), .B2(new_n336), .ZN(new_n340));
  OAI21_X1  g139(.A(KEYINPUT5), .B1(new_n340), .B2(new_n328), .ZN(new_n341));
  OAI21_X1  g140(.A(KEYINPUT79), .B1(new_n338), .B2(new_n341), .ZN(new_n342));
  AOI21_X1  g141(.A(KEYINPUT78), .B1(new_n290), .B2(new_n330), .ZN(new_n343));
  NOR3_X1   g142(.A1(new_n275), .A2(new_n334), .A3(new_n326), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n332), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n275), .A2(new_n326), .ZN(new_n346));
  OAI21_X1  g145(.A(KEYINPUT4), .B1(new_n346), .B2(new_n329), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n345), .A2(new_n347), .A3(new_n327), .ZN(new_n348));
  INV_X1    g147(.A(new_n339), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n349), .B1(new_n343), .B2(new_n344), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(new_n329), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT79), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n348), .A2(new_n351), .A3(new_n352), .A4(KEYINPUT5), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n342), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n332), .B1(new_n335), .B2(new_n336), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT81), .ZN(new_n356));
  NOR3_X1   g155(.A1(new_n275), .A2(KEYINPUT4), .A3(new_n326), .ZN(new_n357));
  OR3_X1    g156(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n329), .A2(KEYINPUT5), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n356), .B1(new_n355), .B2(new_n357), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n358), .A2(new_n327), .A3(new_n359), .A4(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n308), .B1(new_n354), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(KEYINPUT6), .ZN(new_n363));
  AND3_X1   g162(.A1(new_n354), .A2(new_n361), .A3(new_n308), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n364), .A2(new_n362), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT6), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT82), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NOR3_X1   g166(.A1(new_n338), .A2(new_n341), .A3(KEYINPUT79), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT5), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n369), .B1(new_n350), .B2(new_n329), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n352), .B1(new_n370), .B2(new_n348), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n361), .B1(new_n368), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(new_n307), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n354), .A2(new_n361), .A3(new_n308), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n373), .A2(KEYINPUT82), .A3(new_n366), .A4(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n363), .B1(new_n367), .B2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT83), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT72), .ZN(new_n379));
  INV_X1    g178(.A(new_n247), .ZN(new_n380));
  XOR2_X1   g179(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n381));
  NOR2_X1   g180(.A1(G169gat), .A2(G176gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT23), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT65), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n382), .A2(KEYINPUT65), .A3(KEYINPUT23), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT24), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n388), .B1(G183gat), .B2(G190gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(G183gat), .A2(G190gat), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n390), .A2(KEYINPUT24), .ZN(new_n391));
  OAI22_X1  g190(.A1(new_n389), .A2(new_n391), .B1(G183gat), .B2(G190gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n387), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT66), .ZN(new_n394));
  OR3_X1    g193(.A1(new_n382), .A2(new_n394), .A3(KEYINPUT23), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n394), .B1(new_n382), .B2(KEYINPUT23), .ZN(new_n396));
  NAND2_X1  g195(.A1(G169gat), .A2(G176gat), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n381), .B1(new_n393), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT67), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OAI211_X1 g200(.A(KEYINPUT67), .B(new_n381), .C1(new_n393), .C2(new_n398), .ZN(new_n402));
  INV_X1    g201(.A(new_n398), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n390), .A2(KEYINPUT68), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(KEYINPUT24), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n390), .A2(KEYINPUT68), .A3(new_n388), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n405), .B(new_n406), .C1(G183gat), .C2(G190gat), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n403), .A2(new_n407), .A3(KEYINPUT25), .A4(new_n383), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n401), .A2(new_n402), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(G226gat), .A2(G233gat), .ZN(new_n410));
  INV_X1    g209(.A(new_n382), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(KEYINPUT26), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n412), .B(KEYINPUT69), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n413), .B(new_n397), .C1(KEYINPUT26), .C2(new_n411), .ZN(new_n414));
  XOR2_X1   g213(.A(KEYINPUT27), .B(G183gat), .Z(new_n415));
  OAI21_X1  g214(.A(KEYINPUT28), .B1(new_n415), .B2(G190gat), .ZN(new_n416));
  OR3_X1    g215(.A1(new_n415), .A2(KEYINPUT28), .A3(G190gat), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n414), .A2(new_n390), .A3(new_n416), .A4(new_n417), .ZN(new_n418));
  AND3_X1   g217(.A1(new_n409), .A2(new_n410), .A3(new_n418), .ZN(new_n419));
  AOI22_X1  g218(.A1(new_n409), .A2(new_n418), .B1(new_n246), .B2(new_n410), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n380), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n409), .A2(new_n418), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n410), .A2(new_n246), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n409), .A2(new_n410), .A3(new_n418), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n424), .A2(new_n247), .A3(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n379), .B1(new_n421), .B2(new_n426), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n419), .A2(new_n420), .ZN(new_n428));
  AOI21_X1  g227(.A(KEYINPUT72), .B1(new_n428), .B2(new_n247), .ZN(new_n429));
  XNOR2_X1  g228(.A(G8gat), .B(G36gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n430), .B(KEYINPUT73), .ZN(new_n431));
  XNOR2_X1  g230(.A(G64gat), .B(G92gat), .ZN(new_n432));
  XOR2_X1   g231(.A(new_n431), .B(new_n432), .Z(new_n433));
  NOR3_X1   g232(.A1(new_n427), .A2(new_n429), .A3(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(KEYINPUT30), .B1(new_n434), .B2(KEYINPUT74), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n421), .A2(new_n426), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT72), .ZN(new_n437));
  INV_X1    g236(.A(new_n429), .ZN(new_n438));
  INV_X1    g237(.A(new_n433), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT74), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT30), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n433), .B1(new_n427), .B2(new_n429), .ZN(new_n444));
  AND3_X1   g243(.A1(new_n435), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n377), .A2(new_n378), .A3(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n363), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n373), .A2(new_n366), .A3(new_n374), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT82), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n447), .B1(new_n450), .B2(new_n375), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n435), .A2(new_n443), .A3(new_n444), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT83), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n302), .B1(new_n446), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT37), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n437), .A2(new_n438), .A3(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(KEYINPUT37), .B1(new_n427), .B2(new_n429), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n456), .A2(new_n457), .A3(new_n433), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n434), .B1(new_n458), .B2(KEYINPUT38), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n448), .A2(new_n363), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(KEYINPUT38), .B1(new_n436), .B2(KEYINPUT37), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n456), .A2(new_n433), .A3(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n459), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT40), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT39), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n350), .A2(new_n329), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n358), .A2(new_n327), .A3(new_n360), .ZN(new_n468));
  AOI211_X1 g267(.A(new_n466), .B(new_n467), .C1(new_n468), .C2(new_n329), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n468), .A2(new_n466), .A3(new_n329), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(new_n308), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n465), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n467), .B1(new_n468), .B2(new_n329), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT39), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n474), .A2(KEYINPUT40), .A3(new_n308), .A4(new_n470), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n452), .A2(new_n476), .A3(new_n373), .ZN(new_n477));
  AND3_X1   g276(.A1(new_n464), .A2(new_n477), .A3(new_n302), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n422), .A2(new_n326), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n409), .A2(new_n330), .A3(new_n418), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(G227gat), .A2(G233gat), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT33), .ZN(new_n485));
  XNOR2_X1  g284(.A(G15gat), .B(G43gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(G71gat), .B(G99gat), .ZN(new_n487));
  XOR2_X1   g286(.A(new_n486), .B(new_n487), .Z(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n485), .B1(new_n489), .B2(KEYINPUT70), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n490), .B1(KEYINPUT70), .B2(new_n489), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n484), .A2(KEYINPUT32), .A3(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n485), .A2(KEYINPUT32), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n489), .B1(new_n484), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  OR3_X1    g296(.A1(new_n481), .A2(KEYINPUT34), .A3(new_n483), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT34), .B1(new_n481), .B2(new_n483), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT71), .ZN(new_n501));
  OR2_X1    g300(.A1(new_n497), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n497), .A2(new_n501), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n502), .A2(KEYINPUT36), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n496), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n505), .A2(new_n492), .A3(new_n499), .A4(new_n498), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n500), .B1(new_n493), .B2(new_n496), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT36), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n504), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  NOR3_X1   g311(.A1(new_n454), .A2(new_n478), .A3(new_n512), .ZN(new_n513));
  AND3_X1   g312(.A1(new_n302), .A2(new_n506), .A3(new_n507), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n445), .A2(new_n514), .ZN(new_n515));
  AND2_X1   g314(.A1(KEYINPUT87), .A2(KEYINPUT35), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n460), .B1(KEYINPUT87), .B2(KEYINPUT35), .ZN(new_n517));
  NOR3_X1   g316(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n502), .A2(new_n503), .A3(new_n302), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n446), .A2(new_n453), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n518), .B1(new_n520), .B2(KEYINPUT35), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n513), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(G43gat), .B(G50gat), .ZN(new_n523));
  OAI21_X1  g322(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  NOR3_X1   g324(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n527), .B1(G29gat), .B2(G36gat), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT15), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n523), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(G29gat), .ZN(new_n531));
  INV_X1    g330(.A(G36gat), .ZN(new_n532));
  OR3_X1    g331(.A1(new_n531), .A2(new_n532), .A3(KEYINPUT90), .ZN(new_n533));
  OAI21_X1  g332(.A(KEYINPUT90), .B1(new_n531), .B2(new_n532), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n533), .B(new_n534), .C1(new_n525), .C2(new_n526), .ZN(new_n535));
  INV_X1    g334(.A(G43gat), .ZN(new_n536));
  AND2_X1   g335(.A1(new_n536), .A2(G50gat), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n529), .B1(new_n537), .B2(KEYINPUT89), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n538), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n535), .A2(new_n540), .ZN(new_n541));
  OAI22_X1  g340(.A1(new_n530), .A2(new_n539), .B1(new_n523), .B2(new_n541), .ZN(new_n542));
  XOR2_X1   g341(.A(new_n542), .B(KEYINPUT17), .Z(new_n543));
  XNOR2_X1  g342(.A(G15gat), .B(G22gat), .ZN(new_n544));
  OR2_X1    g343(.A1(new_n544), .A2(G1gat), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT16), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n544), .B1(new_n546), .B2(G1gat), .ZN(new_n547));
  INV_X1    g346(.A(G8gat), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n545), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(KEYINPUT92), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT91), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n545), .A2(new_n547), .A3(new_n551), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n552), .B(G8gat), .C1(new_n551), .C2(new_n547), .ZN(new_n553));
  AND2_X1   g352(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n543), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(KEYINPUT93), .B1(new_n554), .B2(new_n542), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(G229gat), .A2(G233gat), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n543), .A2(KEYINPUT93), .A3(new_n554), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT18), .ZN(new_n561));
  OR2_X1    g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  XOR2_X1   g361(.A(new_n554), .B(new_n542), .Z(new_n563));
  XNOR2_X1  g362(.A(new_n558), .B(KEYINPUT13), .ZN(new_n564));
  OR2_X1    g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n560), .A2(new_n561), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n562), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  XOR2_X1   g366(.A(G169gat), .B(G197gat), .Z(new_n568));
  XNOR2_X1  g367(.A(G113gat), .B(G141gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  XOR2_X1   g371(.A(new_n572), .B(KEYINPUT12), .Z(new_n573));
  NAND2_X1  g372(.A1(new_n567), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n573), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n562), .A2(new_n565), .A3(new_n566), .A4(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n235), .B1(new_n522), .B2(new_n578), .ZN(new_n579));
  OAI211_X1 g378(.A(KEYINPUT94), .B(new_n577), .C1(new_n513), .C2(new_n521), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n234), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n212), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n543), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n584));
  OAI211_X1 g383(.A(new_n583), .B(new_n584), .C1(new_n582), .C2(new_n542), .ZN(new_n585));
  XNOR2_X1  g384(.A(G190gat), .B(G218gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT95), .ZN(new_n589));
  XOR2_X1   g388(.A(G134gat), .B(G162gat), .Z(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  OR2_X1    g391(.A1(new_n587), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n587), .A2(new_n592), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT21), .ZN(new_n597));
  OAI211_X1 g396(.A(new_n550), .B(new_n553), .C1(new_n597), .C2(new_n219), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(G183gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n219), .A2(new_n597), .ZN(new_n602));
  INV_X1    g401(.A(G211gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n601), .B(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G127gat), .B(G155gat), .ZN(new_n607));
  NAND2_X1  g406(.A1(G231gat), .A2(G233gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n606), .B(new_n609), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n596), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n581), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(new_n451), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g414(.A(KEYINPUT16), .B(G8gat), .Z(new_n616));
  NAND3_X1  g415(.A1(new_n613), .A2(new_n452), .A3(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT42), .ZN(new_n618));
  OR2_X1    g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g418(.A(G8gat), .B1(new_n612), .B2(new_n445), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n617), .A2(new_n618), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(G1325gat));
  OR2_X1    g421(.A1(new_n612), .A2(new_n508), .ZN(new_n623));
  INV_X1    g422(.A(G15gat), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n511), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(KEYINPUT97), .ZN(new_n626));
  AOI22_X1  g425(.A1(new_n623), .A2(new_n624), .B1(new_n613), .B2(new_n626), .ZN(G1326gat));
  INV_X1    g426(.A(new_n302), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(KEYINPUT43), .B(G22gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(G1327gat));
  INV_X1    g430(.A(new_n610), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n632), .A2(new_n595), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n581), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n635), .A2(new_n531), .A3(new_n451), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT45), .ZN(new_n637));
  NAND2_X1  g436(.A1(KEYINPUT99), .A2(KEYINPUT44), .ZN(new_n638));
  OAI211_X1 g437(.A(new_n596), .B(new_n638), .C1(new_n513), .C2(new_n521), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n520), .A2(KEYINPUT35), .ZN(new_n640));
  INV_X1    g439(.A(new_n518), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n378), .B1(new_n377), .B2(new_n445), .ZN(new_n643));
  NOR3_X1   g442(.A1(new_n451), .A2(new_n452), .A3(KEYINPUT83), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n628), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n464), .A2(new_n477), .A3(new_n302), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n645), .A2(new_n646), .A3(new_n511), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n595), .B1(new_n642), .B2(new_n647), .ZN(new_n648));
  XOR2_X1   g447(.A(KEYINPUT99), .B(KEYINPUT44), .Z(new_n649));
  OAI21_X1  g448(.A(new_n639), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  XOR2_X1   g449(.A(new_n234), .B(KEYINPUT98), .Z(new_n651));
  NOR2_X1   g450(.A1(new_n578), .A2(new_n651), .ZN(new_n652));
  AND3_X1   g451(.A1(new_n650), .A2(new_n610), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(G29gat), .B1(new_n654), .B2(new_n377), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n637), .A2(new_n655), .ZN(G1328gat));
  INV_X1    g455(.A(KEYINPUT100), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n445), .A2(G36gat), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n657), .B1(new_n635), .B2(new_n658), .ZN(new_n659));
  NOR4_X1   g458(.A1(new_n634), .A2(KEYINPUT100), .A3(G36gat), .A4(new_n445), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT46), .ZN(new_n661));
  OR3_X1    g460(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n661), .B1(new_n659), .B2(new_n660), .ZN(new_n663));
  OAI21_X1  g462(.A(G36gat), .B1(new_n654), .B2(new_n445), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(G1329gat));
  OAI21_X1  g464(.A(new_n536), .B1(new_n634), .B2(new_n508), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n653), .A2(G43gat), .A3(new_n512), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g468(.A(KEYINPUT48), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n650), .A2(new_n610), .A3(new_n628), .A4(new_n652), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n670), .B1(new_n671), .B2(G50gat), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT103), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n302), .A2(G50gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(KEYINPUT102), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n581), .A2(new_n633), .A3(new_n675), .ZN(new_n676));
  AND3_X1   g475(.A1(new_n672), .A2(new_n673), .A3(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n673), .B1(new_n672), .B2(new_n676), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT101), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n671), .A2(new_n680), .A3(G50gat), .ZN(new_n681));
  AND2_X1   g480(.A1(new_n681), .A2(new_n676), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n680), .B1(new_n671), .B2(G50gat), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  AOI21_X1  g483(.A(KEYINPUT48), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(KEYINPUT104), .B1(new_n679), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n681), .A2(new_n676), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n670), .B1(new_n687), .B2(new_n683), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT104), .ZN(new_n689));
  OAI211_X1 g488(.A(new_n688), .B(new_n689), .C1(new_n678), .C2(new_n677), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n686), .A2(new_n690), .ZN(G1331gat));
  INV_X1    g490(.A(new_n651), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n522), .A2(new_n577), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(new_n611), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n694), .A2(new_n377), .ZN(new_n695));
  XOR2_X1   g494(.A(KEYINPUT105), .B(G57gat), .Z(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(G1332gat));
  NOR2_X1   g496(.A1(new_n694), .A2(new_n445), .ZN(new_n698));
  NOR2_X1   g497(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n699));
  AND2_X1   g498(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n698), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n701), .B1(new_n698), .B2(new_n699), .ZN(G1333gat));
  NOR2_X1   g501(.A1(new_n694), .A2(new_n508), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n693), .A2(G71gat), .A3(new_n611), .ZN(new_n704));
  OAI22_X1  g503(.A1(new_n703), .A2(G71gat), .B1(new_n511), .B2(new_n704), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g505(.A1(new_n694), .A2(new_n302), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT107), .ZN(new_n708));
  XNOR2_X1  g507(.A(KEYINPUT106), .B(G78gat), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(G1335gat));
  NOR2_X1   g509(.A1(new_n632), .A2(new_n577), .ZN(new_n711));
  AND3_X1   g510(.A1(new_n650), .A2(new_n234), .A3(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(G85gat), .B1(new_n713), .B2(new_n377), .ZN(new_n714));
  OR2_X1    g513(.A1(new_n648), .A2(KEYINPUT108), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n648), .A2(KEYINPUT108), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n715), .A2(new_n711), .A3(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT51), .ZN(new_n718));
  OR2_X1    g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n717), .A2(new_n718), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT109), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(G85gat), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n719), .A2(KEYINPUT109), .A3(new_n720), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n723), .A2(new_n724), .A3(new_n234), .A4(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n714), .B1(new_n726), .B2(new_n377), .ZN(G1336gat));
  NOR3_X1   g526(.A1(new_n692), .A2(new_n445), .A3(G92gat), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n721), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n712), .A2(new_n452), .ZN(new_n730));
  AOI21_X1  g529(.A(KEYINPUT52), .B1(new_n730), .B2(G92gat), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  AOI22_X1  g531(.A1(new_n719), .A2(new_n720), .B1(KEYINPUT110), .B2(new_n728), .ZN(new_n733));
  OR2_X1    g532(.A1(new_n728), .A2(KEYINPUT110), .ZN(new_n734));
  AOI22_X1  g533(.A1(new_n733), .A2(new_n734), .B1(G92gat), .B2(new_n730), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT52), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n732), .B1(new_n735), .B2(new_n736), .ZN(G1337gat));
  OAI21_X1  g536(.A(G99gat), .B1(new_n713), .B2(new_n511), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n723), .A2(new_n207), .A3(new_n234), .A4(new_n725), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n738), .B1(new_n739), .B2(new_n508), .ZN(G1338gat));
  INV_X1    g539(.A(KEYINPUT53), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n713), .A2(new_n302), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n721), .A2(new_n651), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n628), .A2(new_n208), .ZN(new_n744));
  OAI221_X1 g543(.A(new_n741), .B1(new_n208), .B2(new_n742), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  AOI211_X1 g544(.A(new_n692), .B(new_n744), .C1(new_n719), .C2(new_n720), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n742), .A2(new_n208), .ZN(new_n747));
  OAI21_X1  g546(.A(KEYINPUT53), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n745), .A2(new_n748), .ZN(G1339gat));
  NAND2_X1  g548(.A1(new_n563), .A2(new_n564), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT112), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n558), .B1(new_n557), .B2(new_n559), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n572), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n576), .A2(new_n753), .A3(new_n234), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n595), .A2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n233), .ZN(new_n756));
  OAI21_X1  g555(.A(KEYINPUT54), .B1(new_n224), .B2(new_n225), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT54), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n758), .A2(KEYINPUT111), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n757), .B1(new_n227), .B2(new_n759), .ZN(new_n760));
  OR2_X1    g559(.A1(new_n224), .A2(new_n225), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n761), .A2(KEYINPUT111), .A3(KEYINPUT54), .A4(new_n226), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n760), .A2(new_n762), .A3(new_n204), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(KEYINPUT55), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT55), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n760), .A2(new_n762), .A3(new_n765), .A4(new_n204), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n756), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n577), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n755), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n767), .A2(new_n576), .A3(new_n753), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n596), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n769), .A2(new_n610), .A3(new_n771), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n596), .A2(new_n610), .A3(new_n577), .ZN(new_n773));
  INV_X1    g572(.A(new_n234), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(new_n451), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n777), .A2(new_n515), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(G113gat), .B1(new_n779), .B2(new_n578), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n777), .A2(new_n452), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n519), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n577), .A2(new_n314), .ZN(new_n783));
  XOR2_X1   g582(.A(new_n783), .B(KEYINPUT113), .Z(new_n784));
  OAI21_X1  g583(.A(new_n780), .B1(new_n782), .B2(new_n784), .ZN(G1340gat));
  OAI21_X1  g584(.A(G120gat), .B1(new_n779), .B2(new_n692), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n781), .A2(new_n312), .A3(new_n519), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n786), .B1(new_n774), .B2(new_n787), .ZN(G1341gat));
  NOR2_X1   g587(.A1(new_n782), .A2(new_n610), .ZN(new_n789));
  XOR2_X1   g588(.A(new_n789), .B(KEYINPUT114), .Z(new_n790));
  NOR2_X1   g589(.A1(new_n610), .A2(new_n320), .ZN(new_n791));
  AOI22_X1  g590(.A1(new_n790), .A2(new_n320), .B1(new_n778), .B2(new_n791), .ZN(G1342gat));
  NOR3_X1   g591(.A1(new_n782), .A2(G134gat), .A3(new_n595), .ZN(new_n793));
  XNOR2_X1  g592(.A(KEYINPUT115), .B(KEYINPUT56), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n793), .B(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(G134gat), .B1(new_n779), .B2(new_n595), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(G1343gat));
  NOR2_X1   g596(.A1(new_n512), .A2(new_n302), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n781), .A2(new_n798), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n799), .A2(G141gat), .A3(new_n578), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT57), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n632), .B1(new_n755), .B2(new_n768), .ZN(new_n803));
  AOI22_X1  g602(.A1(new_n803), .A2(new_n771), .B1(new_n773), .B2(new_n774), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n802), .B1(new_n804), .B2(new_n302), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n776), .A2(KEYINPUT57), .A3(new_n628), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n512), .A2(new_n377), .A3(new_n452), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(G141gat), .B1(new_n809), .B2(new_n578), .ZN(new_n810));
  XNOR2_X1  g609(.A(KEYINPUT117), .B(KEYINPUT58), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n801), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT116), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n813), .B1(new_n807), .B2(new_n808), .ZN(new_n814));
  INV_X1    g613(.A(new_n808), .ZN(new_n815));
  AOI211_X1 g614(.A(KEYINPUT116), .B(new_n815), .C1(new_n805), .C2(new_n806), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n577), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n800), .B1(new_n817), .B2(G141gat), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT58), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n812), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT118), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  OAI211_X1 g621(.A(KEYINPUT118), .B(new_n812), .C1(new_n818), .C2(new_n819), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(G1344gat));
  AOI21_X1  g623(.A(KEYINPUT119), .B1(new_n805), .B2(new_n806), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT119), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n776), .A2(new_n628), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n827), .B1(new_n828), .B2(new_n802), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n826), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n831), .A2(KEYINPUT59), .A3(new_n234), .A4(new_n808), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n814), .A2(new_n816), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n833), .A2(new_n774), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n832), .B1(new_n834), .B2(KEYINPUT59), .ZN(new_n835));
  INV_X1    g634(.A(new_n799), .ZN(new_n836));
  AOI21_X1  g635(.A(G148gat), .B1(new_n836), .B2(new_n234), .ZN(new_n837));
  AOI22_X1  g636(.A1(new_n835), .A2(G148gat), .B1(KEYINPUT59), .B2(new_n837), .ZN(G1345gat));
  AOI21_X1  g637(.A(G155gat), .B1(new_n836), .B2(new_n632), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n833), .A2(new_n610), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n839), .B1(new_n840), .B2(G155gat), .ZN(G1346gat));
  AOI21_X1  g640(.A(G162gat), .B1(new_n836), .B2(new_n596), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n833), .A2(new_n595), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n842), .B1(new_n843), .B2(G162gat), .ZN(G1347gat));
  NOR2_X1   g643(.A1(new_n445), .A2(new_n451), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n776), .A2(new_n845), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n846), .A2(new_n519), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n847), .B(KEYINPUT120), .ZN(new_n848));
  INV_X1    g647(.A(G169gat), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n848), .A2(new_n849), .A3(new_n577), .ZN(new_n850));
  AND3_X1   g649(.A1(new_n776), .A2(new_n514), .A3(new_n845), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n849), .B1(new_n851), .B2(new_n577), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(KEYINPUT121), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n850), .A2(new_n853), .ZN(G1348gat));
  AOI21_X1  g653(.A(G176gat), .B1(new_n848), .B2(new_n234), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n851), .A2(G176gat), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n855), .B1(new_n651), .B2(new_n856), .ZN(G1349gat));
  NOR2_X1   g656(.A1(new_n610), .A2(new_n415), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n851), .A2(new_n632), .ZN(new_n859));
  AOI22_X1  g658(.A1(new_n847), .A2(new_n858), .B1(new_n859), .B2(G183gat), .ZN(new_n860));
  NOR2_X1   g659(.A1(KEYINPUT122), .A2(KEYINPUT60), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(KEYINPUT122), .A2(KEYINPUT60), .ZN(new_n863));
  XOR2_X1   g662(.A(new_n863), .B(KEYINPUT123), .Z(new_n864));
  XNOR2_X1  g663(.A(new_n862), .B(new_n864), .ZN(G1350gat));
  INV_X1    g664(.A(G190gat), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n866), .B1(new_n851), .B2(new_n596), .ZN(new_n867));
  XNOR2_X1  g666(.A(new_n867), .B(KEYINPUT124), .ZN(new_n868));
  XOR2_X1   g667(.A(new_n868), .B(KEYINPUT61), .Z(new_n869));
  NAND3_X1  g668(.A1(new_n848), .A2(new_n866), .A3(new_n596), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(G1351gat));
  NAND2_X1  g670(.A1(new_n846), .A2(new_n798), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(G197gat), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n873), .A2(new_n874), .A3(new_n577), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n452), .B(new_n511), .C1(new_n825), .C2(new_n829), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n876), .A2(new_n451), .A3(new_n578), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n875), .B1(new_n877), .B2(new_n874), .ZN(G1352gat));
  NOR3_X1   g677(.A1(new_n872), .A2(G204gat), .A3(new_n774), .ZN(new_n879));
  XOR2_X1   g678(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n880));
  OR2_X1    g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n876), .A2(new_n451), .A3(new_n692), .ZN(new_n884));
  INV_X1    g683(.A(G204gat), .ZN(new_n885));
  OAI211_X1 g684(.A(new_n881), .B(new_n883), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n886), .B(KEYINPUT126), .ZN(G1353gat));
  NAND3_X1  g686(.A1(new_n873), .A2(new_n603), .A3(new_n632), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n445), .B1(new_n826), .B2(new_n830), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n889), .A2(new_n377), .A3(new_n632), .A4(new_n511), .ZN(new_n890));
  AND3_X1   g689(.A1(new_n890), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n891));
  AOI21_X1  g690(.A(KEYINPUT63), .B1(new_n890), .B2(G211gat), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n888), .B1(new_n891), .B2(new_n892), .ZN(G1354gat));
  NAND4_X1  g692(.A1(new_n889), .A2(G218gat), .A3(new_n377), .A4(new_n511), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n872), .A2(new_n595), .ZN(new_n895));
  OAI22_X1  g694(.A1(new_n894), .A2(new_n595), .B1(G218gat), .B2(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT127), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n896), .B(new_n897), .ZN(G1355gat));
endmodule


