//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 1 1 1 1 1 1 1 1 1 1 0 0 1 1 1 0 0 0 0 0 0 1 0 1 1 0 0 1 0 0 0 1 1 0 1 1 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:29 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054;
  INV_X1    g000(.A(KEYINPUT76), .ZN(new_n187));
  INV_X1    g001(.A(G119), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G128), .ZN(new_n189));
  INV_X1    g003(.A(G128), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G119), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT24), .B(G110), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  OAI21_X1  g008(.A(KEYINPUT23), .B1(new_n190), .B2(G119), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT73), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT73), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n189), .A2(new_n197), .A3(KEYINPUT23), .ZN(new_n198));
  OR3_X1    g012(.A1(new_n188), .A2(KEYINPUT74), .A3(G128), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n191), .A2(KEYINPUT74), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n196), .A2(new_n198), .A3(new_n199), .A4(new_n200), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n190), .A2(KEYINPUT23), .A3(G119), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n194), .B1(new_n203), .B2(G110), .ZN(new_n204));
  INV_X1    g018(.A(G140), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G125), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n206), .A2(KEYINPUT16), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT75), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  XNOR2_X1  g023(.A(G125), .B(G140), .ZN(new_n210));
  AOI21_X1  g024(.A(KEYINPUT75), .B1(new_n210), .B2(KEYINPUT16), .ZN(new_n211));
  OAI211_X1 g025(.A(G146), .B(new_n209), .C1(new_n211), .C2(new_n207), .ZN(new_n212));
  INV_X1    g026(.A(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n204), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G125), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G140), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n206), .A2(new_n217), .A3(KEYINPUT16), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n207), .B1(new_n218), .B2(new_n208), .ZN(new_n219));
  INV_X1    g033(.A(new_n209), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n213), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(new_n212), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n192), .A2(new_n193), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n223), .B1(new_n203), .B2(G110), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n215), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(KEYINPUT22), .B(G137), .ZN(new_n227));
  INV_X1    g041(.A(G221), .ZN(new_n228));
  INV_X1    g042(.A(G234), .ZN(new_n229));
  NOR3_X1   g043(.A1(new_n228), .A2(new_n229), .A3(G953), .ZN(new_n230));
  XOR2_X1   g044(.A(new_n227), .B(new_n230), .Z(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n226), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(KEYINPUT72), .B(G902), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n215), .A2(new_n225), .A3(new_n231), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT25), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n233), .A2(KEYINPUT25), .A3(new_n234), .A4(new_n235), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G217), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n241), .B1(new_n234), .B2(G234), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n187), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n242), .ZN(new_n244));
  AOI211_X1 g058(.A(KEYINPUT76), .B(new_n244), .C1(new_n238), .C2(new_n239), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n233), .A2(new_n235), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n242), .A2(G902), .ZN(new_n249));
  XNOR2_X1  g063(.A(KEYINPUT77), .B(KEYINPUT78), .ZN(new_n250));
  XOR2_X1   g064(.A(new_n249), .B(new_n250), .Z(new_n251));
  NAND2_X1  g065(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n246), .A2(new_n252), .ZN(new_n253));
  NOR2_X1   g067(.A1(G472), .A2(G902), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT28), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT66), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT2), .ZN(new_n257));
  INV_X1    g071(.A(G113), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n256), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  OAI21_X1  g073(.A(KEYINPUT66), .B1(KEYINPUT2), .B2(G113), .ZN(new_n260));
  AOI22_X1  g074(.A1(new_n259), .A2(new_n260), .B1(KEYINPUT2), .B2(G113), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n188), .A2(G116), .ZN(new_n262));
  INV_X1    g076(.A(G116), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G119), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n261), .B(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(KEYINPUT64), .B1(new_n213), .B2(G143), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT64), .ZN(new_n268));
  INV_X1    g082(.A(G143), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n268), .A2(new_n269), .A3(G146), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n213), .A2(G143), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AND2_X1   g087(.A1(KEYINPUT0), .A2(G128), .ZN(new_n274));
  NOR2_X1   g088(.A1(KEYINPUT0), .A2(G128), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n213), .A2(G143), .ZN(new_n277));
  OAI21_X1  g091(.A(KEYINPUT65), .B1(new_n269), .B2(G146), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT65), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n279), .A2(new_n213), .A3(G143), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n277), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n273), .A2(new_n276), .B1(new_n281), .B2(new_n274), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT11), .ZN(new_n283));
  INV_X1    g097(.A(G134), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n283), .B1(new_n284), .B2(G137), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(G137), .ZN(new_n286));
  INV_X1    g100(.A(G137), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n287), .A2(KEYINPUT11), .A3(G134), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n285), .A2(new_n286), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(G131), .ZN(new_n290));
  INV_X1    g104(.A(G131), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n285), .A2(new_n288), .A3(new_n291), .A4(new_n286), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n277), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n279), .B1(G143), .B2(new_n213), .ZN(new_n295));
  NOR3_X1   g109(.A1(new_n269), .A2(KEYINPUT65), .A3(G146), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT1), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(G128), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n269), .A2(G146), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n300), .B1(new_n267), .B2(new_n270), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n190), .B1(new_n272), .B2(KEYINPUT1), .ZN(new_n302));
  OAI22_X1  g116(.A1(new_n297), .A2(new_n299), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n287), .A2(G134), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n284), .A2(G137), .ZN(new_n305));
  OAI21_X1  g119(.A(G131), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AND2_X1   g120(.A1(new_n292), .A2(new_n306), .ZN(new_n307));
  AOI22_X1  g121(.A1(new_n282), .A2(new_n293), .B1(new_n303), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n266), .B1(new_n308), .B2(KEYINPUT67), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n273), .A2(new_n276), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n281), .A2(new_n274), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n293), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  AOI211_X1 g126(.A(new_n299), .B(new_n277), .C1(new_n278), .C2(new_n280), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n272), .A2(KEYINPUT1), .ZN(new_n314));
  AOI22_X1  g128(.A1(new_n271), .A2(new_n272), .B1(new_n314), .B2(G128), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n307), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n312), .A2(new_n316), .A3(KEYINPUT67), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n255), .B1(new_n309), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT68), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n312), .A2(new_n316), .ZN(new_n321));
  INV_X1    g135(.A(new_n266), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n308), .A2(new_n266), .ZN(new_n324));
  OAI21_X1  g138(.A(KEYINPUT28), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT67), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n321), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n327), .A2(new_n266), .A3(new_n317), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT68), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n328), .A2(new_n329), .A3(new_n255), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n320), .A2(new_n325), .A3(new_n330), .ZN(new_n331));
  NOR2_X1   g145(.A1(G237), .A2(G953), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G210), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n333), .B(KEYINPUT27), .ZN(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT26), .B(G101), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n334), .B(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n331), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT30), .ZN(new_n339));
  AND3_X1   g153(.A1(new_n312), .A2(new_n316), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n339), .B1(new_n312), .B2(new_n316), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n322), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n323), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n342), .A2(new_n343), .A3(new_n336), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(KEYINPUT31), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT31), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n342), .A2(new_n346), .A3(new_n343), .A4(new_n336), .ZN(new_n347));
  AND2_X1   g161(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  AND3_X1   g162(.A1(new_n338), .A2(new_n348), .A3(KEYINPUT69), .ZN(new_n349));
  AOI21_X1  g163(.A(KEYINPUT69), .B1(new_n338), .B2(new_n348), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n254), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(KEYINPUT32), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT32), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n353), .B(new_n254), .C1(new_n349), .C2(new_n350), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n320), .A2(KEYINPUT70), .A3(new_n330), .ZN(new_n356));
  AND2_X1   g170(.A1(new_n356), .A2(new_n325), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT71), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT70), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n322), .B1(new_n321), .B2(new_n326), .ZN(new_n360));
  AOI211_X1 g174(.A(KEYINPUT68), .B(KEYINPUT28), .C1(new_n360), .C2(new_n317), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n329), .B1(new_n328), .B2(new_n255), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n359), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT29), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n337), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n357), .A2(new_n358), .A3(new_n363), .A4(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n361), .A2(new_n362), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n337), .B1(new_n367), .B2(new_n325), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n342), .A2(new_n343), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n369), .A2(new_n336), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n364), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n363), .A2(new_n356), .A3(new_n325), .A4(new_n365), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(KEYINPUT71), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n366), .A2(new_n371), .A3(new_n373), .A4(new_n234), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G472), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n253), .B1(new_n355), .B2(new_n375), .ZN(new_n376));
  XNOR2_X1  g190(.A(KEYINPUT9), .B(G234), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G902), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n228), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(G469), .ZN(new_n382));
  XNOR2_X1  g196(.A(G110), .B(G140), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n383), .B(KEYINPUT79), .ZN(new_n384));
  INV_X1    g198(.A(G953), .ZN(new_n385));
  AND2_X1   g199(.A1(new_n385), .A2(G227), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n384), .B(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n299), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n281), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n390), .B1(new_n281), .B2(new_n302), .ZN(new_n391));
  XNOR2_X1  g205(.A(KEYINPUT80), .B(G104), .ZN(new_n392));
  OAI21_X1  g206(.A(KEYINPUT3), .B1(new_n392), .B2(G107), .ZN(new_n393));
  INV_X1    g207(.A(G101), .ZN(new_n394));
  INV_X1    g208(.A(G104), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(KEYINPUT80), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT80), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G104), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n396), .A2(new_n398), .A3(G107), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT81), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(KEYINPUT3), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT3), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(KEYINPUT81), .ZN(new_n403));
  INV_X1    g217(.A(G107), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n401), .A2(new_n403), .A3(G104), .A4(new_n404), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n393), .A2(new_n394), .A3(new_n399), .A4(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(G107), .B1(new_n396), .B2(new_n398), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n404), .A2(G104), .ZN(new_n408));
  OAI21_X1  g222(.A(G101), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  AND3_X1   g223(.A1(new_n391), .A2(new_n406), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n303), .B1(new_n406), .B2(new_n409), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n293), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT12), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n406), .A2(new_n409), .ZN(new_n415));
  INV_X1    g229(.A(new_n303), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n391), .A2(new_n406), .A3(new_n409), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n419), .A2(KEYINPUT12), .A3(new_n293), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n414), .A2(new_n420), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n399), .B(new_n405), .C1(new_n407), .C2(new_n402), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(G101), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(KEYINPUT82), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT82), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n422), .A2(new_n425), .A3(G101), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n424), .A2(KEYINPUT4), .A3(new_n426), .A4(new_n406), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT4), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n422), .A2(new_n428), .A3(G101), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT83), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n422), .A2(KEYINPUT83), .A3(new_n428), .A4(G101), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n427), .A2(new_n282), .A3(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n293), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT10), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n416), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n415), .ZN(new_n438));
  AOI22_X1  g252(.A1(new_n437), .A2(new_n438), .B1(new_n418), .B2(new_n436), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n434), .A2(new_n435), .A3(new_n439), .ZN(new_n440));
  AND3_X1   g254(.A1(new_n421), .A2(KEYINPUT84), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(KEYINPUT84), .B1(new_n421), .B2(new_n440), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n388), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  AND3_X1   g257(.A1(new_n434), .A2(new_n435), .A3(new_n439), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n435), .B1(new_n434), .B2(new_n439), .ZN(new_n445));
  NOR3_X1   g259(.A1(new_n444), .A2(new_n445), .A3(new_n388), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n443), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n382), .B1(new_n448), .B2(new_n379), .ZN(new_n449));
  INV_X1    g263(.A(new_n234), .ZN(new_n450));
  XOR2_X1   g264(.A(KEYINPUT85), .B(G469), .Z(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n388), .B1(new_n444), .B2(new_n445), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n421), .A2(new_n387), .A3(new_n440), .ZN(new_n454));
  AOI211_X1 g268(.A(new_n450), .B(new_n452), .C1(new_n453), .C2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n381), .B1(new_n449), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(G210), .B1(G237), .B2(G902), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT88), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n416), .A2(new_n216), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n310), .A2(new_n311), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(G125), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n459), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n282), .A2(new_n216), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n464), .A2(KEYINPUT88), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(G224), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n467), .A2(G953), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n466), .B(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n427), .A2(new_n322), .A3(new_n433), .ZN(new_n470));
  INV_X1    g284(.A(new_n265), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n263), .A2(G119), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT5), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n258), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n262), .A2(new_n264), .A3(KEYINPUT5), .ZN(new_n475));
  AOI22_X1  g289(.A1(new_n261), .A2(new_n471), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n406), .A2(new_n476), .A3(new_n409), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n477), .B(KEYINPUT86), .ZN(new_n478));
  XNOR2_X1  g292(.A(G110), .B(G122), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n470), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(KEYINPUT6), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n470), .A2(new_n478), .ZN(new_n482));
  XOR2_X1   g296(.A(new_n479), .B(KEYINPUT87), .Z(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n482), .A2(KEYINPUT6), .A3(new_n483), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n469), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n468), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n466), .A2(KEYINPUT7), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n460), .A2(new_n462), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT7), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n490), .B1(new_n491), .B2(new_n468), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n479), .B(KEYINPUT8), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n438), .A2(new_n476), .ZN(new_n494));
  INV_X1    g308(.A(new_n477), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n489), .A2(new_n492), .A3(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n480), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n379), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n458), .B1(new_n487), .B2(new_n499), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n466), .B(new_n488), .ZN(new_n501));
  AOI22_X1  g315(.A1(new_n480), .A2(KEYINPUT6), .B1(new_n482), .B2(new_n483), .ZN(new_n502));
  AND3_X1   g316(.A1(new_n482), .A2(KEYINPUT6), .A3(new_n483), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n496), .A2(new_n492), .ZN(new_n505));
  NOR4_X1   g319(.A1(new_n463), .A2(new_n465), .A3(new_n491), .A4(new_n468), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(G902), .B1(new_n507), .B2(new_n480), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n504), .A2(new_n457), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n500), .A2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(G952), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n511), .A2(G953), .ZN(new_n512));
  INV_X1    g326(.A(G237), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n512), .B1(new_n229), .B2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  AOI211_X1 g329(.A(new_n385), .B(new_n234), .C1(G234), .C2(G237), .ZN(new_n516));
  XNOR2_X1  g330(.A(KEYINPUT21), .B(G898), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(G214), .B1(G237), .B2(G902), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n332), .A2(G214), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n269), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n332), .A2(G143), .A3(G214), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n524), .A2(KEYINPUT18), .A3(G131), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n210), .B(new_n213), .ZN(new_n526));
  NAND2_X1  g340(.A1(KEYINPUT18), .A2(G131), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n522), .A2(new_n523), .A3(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n525), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(KEYINPUT90), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT90), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n525), .A2(new_n526), .A3(new_n531), .A4(new_n528), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n524), .A2(G131), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT17), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n522), .A2(new_n291), .A3(new_n523), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n524), .A2(KEYINPUT17), .A3(G131), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n537), .A2(new_n221), .A3(new_n212), .A4(new_n538), .ZN(new_n539));
  XNOR2_X1  g353(.A(G113), .B(G122), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n540), .B(new_n395), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n533), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n541), .B1(new_n533), .B2(new_n539), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n379), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(G475), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n210), .B(KEYINPUT19), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(KEYINPUT91), .B1(new_n548), .B2(G146), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT91), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n547), .A2(new_n550), .A3(new_n213), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n534), .A2(new_n536), .ZN(new_n553));
  AND2_X1   g367(.A1(new_n553), .A2(new_n212), .ZN(new_n554));
  AOI22_X1  g368(.A1(new_n552), .A2(new_n554), .B1(new_n532), .B2(new_n530), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n542), .B1(new_n555), .B2(new_n541), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT20), .ZN(new_n557));
  NOR2_X1   g371(.A1(G475), .A2(G902), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  XOR2_X1   g374(.A(KEYINPUT89), .B(KEYINPUT20), .Z(new_n561));
  AOI21_X1  g375(.A(new_n561), .B1(new_n556), .B2(new_n558), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n546), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  XNOR2_X1  g377(.A(G116), .B(G122), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT14), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n263), .A2(KEYINPUT14), .A3(G122), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n566), .A2(G107), .A3(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n564), .A2(new_n404), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n269), .A2(G128), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n190), .A2(G143), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n571), .A2(new_n572), .A3(new_n284), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n284), .B1(new_n571), .B2(new_n572), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n570), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(KEYINPUT93), .B1(new_n569), .B2(new_n576), .ZN(new_n577));
  OR2_X1    g391(.A1(new_n574), .A2(new_n575), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT93), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n578), .A2(new_n579), .A3(new_n568), .A4(new_n570), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n564), .B(new_n404), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT13), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n571), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n572), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n571), .A2(new_n583), .ZN(new_n586));
  OAI21_X1  g400(.A(G134), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n582), .A2(new_n587), .A3(new_n573), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT92), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n582), .A2(new_n587), .A3(KEYINPUT92), .A4(new_n573), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n581), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NOR3_X1   g406(.A1(new_n377), .A2(new_n241), .A3(G953), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n581), .A2(new_n590), .A3(new_n591), .A4(new_n593), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n450), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(KEYINPUT94), .ZN(new_n598));
  INV_X1    g412(.A(G478), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n599), .A2(KEYINPUT15), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n597), .B(KEYINPUT94), .C1(KEYINPUT15), .C2(new_n599), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n563), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n510), .A2(new_n519), .A3(new_n520), .A4(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n456), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n376), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(G101), .ZN(G3));
  INV_X1    g422(.A(new_n252), .ZN(new_n609));
  NOR3_X1   g423(.A1(new_n243), .A2(new_n245), .A3(new_n609), .ZN(new_n610));
  OAI211_X1 g424(.A(new_n610), .B(new_n381), .C1(new_n449), .C2(new_n455), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT69), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n336), .B1(new_n367), .B2(new_n325), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n345), .A2(new_n347), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n612), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n338), .A2(new_n348), .A3(KEYINPUT69), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n450), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(G472), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n351), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n611), .A2(new_n619), .ZN(new_n620));
  NOR3_X1   g434(.A1(new_n487), .A2(new_n499), .A3(new_n458), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n457), .B1(new_n504), .B2(new_n508), .ZN(new_n622));
  OAI211_X1 g436(.A(new_n519), .B(new_n520), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n595), .A2(new_n596), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(KEYINPUT33), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT33), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n595), .A2(new_n626), .A3(new_n596), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n450), .A2(new_n599), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n597), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n599), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n563), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n623), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n620), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT34), .B(G104), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G6));
  INV_X1    g452(.A(new_n562), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT95), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n556), .A2(new_n561), .A3(new_n558), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  AOI22_X1  g456(.A1(new_n562), .A2(KEYINPUT95), .B1(G475), .B2(new_n545), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n642), .A2(new_n603), .A3(new_n643), .ZN(new_n644));
  OAI21_X1  g458(.A(KEYINPUT96), .B1(new_n623), .B2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n520), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n646), .B1(new_n500), .B2(new_n509), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT96), .ZN(new_n648));
  INV_X1    g462(.A(new_n644), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n647), .A2(new_n648), .A3(new_n649), .A4(new_n519), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n645), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n620), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(new_n404), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT97), .B(KEYINPUT35), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G9));
  INV_X1    g469(.A(new_n243), .ZN(new_n656));
  INV_X1    g470(.A(new_n245), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n232), .A2(KEYINPUT36), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n226), .B(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n251), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n656), .A2(new_n657), .A3(new_n660), .ZN(new_n661));
  OAI211_X1 g475(.A(new_n351), .B(new_n661), .C1(new_n617), .C2(new_n618), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n662), .A2(new_n456), .A3(new_n605), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT98), .ZN(new_n664));
  XNOR2_X1  g478(.A(KEYINPUT37), .B(G110), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G12));
  NAND2_X1  g480(.A1(new_n615), .A2(new_n616), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n353), .B1(new_n667), .B2(new_n254), .ZN(new_n668));
  INV_X1    g482(.A(new_n354), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n375), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  OAI211_X1 g484(.A(new_n661), .B(new_n381), .C1(new_n449), .C2(new_n455), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(G900), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n515), .B1(new_n516), .B2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n647), .A2(new_n649), .A3(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n670), .A2(new_n672), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G128), .ZN(G30));
  XNOR2_X1  g493(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n510), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n500), .A2(new_n509), .A3(new_n680), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n660), .ZN(new_n685));
  NOR3_X1   g499(.A1(new_n243), .A2(new_n245), .A3(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n603), .ZN(new_n687));
  AOI22_X1  g501(.A1(new_n639), .A2(new_n559), .B1(G475), .B2(new_n545), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n686), .A2(new_n689), .A3(new_n520), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n684), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g505(.A(new_n674), .B(KEYINPUT39), .Z(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g507(.A(KEYINPUT40), .B1(new_n456), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n369), .A2(new_n336), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n323), .A2(new_n324), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n379), .B1(new_n698), .B2(new_n336), .ZN(new_n699));
  OAI21_X1  g513(.A(G472), .B1(new_n696), .B2(new_n699), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n700), .B1(new_n668), .B2(new_n669), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT84), .ZN(new_n702));
  AOI21_X1  g516(.A(KEYINPUT12), .B1(new_n419), .B2(new_n293), .ZN(new_n703));
  AOI211_X1 g517(.A(new_n413), .B(new_n435), .C1(new_n417), .C2(new_n418), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n702), .B1(new_n444), .B2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n421), .A2(KEYINPUT84), .A3(new_n440), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n387), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n379), .B1(new_n708), .B2(new_n446), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(G469), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n450), .B1(new_n453), .B2(new_n454), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(new_n451), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n380), .B1(new_n710), .B2(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT40), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n713), .A2(new_n714), .A3(new_n692), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n691), .A2(new_n694), .A3(new_n701), .A4(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT100), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G143), .ZN(G45));
  NOR2_X1   g533(.A1(new_n634), .A2(new_n674), .ZN(new_n720));
  AND2_X1   g534(.A1(new_n720), .A2(new_n647), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n670), .A2(new_n672), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G146), .ZN(G48));
  NOR2_X1   g537(.A1(new_n711), .A2(new_n382), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n724), .A2(new_n455), .A3(new_n380), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n670), .A2(new_n635), .A3(new_n610), .A4(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(KEYINPUT41), .B(G113), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G15));
  NAND4_X1  g542(.A1(new_n651), .A2(new_n670), .A3(new_n610), .A4(new_n725), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G116), .ZN(G18));
  NOR3_X1   g544(.A1(new_n563), .A2(new_n603), .A3(new_n518), .ZN(new_n731));
  AND4_X1   g545(.A1(new_n647), .A2(new_n725), .A3(new_n661), .A4(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n670), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G119), .ZN(G21));
  INV_X1    g548(.A(KEYINPUT101), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n735), .B1(new_n246), .B2(new_n252), .ZN(new_n736));
  NOR4_X1   g550(.A1(new_n243), .A2(new_n245), .A3(KEYINPUT101), .A4(new_n609), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n336), .B1(new_n357), .B2(new_n363), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n254), .B1(new_n739), .B2(new_n614), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n740), .B1(new_n617), .B2(new_n618), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n647), .A2(new_n689), .ZN(new_n743));
  OAI211_X1 g557(.A(new_n712), .B(new_n381), .C1(new_n382), .C2(new_n711), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n743), .A2(new_n518), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G122), .ZN(G24));
  OAI211_X1 g561(.A(new_n740), .B(new_n661), .C1(new_n617), .C2(new_n618), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n720), .A2(new_n647), .A3(new_n725), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(new_n216), .ZN(G27));
  NOR3_X1   g565(.A1(new_n621), .A2(new_n622), .A3(new_n646), .ZN(new_n752));
  NAND2_X1  g566(.A1(G469), .A2(G902), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(KEYINPUT102), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n754), .B1(new_n711), .B2(new_n451), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n443), .A2(G469), .A3(new_n447), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n380), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  AND3_X1   g571(.A1(new_n752), .A2(new_n720), .A3(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(new_n738), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n670), .A2(KEYINPUT42), .A3(new_n758), .A4(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT103), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n670), .A2(new_n761), .A3(new_n758), .A4(new_n610), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT42), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n761), .B1(new_n376), .B2(new_n758), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n760), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G131), .ZN(G33));
  NAND4_X1  g581(.A1(new_n642), .A2(new_n603), .A3(new_n643), .A4(new_n675), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT104), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n752), .A2(new_n757), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(new_n670), .A3(new_n610), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G134), .ZN(G36));
  INV_X1    g588(.A(KEYINPUT45), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n775), .B1(new_n708), .B2(new_n446), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n443), .A2(KEYINPUT45), .A3(new_n447), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n776), .A2(new_n777), .A3(G469), .ZN(new_n778));
  INV_X1    g592(.A(new_n754), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n778), .A2(KEYINPUT46), .A3(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(KEYINPUT46), .B1(new_n778), .B2(new_n779), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT105), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n712), .B(new_n780), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n781), .A2(new_n782), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n381), .B(new_n692), .C1(new_n783), .C2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT106), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n787), .A2(KEYINPUT43), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n688), .A2(new_n633), .A3(new_n789), .ZN(new_n790));
  XOR2_X1   g604(.A(KEYINPUT106), .B(KEYINPUT43), .Z(new_n791));
  AOI22_X1  g605(.A1(new_n628), .A2(new_n629), .B1(new_n599), .B2(new_n631), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n791), .B1(new_n563), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT107), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n790), .A2(new_n793), .A3(KEYINPUT107), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n686), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n798), .A2(KEYINPUT44), .A3(new_n619), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT44), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n790), .A2(new_n793), .A3(KEYINPUT107), .ZN(new_n801));
  AOI21_X1  g615(.A(KEYINPUT107), .B1(new_n790), .B2(new_n793), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n661), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n234), .B1(new_n349), .B2(new_n350), .ZN(new_n804));
  AOI22_X1  g618(.A1(new_n804), .A2(G472), .B1(new_n667), .B2(new_n254), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n800), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n786), .A2(new_n752), .A3(new_n799), .A4(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(KEYINPUT108), .B(G137), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n807), .B(new_n808), .ZN(G39));
  OAI21_X1  g623(.A(new_n381), .B1(new_n783), .B2(new_n784), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT47), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  OAI211_X1 g626(.A(KEYINPUT47), .B(new_n381), .C1(new_n783), .C2(new_n784), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  AOI22_X1  g628(.A1(new_n352), .A2(new_n354), .B1(G472), .B2(new_n374), .ZN(new_n815));
  AND4_X1   g629(.A1(new_n815), .A2(new_n253), .A3(new_n720), .A4(new_n752), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(G140), .ZN(G42));
  NOR2_X1   g632(.A1(new_n724), .A2(new_n455), .ZN(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n820), .A2(KEYINPUT49), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n820), .A2(KEYINPUT49), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n688), .A2(new_n633), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n381), .A2(new_n520), .ZN(new_n824));
  NOR4_X1   g638(.A1(new_n821), .A2(new_n822), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n825), .A2(new_n684), .A3(new_n759), .ZN(new_n826));
  OR2_X1    g640(.A1(new_n826), .A2(new_n701), .ZN(new_n827));
  AOI22_X1  g641(.A1(new_n742), .A2(new_n745), .B1(new_n670), .B2(new_n732), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n828), .A2(new_n729), .A3(new_n726), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n766), .A2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT114), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT110), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n815), .A2(new_n671), .A3(new_n676), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n833), .B1(new_n834), .B2(new_n750), .ZN(new_n835));
  INV_X1    g649(.A(new_n750), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n678), .A2(new_n836), .A3(KEYINPUT110), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT52), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n757), .A2(new_n686), .A3(new_n675), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n839), .A2(new_n743), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n838), .B1(new_n840), .B2(new_n701), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n835), .A2(new_n722), .A3(new_n837), .A4(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n840), .A2(new_n701), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n678), .A2(new_n722), .A3(new_n836), .A4(new_n843), .ZN(new_n844));
  XNOR2_X1  g658(.A(KEYINPUT111), .B(KEYINPUT52), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n842), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n687), .A2(new_n563), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n647), .A2(new_n519), .A3(new_n848), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n619), .A2(new_n611), .A3(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(KEYINPUT109), .B1(new_n850), .B2(new_n663), .ZN(new_n851));
  INV_X1    g665(.A(new_n849), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n852), .A2(new_n805), .A3(new_n713), .A4(new_n610), .ZN(new_n853));
  INV_X1    g667(.A(new_n662), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n606), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT109), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n853), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  AOI22_X1  g671(.A1(new_n376), .A2(new_n606), .B1(new_n620), .B2(new_n635), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n851), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT53), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n500), .A2(new_n520), .A3(new_n509), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n642), .A2(new_n643), .ZN(new_n862));
  NOR4_X1   g676(.A1(new_n861), .A2(new_n603), .A3(new_n862), .A4(new_n674), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n670), .A2(new_n672), .A3(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n748), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(new_n758), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n773), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n859), .A2(new_n860), .A3(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n766), .A2(new_n829), .A3(KEYINPUT114), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n832), .A2(new_n847), .A3(new_n868), .A4(new_n869), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n851), .A2(new_n857), .A3(new_n858), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n773), .A2(new_n864), .A3(new_n866), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n871), .A2(new_n766), .A3(new_n829), .A4(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n844), .A2(new_n838), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n671), .B1(new_n355), .B2(new_n375), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n750), .B1(new_n875), .B2(new_n677), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n876), .A2(KEYINPUT52), .A3(new_n722), .A4(new_n843), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n860), .B1(new_n873), .B2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT54), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n870), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  AOI211_X1 g695(.A(new_n520), .B(new_n744), .C1(new_n682), .C2(new_n683), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n514), .B1(new_n790), .B2(new_n793), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n742), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT50), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n742), .A2(new_n882), .A3(KEYINPUT50), .A4(new_n883), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n861), .A2(new_n744), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(new_n883), .ZN(new_n890));
  OR3_X1    g704(.A1(new_n890), .A2(KEYINPUT116), .A3(new_n748), .ZN(new_n891));
  OAI21_X1  g705(.A(KEYINPUT116), .B1(new_n890), .B2(new_n748), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n889), .A2(new_n610), .A3(new_n515), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n701), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n633), .A2(new_n563), .ZN(new_n895));
  AOI22_X1  g709(.A1(new_n891), .A2(new_n892), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n888), .A2(KEYINPUT51), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n819), .A2(new_n380), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n812), .A2(new_n813), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n742), .A2(new_n883), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n900), .A2(new_n861), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n897), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n894), .A2(new_n563), .A3(new_n633), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n742), .A2(new_n647), .A3(new_n725), .A4(new_n883), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n903), .A2(new_n904), .A3(new_n512), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n670), .A2(new_n759), .ZN(new_n906));
  OR3_X1    g720(.A1(new_n906), .A2(KEYINPUT117), .A3(new_n890), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT48), .ZN(new_n908));
  OAI21_X1  g722(.A(KEYINPUT117), .B1(new_n906), .B2(new_n890), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n908), .B1(new_n907), .B2(new_n909), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n905), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n902), .A2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT115), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n899), .A2(new_n914), .A3(new_n901), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n914), .B1(new_n899), .B2(new_n901), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n888), .A2(new_n896), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n913), .B1(new_n918), .B2(KEYINPUT51), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n872), .A2(new_n857), .A3(new_n851), .A4(new_n858), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n830), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n874), .A2(new_n877), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n921), .A2(KEYINPUT113), .A3(KEYINPUT53), .A4(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n828), .A2(new_n729), .A3(new_n726), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n670), .A2(new_n610), .A3(new_n758), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(KEYINPUT103), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n926), .A2(new_n763), .A3(new_n762), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n924), .B1(new_n927), .B2(new_n760), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n859), .A2(new_n867), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n928), .A2(new_n929), .A3(new_n922), .A4(KEYINPUT53), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT113), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n923), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n847), .A2(new_n928), .A3(new_n929), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT112), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n934), .A2(new_n935), .A3(new_n860), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n935), .B1(new_n934), .B2(new_n860), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n933), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  AOI211_X1 g752(.A(new_n881), .B(new_n919), .C1(new_n938), .C2(KEYINPUT54), .ZN(new_n939));
  NOR2_X1   g753(.A1(G952), .A2(G953), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n827), .B1(new_n939), .B2(new_n940), .ZN(G75));
  NOR2_X1   g755(.A1(new_n385), .A2(G952), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n870), .A2(new_n879), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n450), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n945), .A2(new_n457), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n502), .A2(new_n503), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n469), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n948), .A2(new_n504), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT55), .ZN(new_n950));
  OR2_X1    g764(.A1(new_n950), .A2(KEYINPUT56), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n943), .B1(new_n946), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g766(.A(KEYINPUT118), .B1(new_n945), .B2(new_n457), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT56), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n234), .B1(new_n870), .B2(new_n879), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT118), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n955), .A2(new_n956), .A3(new_n458), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n953), .A2(new_n954), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n952), .B1(new_n950), .B2(new_n958), .ZN(G51));
  NAND2_X1  g773(.A1(new_n453), .A2(new_n454), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT119), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n880), .B1(new_n870), .B2(new_n879), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n881), .A2(new_n962), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n754), .B(KEYINPUT57), .Z(new_n964));
  OAI21_X1  g778(.A(new_n961), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n778), .B(KEYINPUT120), .Z(new_n966));
  NAND2_X1  g780(.A1(new_n955), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n942), .B1(new_n965), .B2(new_n967), .ZN(G54));
  AND2_X1   g782(.A1(KEYINPUT58), .A2(G475), .ZN(new_n969));
  AND3_X1   g783(.A1(new_n955), .A2(new_n556), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n556), .B1(new_n955), .B2(new_n969), .ZN(new_n971));
  NOR3_X1   g785(.A1(new_n970), .A2(new_n971), .A3(new_n942), .ZN(G60));
  XOR2_X1   g786(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n973));
  NOR2_X1   g787(.A1(new_n599), .A2(new_n379), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n973), .B(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n628), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n943), .B1(new_n963), .B2(new_n976), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n842), .A2(new_n846), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n860), .B1(new_n978), .B2(new_n873), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(KEYINPUT112), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n934), .A2(new_n935), .A3(new_n860), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n880), .B1(new_n982), .B2(new_n933), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n975), .B1(new_n983), .B2(new_n881), .ZN(new_n984));
  INV_X1    g798(.A(new_n628), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n977), .B1(new_n984), .B2(new_n985), .ZN(G63));
  XNOR2_X1  g800(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n241), .A2(new_n379), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n987), .B(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n944), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n942), .B1(new_n990), .B2(new_n247), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT61), .ZN(new_n992));
  INV_X1    g806(.A(new_n989), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n993), .B1(new_n870), .B2(new_n879), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(new_n659), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n991), .A2(KEYINPUT123), .A3(new_n992), .A4(new_n995), .ZN(new_n996));
  OR2_X1    g810(.A1(new_n992), .A2(KEYINPUT123), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n992), .A2(KEYINPUT123), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n943), .B1(new_n994), .B2(new_n248), .ZN(new_n999));
  AND3_X1   g813(.A1(new_n944), .A2(new_n659), .A3(new_n989), .ZN(new_n1000));
  OAI211_X1 g814(.A(new_n997), .B(new_n998), .C1(new_n999), .C2(new_n1000), .ZN(new_n1001));
  AND2_X1   g815(.A1(new_n996), .A2(new_n1001), .ZN(G66));
  OAI21_X1  g816(.A(G953), .B1(new_n517), .B2(new_n467), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n859), .A2(new_n924), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n1003), .B1(new_n1004), .B2(G953), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n947), .B1(G898), .B2(new_n385), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1005), .B(new_n1006), .ZN(G69));
  INV_X1    g821(.A(KEYINPUT62), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n678), .A2(new_n836), .ZN(new_n1009));
  AOI22_X1  g823(.A1(new_n1009), .A2(new_n833), .B1(new_n875), .B2(new_n721), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n718), .A2(new_n1008), .A3(new_n837), .A4(new_n1010), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1011), .A2(KEYINPUT124), .ZN(new_n1012));
  AND3_X1   g826(.A1(new_n835), .A2(new_n722), .A3(new_n837), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT124), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n1013), .A2(new_n1014), .A3(new_n1008), .A4(new_n718), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1012), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g830(.A(new_n848), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n861), .B1(new_n1017), .B2(new_n634), .ZN(new_n1018));
  NAND4_X1  g832(.A1(new_n376), .A2(new_n713), .A3(new_n692), .A4(new_n1018), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n817), .A2(new_n807), .A3(new_n1019), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n1008), .B1(new_n1013), .B2(new_n718), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1016), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1023), .A2(new_n385), .ZN(new_n1024));
  NOR2_X1   g838(.A1(new_n340), .A2(new_n341), .ZN(new_n1025));
  XNOR2_X1  g839(.A(new_n1025), .B(new_n547), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g841(.A(KEYINPUT125), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n385), .B1(G227), .B2(G900), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n1026), .B1(G900), .B2(G953), .ZN(new_n1030));
  INV_X1    g844(.A(new_n1030), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n817), .A2(new_n766), .A3(new_n773), .ZN(new_n1032));
  NOR3_X1   g846(.A1(new_n785), .A2(new_n743), .A3(new_n906), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1013), .A2(new_n807), .ZN(new_n1034));
  NOR3_X1   g848(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1031), .B1(new_n1035), .B2(new_n385), .ZN(new_n1036));
  INV_X1    g850(.A(new_n1036), .ZN(new_n1037));
  NAND4_X1  g851(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .A4(new_n1037), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1029), .A2(new_n1028), .ZN(new_n1039));
  OR2_X1    g853(.A1(new_n1029), .A2(new_n1028), .ZN(new_n1040));
  INV_X1    g854(.A(new_n1026), .ZN(new_n1041));
  AOI21_X1  g855(.A(new_n1041), .B1(new_n1023), .B2(new_n385), .ZN(new_n1042));
  OAI211_X1 g856(.A(new_n1039), .B(new_n1040), .C1(new_n1042), .C2(new_n1036), .ZN(new_n1043));
  AND2_X1   g857(.A1(new_n1038), .A2(new_n1043), .ZN(G72));
  NAND3_X1  g858(.A1(new_n1016), .A2(new_n1022), .A3(new_n1004), .ZN(new_n1045));
  XNOR2_X1  g859(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1046));
  NOR2_X1   g860(.A1(new_n618), .A2(new_n379), .ZN(new_n1047));
  XOR2_X1   g861(.A(new_n1046), .B(new_n1047), .Z(new_n1048));
  INV_X1    g862(.A(new_n1048), .ZN(new_n1049));
  AOI21_X1  g863(.A(new_n695), .B1(new_n1045), .B2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g864(.A(new_n1048), .B1(new_n1035), .B2(new_n1004), .ZN(new_n1051));
  XOR2_X1   g865(.A(new_n370), .B(KEYINPUT127), .Z(new_n1052));
  OAI21_X1  g866(.A(new_n943), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NOR3_X1   g867(.A1(new_n696), .A2(new_n370), .A3(new_n1048), .ZN(new_n1054));
  AOI211_X1 g868(.A(new_n1050), .B(new_n1053), .C1(new_n938), .C2(new_n1054), .ZN(G57));
endmodule


