//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 1 0 1 0 1 0 0 1 1 0 0 1 0 0 0 1 0 1 0 0 1 0 0 0 0 0 1 1 1 1 0 0 0 0 0 0 0 0 0 1 1 0 1 1 0 1 0 0 0 0 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:44 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n449, new_n450, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n570, new_n572, new_n573,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n583, new_n584, new_n585, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n615, new_n616,
    new_n617, new_n620, new_n622, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n882, new_n883, new_n884, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1204, new_n1205, new_n1206;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT64), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XNOR2_X1  g013(.A(KEYINPUT65), .B(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  INV_X1    g023(.A(G567), .ZN(new_n449));
  NOR2_X1   g024(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT66), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g027(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NOR4_X1   g029(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(new_n454), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G2106), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n455), .A2(new_n449), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT68), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n466), .A2(new_n463), .A3(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n465), .A2(G137), .A3(new_n467), .A4(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(G101), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(G2105), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n464), .A2(new_n469), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT67), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n473), .A2(new_n474), .A3(G125), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n464), .A2(new_n469), .ZN(new_n477));
  INV_X1    g052(.A(G125), .ZN(new_n478));
  OAI21_X1  g053(.A(KEYINPUT67), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n475), .A2(new_n476), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n472), .B1(new_n480), .B2(G2105), .ZN(G160));
  NAND3_X1  g056(.A1(new_n465), .A2(new_n467), .A3(new_n469), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT69), .ZN(new_n483));
  INV_X1    g058(.A(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(G136), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n484), .A2(G112), .ZN(new_n487));
  OAI21_X1  g062(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n488));
  OAI22_X1  g063(.A1(new_n485), .A2(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n483), .A2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT70), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n483), .A2(KEYINPUT70), .A3(G2105), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n489), .B1(new_n494), .B2(G124), .ZN(G162));
  INV_X1    g070(.A(G138), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n465), .A2(new_n467), .A3(new_n469), .A4(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  NOR3_X1   g074(.A1(new_n496), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n473), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT72), .ZN(new_n503));
  OR2_X1    g078(.A1(G102), .A2(G2105), .ZN(new_n504));
  INV_X1    g079(.A(G114), .ZN(new_n505));
  AND3_X1   g080(.A1(new_n505), .A2(KEYINPUT71), .A3(G2105), .ZN(new_n506));
  AOI21_X1  g081(.A(KEYINPUT71), .B1(new_n505), .B2(G2105), .ZN(new_n507));
  OAI211_X1 g082(.A(G2104), .B(new_n504), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(G126), .A2(G2105), .ZN(new_n509));
  OR2_X1    g084(.A1(new_n482), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g085(.A1(new_n502), .A2(new_n503), .A3(new_n508), .A4(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n498), .A2(KEYINPUT4), .B1(new_n473), .B2(new_n500), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n508), .B1(new_n482), .B2(new_n509), .ZN(new_n513));
  OAI21_X1  g088(.A(KEYINPUT72), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(G164));
  NOR2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  AND2_X1   g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  AND2_X1   g093(.A1(KEYINPUT5), .A2(G543), .ZN(new_n519));
  NOR2_X1   g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  OAI22_X1  g095(.A1(new_n517), .A2(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT73), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  XNOR2_X1  g098(.A(KEYINPUT6), .B(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT5), .B(G543), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n524), .A2(new_n525), .A3(KEYINPUT73), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G88), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n524), .A2(G543), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(G75), .A2(G543), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n519), .A2(new_n520), .ZN(new_n532));
  INV_X1    g107(.A(G62), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  AOI22_X1  g109(.A1(G50), .A2(new_n530), .B1(new_n534), .B2(G651), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n528), .A2(new_n535), .ZN(G303));
  INV_X1    g111(.A(G303), .ZN(G166));
  XNOR2_X1  g112(.A(KEYINPUT74), .B(G89), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n523), .A2(new_n526), .A3(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT7), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n539), .A2(KEYINPUT75), .A3(new_n541), .ZN(new_n542));
  AND2_X1   g117(.A1(G63), .A2(G651), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n530), .A2(G51), .B1(new_n525), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g120(.A(KEYINPUT75), .B1(new_n539), .B2(new_n541), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n545), .A2(new_n546), .ZN(G168));
  AOI22_X1  g122(.A1(new_n525), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n548));
  INV_X1    g123(.A(G651), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT76), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n550), .A2(new_n551), .B1(G52), .B2(new_n530), .ZN(new_n552));
  XNOR2_X1  g127(.A(KEYINPUT77), .B(G90), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n527), .A2(new_n553), .ZN(new_n554));
  OAI21_X1  g129(.A(KEYINPUT76), .B1(new_n548), .B2(new_n549), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n552), .A2(new_n554), .A3(new_n555), .ZN(G301));
  INV_X1    g131(.A(G301), .ZN(G171));
  AOI22_X1  g132(.A1(new_n525), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n558));
  OR2_X1    g133(.A1(new_n558), .A2(new_n549), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n523), .A2(G81), .A3(new_n526), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n530), .A2(G43), .ZN(new_n561));
  AND3_X1   g136(.A1(new_n560), .A2(KEYINPUT78), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g137(.A(KEYINPUT78), .B1(new_n560), .B2(new_n561), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n559), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT79), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OAI211_X1 g141(.A(KEYINPUT79), .B(new_n559), .C1(new_n562), .C2(new_n563), .ZN(new_n567));
  AND2_X1   g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G860), .ZN(G153));
  NAND4_X1  g144(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n570));
  XOR2_X1   g145(.A(new_n570), .B(KEYINPUT80), .Z(G176));
  NAND2_X1  g146(.A1(G1), .A2(G3), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT8), .ZN(new_n573));
  NAND4_X1  g148(.A1(G319), .A2(G483), .A3(G661), .A4(new_n573), .ZN(G188));
  NAND2_X1  g149(.A1(new_n527), .A2(G91), .ZN(new_n575));
  INV_X1    g150(.A(G53), .ZN(new_n576));
  OR3_X1    g151(.A1(new_n529), .A2(KEYINPUT9), .A3(new_n576), .ZN(new_n577));
  OAI21_X1  g152(.A(KEYINPUT9), .B1(new_n529), .B2(new_n576), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n525), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n580), .A2(new_n549), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n575), .A2(new_n579), .A3(new_n581), .ZN(G299));
  NAND2_X1  g157(.A1(new_n539), .A2(new_n541), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT75), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n585), .A2(new_n542), .A3(new_n544), .ZN(G286));
  NAND2_X1  g161(.A1(new_n527), .A2(G87), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n525), .A2(G74), .ZN(new_n588));
  AOI22_X1  g163(.A1(G49), .A2(new_n530), .B1(new_n588), .B2(G651), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n587), .A2(new_n589), .ZN(G288));
  NAND2_X1  g165(.A1(G73), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G61), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n532), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(G651), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n594), .B(KEYINPUT81), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n527), .A2(G86), .B1(G48), .B2(new_n530), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(G305));
  NAND2_X1  g172(.A1(new_n530), .A2(G47), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n525), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n523), .A2(new_n526), .ZN(new_n600));
  INV_X1    g175(.A(G85), .ZN(new_n601));
  OAI221_X1 g176(.A(new_n598), .B1(new_n549), .B2(new_n599), .C1(new_n600), .C2(new_n601), .ZN(G290));
  NAND2_X1  g177(.A1(G301), .A2(G868), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n525), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n604));
  INV_X1    g179(.A(G54), .ZN(new_n605));
  OAI22_X1  g180(.A1(new_n604), .A2(new_n549), .B1(new_n605), .B2(new_n529), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n527), .A2(KEYINPUT10), .A3(G92), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT10), .ZN(new_n608));
  INV_X1    g183(.A(G92), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n600), .B2(new_n609), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n606), .B1(new_n607), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n603), .B1(G868), .B2(new_n611), .ZN(G284));
  OAI21_X1  g187(.A(new_n603), .B1(G868), .B2(new_n611), .ZN(G321));
  NAND2_X1  g188(.A1(G286), .A2(G868), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n614), .A2(KEYINPUT82), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(KEYINPUT82), .ZN(new_n616));
  AND3_X1   g191(.A1(new_n575), .A2(new_n579), .A3(new_n581), .ZN(new_n617));
  OAI211_X1 g192(.A(new_n615), .B(new_n616), .C1(G868), .C2(new_n617), .ZN(G297));
  OAI211_X1 g193(.A(new_n615), .B(new_n616), .C1(G868), .C2(new_n617), .ZN(G280));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n611), .B1(new_n620), .B2(G860), .ZN(G148));
  NAND2_X1  g196(.A1(new_n611), .A2(new_n620), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G868), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(new_n568), .B2(G868), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT83), .Z(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g201(.A1(new_n463), .A2(G2105), .ZN(new_n627));
  INV_X1    g202(.A(new_n627), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n477), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n629), .B(new_n630), .Z(new_n631));
  INV_X1    g206(.A(new_n631), .ZN(new_n632));
  INV_X1    g207(.A(KEYINPUT13), .ZN(new_n633));
  INV_X1    g208(.A(KEYINPUT85), .ZN(new_n634));
  AOI22_X1  g209(.A1(new_n632), .A2(new_n633), .B1(new_n634), .B2(G2100), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n635), .B1(new_n633), .B2(new_n632), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n634), .A2(G2100), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n494), .A2(G123), .ZN(new_n639));
  INV_X1    g214(.A(G2096), .ZN(new_n640));
  OAI21_X1  g215(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n641));
  INV_X1    g216(.A(G111), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n641), .B1(new_n642), .B2(G2105), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n482), .A2(KEYINPUT69), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n482), .A2(KEYINPUT69), .ZN(new_n645));
  AOI21_X1  g220(.A(G2105), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n643), .B1(new_n646), .B2(G135), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n639), .A2(new_n640), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n639), .A2(new_n647), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(G2096), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n638), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(KEYINPUT86), .Z(G156));
  INV_X1    g227(.A(KEYINPUT14), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2427), .B(G2438), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2430), .ZN(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT15), .B(G2435), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n653), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n657), .B1(new_n656), .B2(new_n655), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2451), .B(G2454), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT16), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1341), .B(G1348), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n658), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2443), .B(G2446), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n663), .A2(new_n664), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n665), .A2(new_n666), .A3(G14), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT87), .Z(G401));
  INV_X1    g243(.A(KEYINPUT18), .ZN(new_n669));
  XOR2_X1   g244(.A(G2084), .B(G2090), .Z(new_n670));
  XNOR2_X1  g245(.A(G2067), .B(G2678), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n672), .A2(KEYINPUT17), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n670), .A2(new_n671), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n669), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT88), .B(G2100), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G2072), .B(G2078), .Z(new_n678));
  AOI21_X1  g253(.A(new_n678), .B1(new_n672), .B2(KEYINPUT18), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(new_n640), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n677), .B(new_n680), .ZN(G227));
  XNOR2_X1  g256(.A(G1971), .B(G1976), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1956), .B(G2474), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1961), .B(G1966), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT90), .B(KEYINPUT20), .Z(new_n689));
  OR2_X1    g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n688), .A2(new_n689), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n685), .A2(new_n686), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n684), .A2(new_n693), .ZN(new_n694));
  OR3_X1    g269(.A1(new_n684), .A2(new_n687), .A3(new_n693), .ZN(new_n695));
  NAND4_X1  g270(.A1(new_n690), .A2(new_n691), .A3(new_n694), .A4(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(G1991), .B(G1996), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(G1981), .B(G1986), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT91), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n698), .B(new_n702), .ZN(G229));
  NOR2_X1   g278(.A1(G16), .A2(G23), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT94), .ZN(new_n705));
  INV_X1    g280(.A(G16), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n705), .B1(G288), .B2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT95), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT33), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(G1976), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n709), .B(KEYINPUT33), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G1976), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n706), .A2(G22), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G166), .B2(new_n706), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(G1971), .ZN(new_n718));
  AND2_X1   g293(.A1(new_n706), .A2(G6), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G305), .B2(G16), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT32), .B(G1981), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  AND2_X1   g297(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n720), .A2(new_n722), .ZN(new_n724));
  NOR3_X1   g299(.A1(new_n718), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n713), .A2(new_n715), .A3(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(KEYINPUT96), .B1(new_n726), .B2(KEYINPUT34), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT34), .ZN(new_n729));
  NAND4_X1  g304(.A1(new_n713), .A2(new_n715), .A3(new_n729), .A4(new_n725), .ZN(new_n730));
  INV_X1    g305(.A(G29), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G25), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT92), .ZN(new_n733));
  AOI211_X1 g308(.A(new_n491), .B(new_n484), .C1(new_n644), .C2(new_n645), .ZN(new_n734));
  AOI21_X1  g309(.A(KEYINPUT70), .B1(new_n483), .B2(G2105), .ZN(new_n735));
  OAI21_X1  g310(.A(G119), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g311(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n737));
  INV_X1    g312(.A(G107), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n737), .B1(new_n738), .B2(G2105), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n646), .B2(G131), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n736), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n733), .B1(new_n741), .B2(G29), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT35), .B(G1991), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT93), .Z(new_n744));
  INV_X1    g319(.A(new_n744), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n742), .A2(new_n745), .ZN(new_n747));
  MUX2_X1   g322(.A(G24), .B(G290), .S(G16), .Z(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G1986), .ZN(new_n749));
  NOR3_X1   g324(.A1(new_n746), .A2(new_n747), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n730), .A2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n726), .A2(KEYINPUT96), .A3(KEYINPUT34), .ZN(new_n753));
  AND2_X1   g328(.A1(KEYINPUT97), .A2(KEYINPUT36), .ZN(new_n754));
  NAND4_X1  g329(.A1(new_n728), .A2(new_n752), .A3(new_n753), .A4(new_n754), .ZN(new_n755));
  AND3_X1   g330(.A1(new_n726), .A2(KEYINPUT96), .A3(KEYINPUT34), .ZN(new_n756));
  NOR3_X1   g331(.A1(new_n756), .A2(new_n727), .A3(new_n751), .ZN(new_n757));
  NOR2_X1   g332(.A1(KEYINPUT97), .A2(KEYINPUT36), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n754), .A2(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n755), .B1(new_n757), .B2(new_n760), .ZN(new_n761));
  AND2_X1   g336(.A1(new_n646), .A2(G139), .ZN(new_n762));
  NAND2_X1  g337(.A1(G115), .A2(G2104), .ZN(new_n763));
  INV_X1    g338(.A(G127), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n763), .B1(new_n477), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n765), .A2(G2105), .ZN(new_n766));
  OR2_X1    g341(.A1(new_n766), .A2(KEYINPUT100), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n484), .A2(G103), .A3(G2104), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT25), .Z(new_n769));
  NAND2_X1  g344(.A1(new_n766), .A2(KEYINPUT100), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n767), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT101), .ZN(new_n772));
  NOR3_X1   g347(.A1(new_n762), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n772), .B1(new_n762), .B2(new_n771), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n774), .A2(G29), .A3(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(G29), .A2(G33), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT99), .Z(new_n778));
  NAND2_X1  g353(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n779), .A2(G2072), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n779), .A2(G2072), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n731), .A2(G32), .ZN(new_n783));
  NAND3_X1  g358(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT105), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT26), .Z(new_n786));
  AND2_X1   g361(.A1(new_n627), .A2(G105), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n646), .A2(KEYINPUT103), .A3(G141), .ZN(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  AOI21_X1  g365(.A(KEYINPUT103), .B1(new_n646), .B2(G141), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n788), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT104), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n734), .A2(new_n735), .ZN(new_n794));
  INV_X1    g369(.A(G129), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n793), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  OAI211_X1 g371(.A(KEYINPUT104), .B(G129), .C1(new_n734), .C2(new_n735), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n792), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n783), .B1(new_n798), .B2(new_n731), .ZN(new_n799));
  XNOR2_X1  g374(.A(KEYINPUT27), .B(G1996), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT106), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(G34), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n803), .A2(KEYINPUT24), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n803), .A2(KEYINPUT24), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n731), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G160), .B2(new_n731), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT102), .ZN(new_n808));
  INV_X1    g383(.A(G2084), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n782), .A2(new_n802), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n811), .A2(KEYINPUT107), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT107), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n782), .A2(new_n813), .A3(new_n802), .A4(new_n810), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(G2090), .ZN(new_n816));
  NOR2_X1   g391(.A1(G162), .A2(new_n731), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n731), .A2(G35), .ZN(new_n818));
  OR3_X1    g393(.A1(new_n817), .A2(KEYINPUT29), .A3(new_n818), .ZN(new_n819));
  OAI21_X1  g394(.A(KEYINPUT29), .B1(new_n817), .B2(new_n818), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n816), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n821), .A2(KEYINPUT109), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n706), .A2(G20), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT23), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(new_n617), .B2(new_n706), .ZN(new_n825));
  INV_X1    g400(.A(G1956), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n821), .A2(KEYINPUT109), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n822), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(KEYINPUT110), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT110), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n822), .A2(new_n831), .A3(new_n827), .A4(new_n828), .ZN(new_n832));
  NOR2_X1   g407(.A1(G5), .A2(G16), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT108), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(G301), .B2(new_n706), .ZN(new_n835));
  INV_X1    g410(.A(G1961), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n835), .A2(new_n836), .ZN(new_n838));
  XOR2_X1   g413(.A(KEYINPUT31), .B(G11), .Z(new_n839));
  INV_X1    g414(.A(G28), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n840), .A2(KEYINPUT30), .ZN(new_n841));
  AOI21_X1  g416(.A(G29), .B1(new_n840), .B2(KEYINPUT30), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n839), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n837), .A2(new_n838), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n706), .A2(G4), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(new_n611), .B2(new_n706), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(G1348), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n649), .A2(new_n731), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n731), .A2(G27), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n849), .B1(G164), .B2(new_n731), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n850), .A2(G2078), .ZN(new_n851));
  NOR4_X1   g426(.A1(new_n844), .A2(new_n847), .A3(new_n848), .A4(new_n851), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n819), .A2(new_n816), .A3(new_n820), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n799), .A2(new_n801), .ZN(new_n854));
  NOR2_X1   g429(.A1(G16), .A2(G21), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n855), .B1(G168), .B2(G16), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n856), .A2(G1966), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n808), .A2(new_n809), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n850), .A2(G2078), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n856), .A2(G1966), .ZN(new_n860));
  AND4_X1   g435(.A1(new_n857), .A2(new_n858), .A3(new_n859), .A4(new_n860), .ZN(new_n861));
  NAND4_X1  g436(.A1(new_n852), .A2(new_n853), .A3(new_n854), .A4(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n731), .A2(G26), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n863), .B(KEYINPUT98), .Z(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT28), .ZN(new_n865));
  OAI21_X1  g440(.A(G128), .B1(new_n734), .B2(new_n735), .ZN(new_n866));
  OAI21_X1  g441(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n867));
  INV_X1    g442(.A(G116), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n867), .B1(new_n868), .B2(G2105), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n869), .B1(new_n646), .B2(G140), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n866), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n865), .B1(new_n871), .B2(G29), .ZN(new_n872));
  INV_X1    g447(.A(G2067), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n872), .B(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n706), .A2(G19), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n875), .B1(new_n568), .B2(new_n706), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n876), .A2(G1341), .ZN(new_n877));
  AND2_X1   g452(.A1(new_n876), .A2(G1341), .ZN(new_n878));
  NOR4_X1   g453(.A1(new_n862), .A2(new_n874), .A3(new_n877), .A4(new_n878), .ZN(new_n879));
  NAND4_X1  g454(.A1(new_n815), .A2(new_n830), .A3(new_n832), .A4(new_n879), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n761), .A2(new_n880), .ZN(G311));
  AND3_X1   g456(.A1(new_n815), .A2(new_n879), .A3(new_n832), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n728), .A2(new_n752), .A3(new_n753), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(new_n759), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n882), .A2(new_n884), .A3(new_n830), .A4(new_n755), .ZN(G150));
  AOI22_X1  g460(.A1(new_n525), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n886), .A2(new_n549), .ZN(new_n887));
  INV_X1    g462(.A(G55), .ZN(new_n888));
  INV_X1    g463(.A(G93), .ZN(new_n889));
  OAI221_X1 g464(.A(new_n887), .B1(new_n888), .B2(new_n529), .C1(new_n600), .C2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(G860), .ZN(new_n891));
  XOR2_X1   g466(.A(new_n891), .B(KEYINPUT37), .Z(new_n892));
  INV_X1    g467(.A(KEYINPUT111), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n566), .A2(new_n893), .A3(new_n567), .A4(new_n890), .ZN(new_n894));
  INV_X1    g469(.A(new_n890), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n564), .A2(new_n895), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n566), .A2(new_n567), .A3(new_n890), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(KEYINPUT111), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n611), .A2(G559), .ZN(new_n901));
  XOR2_X1   g476(.A(new_n901), .B(KEYINPUT38), .Z(new_n902));
  XNOR2_X1  g477(.A(new_n900), .B(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  AND2_X1   g479(.A1(new_n904), .A2(KEYINPUT39), .ZN(new_n905));
  INV_X1    g480(.A(G860), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n906), .B1(new_n904), .B2(KEYINPUT39), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n892), .B1(new_n905), .B2(new_n907), .ZN(G145));
  XNOR2_X1  g483(.A(new_n649), .B(G160), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(G162), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n741), .A2(new_n631), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n736), .A2(new_n632), .A3(new_n740), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n646), .A2(G142), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(KEYINPUT113), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n494), .A2(G130), .ZN(new_n916));
  OR2_X1    g491(.A1(G106), .A2(G2105), .ZN(new_n917));
  OAI211_X1 g492(.A(new_n917), .B(G2104), .C1(G118), .C2(new_n484), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n915), .A2(new_n916), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n913), .A2(new_n919), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n916), .A2(new_n918), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n921), .A2(new_n915), .A3(new_n911), .A4(new_n912), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT112), .ZN(new_n924));
  INV_X1    g499(.A(new_n775), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n924), .B1(new_n925), .B2(new_n773), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n774), .A2(KEYINPUT112), .A3(new_n775), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n512), .A2(new_n513), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n866), .A2(new_n930), .A3(new_n870), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n930), .B1(new_n866), .B2(new_n870), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n788), .ZN(new_n934));
  INV_X1    g509(.A(new_n791), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n934), .B1(new_n935), .B2(new_n789), .ZN(new_n936));
  AOI21_X1  g511(.A(KEYINPUT104), .B1(new_n494), .B2(G129), .ZN(new_n937));
  INV_X1    g512(.A(new_n797), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n933), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(G128), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n941), .B1(new_n492), .B2(new_n493), .ZN(new_n942));
  INV_X1    g517(.A(new_n870), .ZN(new_n943));
  OAI22_X1  g518(.A1(new_n942), .A2(new_n943), .B1(new_n512), .B2(new_n513), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n866), .A2(new_n930), .A3(new_n870), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n946), .A2(new_n798), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n929), .B1(new_n940), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n933), .A2(new_n939), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n946), .A2(new_n798), .ZN(new_n950));
  INV_X1    g525(.A(new_n927), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n923), .B1(new_n948), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT114), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n948), .A2(new_n923), .A3(new_n952), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n953), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n952), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n928), .B1(new_n949), .B2(new_n950), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NOR3_X1   g534(.A1(new_n959), .A2(KEYINPUT114), .A3(new_n923), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n910), .B1(new_n956), .B2(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n910), .B1(new_n959), .B2(new_n923), .ZN(new_n962));
  INV_X1    g537(.A(new_n953), .ZN(new_n963));
  AOI21_X1  g538(.A(G37), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n961), .A2(KEYINPUT40), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(KEYINPUT40), .B1(new_n961), .B2(new_n964), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n965), .A2(new_n966), .ZN(G395));
  INV_X1    g542(.A(KEYINPUT116), .ZN(new_n968));
  XNOR2_X1  g543(.A(G288), .B(new_n968), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n969), .B(G305), .ZN(new_n970));
  XNOR2_X1  g545(.A(G303), .B(G290), .ZN(new_n971));
  XOR2_X1   g546(.A(new_n970), .B(new_n971), .Z(new_n972));
  INV_X1    g547(.A(KEYINPUT117), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n972), .A2(new_n973), .A3(KEYINPUT42), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n970), .B(new_n971), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n973), .A2(KEYINPUT42), .ZN(new_n976));
  OR2_X1    g551(.A1(new_n973), .A2(KEYINPUT42), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n974), .A2(new_n978), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n900), .B(new_n622), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT41), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT115), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n617), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(G299), .A2(KEYINPUT115), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n983), .A2(new_n611), .A3(new_n984), .ZN(new_n985));
  NOR3_X1   g560(.A1(new_n617), .A2(new_n611), .A3(new_n982), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n981), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n986), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n983), .A2(new_n611), .A3(new_n984), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n988), .A2(new_n989), .A3(KEYINPUT41), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n980), .A2(new_n991), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n985), .A2(new_n986), .ZN(new_n993));
  OR2_X1    g568(.A1(new_n980), .A2(new_n993), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n979), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n979), .B1(new_n994), .B2(new_n992), .ZN(new_n996));
  OAI21_X1  g571(.A(G868), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n997), .B1(G868), .B2(new_n895), .ZN(G295));
  OAI21_X1  g573(.A(new_n997), .B1(G868), .B2(new_n895), .ZN(G331));
  NAND2_X1  g574(.A1(G168), .A2(G301), .ZN(new_n1000));
  NAND2_X1  g575(.A1(G171), .A2(G286), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  AND2_X1   g578(.A1(new_n898), .A2(KEYINPUT111), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n894), .A2(new_n896), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1003), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n899), .A2(new_n896), .A3(new_n894), .A4(new_n1002), .ZN(new_n1007));
  AND3_X1   g582(.A1(new_n1006), .A2(new_n993), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n991), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n972), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT43), .ZN(new_n1011));
  AND2_X1   g586(.A1(new_n987), .A2(new_n990), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1002), .B1(new_n897), .B2(new_n899), .ZN(new_n1013));
  AND4_X1   g588(.A1(new_n899), .A2(new_n896), .A3(new_n894), .A4(new_n1002), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1012), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1006), .A2(new_n993), .A3(new_n1007), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1015), .A2(new_n975), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G37), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1010), .A2(new_n1011), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT118), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1021));
  AOI21_X1  g596(.A(G37), .B1(new_n1021), .B2(new_n972), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT118), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n1022), .A2(new_n1023), .A3(new_n1011), .A4(new_n1017), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1010), .A2(new_n1018), .A3(new_n1017), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT43), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1020), .A2(new_n1024), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT44), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1026), .A2(KEYINPUT44), .A3(new_n1019), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(G397));
  XNOR2_X1  g606(.A(new_n939), .B(G1996), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n871), .A2(G2067), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n866), .A2(new_n873), .A3(new_n870), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n741), .A2(new_n744), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n1034), .ZN(new_n1039));
  AND2_X1   g614(.A1(G160), .A2(G40), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT45), .ZN(new_n1041));
  INV_X1    g616(.A(G1384), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1042), .B1(new_n512), .B2(new_n513), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1040), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  AND3_X1   g620(.A1(new_n1039), .A2(KEYINPUT126), .A3(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT126), .B1(new_n1039), .B2(new_n1045), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1044), .A2(G1996), .ZN(new_n1048));
  XOR2_X1   g623(.A(new_n1048), .B(KEYINPUT46), .Z(new_n1049));
  OAI21_X1  g624(.A(new_n1045), .B1(new_n1035), .B2(new_n939), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  XNOR2_X1  g626(.A(new_n1051), .B(KEYINPUT47), .ZN(new_n1052));
  XNOR2_X1  g627(.A(new_n741), .B(new_n745), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1044), .B1(new_n1036), .B2(new_n1053), .ZN(new_n1054));
  NOR3_X1   g629(.A1(new_n1044), .A2(G1986), .A3(G290), .ZN(new_n1055));
  XNOR2_X1  g630(.A(new_n1055), .B(KEYINPUT48), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1052), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  NOR3_X1   g632(.A1(new_n1046), .A2(new_n1047), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(G1966), .ZN(new_n1059));
  AOI21_X1  g634(.A(G1384), .B1(new_n511), .B2(new_n514), .ZN(new_n1060));
  AND2_X1   g635(.A1(new_n1060), .A2(KEYINPUT45), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1043), .A2(new_n1041), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1040), .A2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1059), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT50), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1065), .B(new_n1042), .C1(new_n512), .C2(new_n513), .ZN(new_n1066));
  AND3_X1   g641(.A1(new_n1066), .A2(G40), .A3(G160), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1067), .B(new_n809), .C1(new_n1060), .C2(new_n1065), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1064), .A2(G168), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(G8), .ZN(new_n1070));
  AOI21_X1  g645(.A(G168), .B1(new_n1064), .B2(new_n1068), .ZN(new_n1071));
  OAI21_X1  g646(.A(KEYINPUT51), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT51), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1069), .A2(new_n1073), .A3(G8), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(KEYINPUT62), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT62), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1072), .A2(new_n1074), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(G8), .ZN(new_n1079));
  NOR2_X1   g654(.A1(G166), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(KEYINPUT119), .A2(KEYINPUT55), .ZN(new_n1081));
  OR2_X1    g656(.A1(KEYINPUT119), .A2(KEYINPUT55), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1080), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  AND2_X1   g658(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1043), .ZN(new_n1086));
  OAI211_X1 g661(.A(G40), .B(G160), .C1(new_n1086), .C2(new_n1065), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1087), .B1(new_n1065), .B2(new_n1060), .ZN(new_n1088));
  INV_X1    g663(.A(G1971), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1086), .A2(KEYINPUT45), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1040), .B(new_n1090), .C1(new_n1060), .C2(KEYINPUT45), .ZN(new_n1091));
  AOI22_X1  g666(.A1(new_n1088), .A2(new_n816), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1085), .B1(new_n1092), .B2(new_n1079), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1091), .A2(new_n1089), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1067), .B(new_n816), .C1(new_n1060), .C2(new_n1065), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1079), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1040), .A2(new_n1086), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n587), .A2(G1976), .A3(new_n589), .ZN(new_n1099));
  AOI21_X1  g674(.A(KEYINPUT52), .B1(G288), .B2(new_n712), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1098), .A2(G8), .A3(new_n1099), .A4(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(G160), .A2(G40), .ZN(new_n1102));
  OAI211_X1 g677(.A(G8), .B(new_n1099), .C1(new_n1102), .C2(new_n1043), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT52), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n530), .A2(G48), .ZN(new_n1106));
  INV_X1    g681(.A(G86), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1106), .B(new_n594), .C1(new_n600), .C2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(G1981), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1109), .A2(KEYINPUT120), .ZN(new_n1110));
  AND2_X1   g685(.A1(new_n1109), .A2(KEYINPUT120), .ZN(new_n1111));
  INV_X1    g686(.A(G1981), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n595), .A2(new_n596), .A3(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1110), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT49), .ZN(new_n1115));
  OR2_X1    g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1098), .A2(G8), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1117), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1105), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1093), .A2(new_n1097), .A3(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n515), .A2(new_n1042), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(new_n1041), .ZN(new_n1122));
  INV_X1    g697(.A(G2078), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1122), .A2(new_n1123), .A3(new_n1040), .A4(new_n1090), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT53), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1067), .B1(new_n1060), .B2(new_n1065), .ZN(new_n1126));
  AOI22_X1  g701(.A1(new_n1124), .A2(new_n1125), .B1(new_n1126), .B2(new_n836), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1102), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1128), .B(new_n1123), .C1(new_n1041), .C2(new_n1121), .ZN(new_n1129));
  AND2_X1   g704(.A1(new_n1129), .A2(KEYINPUT124), .ZN(new_n1130));
  OAI21_X1  g705(.A(KEYINPUT53), .B1(new_n1129), .B2(KEYINPUT124), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1127), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(G171), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1120), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1076), .A2(new_n1078), .A3(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1113), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1137));
  NOR2_X1   g712(.A1(G288), .A2(G1976), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1136), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1119), .ZN(new_n1140));
  OAI22_X1  g715(.A1(new_n1139), .A2(new_n1117), .B1(new_n1140), .B2(new_n1097), .ZN(new_n1141));
  NAND2_X1  g716(.A1(G168), .A2(G8), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1142), .B1(new_n1064), .B2(new_n1068), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1093), .A2(new_n1097), .A3(new_n1119), .A4(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT63), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  OR3_X1    g721(.A1(new_n1096), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1147));
  AND2_X1   g722(.A1(new_n1143), .A2(KEYINPUT63), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1147), .A2(new_n1097), .A3(new_n1148), .A4(new_n1119), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1141), .B1(new_n1146), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1135), .A2(new_n1150), .ZN(new_n1151));
  XOR2_X1   g726(.A(KEYINPUT56), .B(G2072), .Z(new_n1152));
  OR2_X1    g727(.A1(new_n1091), .A2(new_n1152), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1121), .A2(KEYINPUT50), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n826), .B1(new_n1154), .B2(new_n1087), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n617), .B(KEYINPUT57), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1153), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  XOR2_X1   g732(.A(new_n1157), .B(KEYINPUT121), .Z(new_n1158));
  NAND2_X1  g733(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1156), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(new_n611), .ZN(new_n1162));
  INV_X1    g737(.A(G1348), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1098), .ZN(new_n1164));
  AOI22_X1  g739(.A1(new_n1163), .A2(new_n1126), .B1(new_n1164), .B2(new_n873), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1161), .B1(new_n1162), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1158), .A2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(KEYINPUT61), .B1(new_n1158), .B2(new_n1161), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1165), .A2(KEYINPUT60), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(KEYINPUT123), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT123), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1165), .A2(new_n1171), .A3(KEYINPUT60), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n611), .B1(new_n1165), .B2(KEYINPUT60), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  XNOR2_X1  g750(.A(KEYINPUT58), .B(G1341), .ZN(new_n1176));
  OAI22_X1  g751(.A1(new_n1091), .A2(G1996), .B1(new_n1164), .B2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1177), .A2(KEYINPUT122), .A3(new_n568), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n1178), .B(KEYINPUT59), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1174), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1180), .A2(new_n1170), .A3(new_n1172), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1161), .A2(KEYINPUT61), .A3(new_n1157), .ZN(new_n1182));
  NAND4_X1  g757(.A1(new_n1175), .A2(new_n1179), .A3(new_n1181), .A4(new_n1182), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1167), .B1(new_n1168), .B2(new_n1183), .ZN(new_n1184));
  AND2_X1   g759(.A1(new_n1097), .A2(new_n1119), .ZN(new_n1185));
  XNOR2_X1  g760(.A(G301), .B(KEYINPUT54), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1132), .A2(new_n1186), .ZN(new_n1187));
  AOI211_X1 g762(.A(new_n1125), .B(G2078), .C1(new_n1086), .C2(KEYINPUT45), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1186), .B1(new_n1128), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1127), .A2(new_n1189), .ZN(new_n1190));
  NAND4_X1  g765(.A1(new_n1185), .A2(new_n1187), .A3(new_n1093), .A4(new_n1190), .ZN(new_n1191));
  AND2_X1   g766(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1192));
  OAI21_X1  g767(.A(KEYINPUT125), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  AND4_X1   g768(.A1(new_n1093), .A2(new_n1190), .A3(new_n1097), .A4(new_n1119), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT125), .ZN(new_n1195));
  NAND4_X1  g770(.A1(new_n1194), .A2(new_n1075), .A3(new_n1195), .A4(new_n1187), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1193), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1151), .B1(new_n1184), .B2(new_n1197), .ZN(new_n1198));
  AND2_X1   g773(.A1(new_n1036), .A2(new_n1053), .ZN(new_n1199));
  XOR2_X1   g774(.A(G290), .B(G1986), .Z(new_n1200));
  AOI21_X1  g775(.A(new_n1044), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1058), .B1(new_n1198), .B2(new_n1201), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g777(.A(new_n667), .ZN(new_n1204));
  OR4_X1    g778(.A1(new_n461), .A2(G229), .A3(new_n1204), .A4(G227), .ZN(new_n1205));
  AOI21_X1  g779(.A(new_n1205), .B1(new_n961), .B2(new_n964), .ZN(new_n1206));
  AND2_X1   g780(.A1(new_n1206), .A2(new_n1027), .ZN(G308));
  NAND2_X1  g781(.A1(new_n1206), .A2(new_n1027), .ZN(G225));
endmodule


