

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588;

  NOR2_X1 U324 ( .A1(n531), .A2(n461), .ZN(n575) );
  XOR2_X1 U325 ( .A(G50GAT), .B(G36GAT), .Z(n292) );
  XNOR2_X1 U326 ( .A(n390), .B(n292), .ZN(n296) );
  XNOR2_X1 U327 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U328 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U329 ( .A(n340), .B(n339), .ZN(n344) );
  XNOR2_X1 U330 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U331 ( .A(n305), .B(n304), .ZN(n310) );
  INV_X1 U332 ( .A(G218GAT), .ZN(n454) );
  NOR2_X1 U333 ( .A1(n452), .A2(n469), .ZN(n586) );
  XNOR2_X1 U334 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U335 ( .A(n466), .B(G190GAT), .ZN(n467) );
  XNOR2_X1 U336 ( .A(n457), .B(n456), .ZN(G1355GAT) );
  XNOR2_X1 U337 ( .A(n468), .B(n467), .ZN(G1351GAT) );
  XOR2_X1 U338 ( .A(G190GAT), .B(KEYINPUT80), .Z(n390) );
  XOR2_X1 U339 ( .A(G92GAT), .B(G106GAT), .Z(n294) );
  XNOR2_X1 U340 ( .A(G218GAT), .B(G162GAT), .ZN(n293) );
  XNOR2_X1 U341 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U342 ( .A(G99GAT), .B(G85GAT), .Z(n333) );
  XOR2_X1 U343 ( .A(n297), .B(n333), .Z(n305) );
  XOR2_X1 U344 ( .A(G29GAT), .B(G43GAT), .Z(n299) );
  XNOR2_X1 U345 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n298) );
  XNOR2_X1 U346 ( .A(n299), .B(n298), .ZN(n324) );
  XOR2_X1 U347 ( .A(G134GAT), .B(KEYINPUT78), .Z(n409) );
  XNOR2_X1 U348 ( .A(n324), .B(n409), .ZN(n303) );
  XOR2_X1 U349 ( .A(KEYINPUT11), .B(KEYINPUT77), .Z(n301) );
  NAND2_X1 U350 ( .A1(G232GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U351 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U352 ( .A(KEYINPUT67), .B(KEYINPUT9), .Z(n307) );
  XNOR2_X1 U353 ( .A(KEYINPUT65), .B(KEYINPUT79), .ZN(n306) );
  XNOR2_X1 U354 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U355 ( .A(n308), .B(KEYINPUT10), .ZN(n309) );
  XNOR2_X1 U356 ( .A(n310), .B(n309), .ZN(n552) );
  XOR2_X1 U357 ( .A(n552), .B(KEYINPUT101), .Z(n311) );
  XNOR2_X1 U358 ( .A(n311), .B(KEYINPUT36), .ZN(n496) );
  XOR2_X1 U359 ( .A(KEYINPUT68), .B(KEYINPUT70), .Z(n313) );
  NAND2_X1 U360 ( .A1(G229GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U361 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U362 ( .A(n314), .B(KEYINPUT29), .Z(n318) );
  XNOR2_X1 U363 ( .A(G169GAT), .B(G36GAT), .ZN(n315) );
  XNOR2_X1 U364 ( .A(n315), .B(G8GAT), .ZN(n380) );
  XNOR2_X1 U365 ( .A(G15GAT), .B(G1GAT), .ZN(n316) );
  XNOR2_X1 U366 ( .A(n316), .B(KEYINPUT71), .ZN(n356) );
  XNOR2_X1 U367 ( .A(n380), .B(n356), .ZN(n317) );
  XNOR2_X1 U368 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U369 ( .A(KEYINPUT30), .B(KEYINPUT69), .Z(n320) );
  XNOR2_X1 U370 ( .A(G197GAT), .B(G113GAT), .ZN(n319) );
  XNOR2_X1 U371 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U372 ( .A(n322), .B(n321), .Z(n326) );
  XNOR2_X1 U373 ( .A(G50GAT), .B(G22GAT), .ZN(n323) );
  XNOR2_X1 U374 ( .A(n323), .B(G141GAT), .ZN(n429) );
  XNOR2_X1 U375 ( .A(n324), .B(n429), .ZN(n325) );
  XNOR2_X1 U376 ( .A(n326), .B(n325), .ZN(n577) );
  INV_X1 U377 ( .A(G92GAT), .ZN(n327) );
  NAND2_X1 U378 ( .A1(G64GAT), .A2(n327), .ZN(n330) );
  INV_X1 U379 ( .A(G64GAT), .ZN(n328) );
  NAND2_X1 U380 ( .A1(n328), .A2(G92GAT), .ZN(n329) );
  NAND2_X1 U381 ( .A1(n330), .A2(n329), .ZN(n332) );
  XNOR2_X1 U382 ( .A(G176GAT), .B(G204GAT), .ZN(n331) );
  XNOR2_X1 U383 ( .A(n332), .B(n331), .ZN(n381) );
  XNOR2_X1 U384 ( .A(n381), .B(n333), .ZN(n335) );
  AND2_X1 U385 ( .A1(G230GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U386 ( .A(n335), .B(n334), .ZN(n340) );
  XNOR2_X1 U387 ( .A(G106GAT), .B(G78GAT), .ZN(n336) );
  XNOR2_X1 U388 ( .A(n336), .B(G148GAT), .ZN(n426) );
  XNOR2_X1 U389 ( .A(n426), .B(KEYINPUT75), .ZN(n338) );
  INV_X1 U390 ( .A(KEYINPUT74), .ZN(n337) );
  XOR2_X1 U391 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n342) );
  XNOR2_X1 U392 ( .A(KEYINPUT31), .B(KEYINPUT73), .ZN(n341) );
  XOR2_X1 U393 ( .A(n342), .B(n341), .Z(n343) );
  XNOR2_X1 U394 ( .A(n344), .B(n343), .ZN(n346) );
  XOR2_X1 U395 ( .A(G120GAT), .B(G71GAT), .Z(n435) );
  XOR2_X1 U396 ( .A(G57GAT), .B(KEYINPUT13), .Z(n352) );
  XNOR2_X1 U397 ( .A(n435), .B(n352), .ZN(n345) );
  XNOR2_X1 U398 ( .A(n346), .B(n345), .ZN(n582) );
  INV_X1 U399 ( .A(KEYINPUT64), .ZN(n347) );
  XNOR2_X1 U400 ( .A(n582), .B(n347), .ZN(n348) );
  XOR2_X1 U401 ( .A(KEYINPUT41), .B(n348), .Z(n543) );
  INV_X1 U402 ( .A(n543), .ZN(n564) );
  NAND2_X1 U403 ( .A1(n577), .A2(n564), .ZN(n349) );
  XNOR2_X1 U404 ( .A(n349), .B(KEYINPUT46), .ZN(n370) );
  INV_X1 U405 ( .A(n552), .ZN(n568) );
  XOR2_X1 U406 ( .A(G155GAT), .B(G211GAT), .Z(n351) );
  XNOR2_X1 U407 ( .A(G127GAT), .B(G183GAT), .ZN(n350) );
  XNOR2_X1 U408 ( .A(n351), .B(n350), .ZN(n353) );
  XOR2_X1 U409 ( .A(n353), .B(n352), .Z(n355) );
  XNOR2_X1 U410 ( .A(G22GAT), .B(G78GAT), .ZN(n354) );
  XNOR2_X1 U411 ( .A(n355), .B(n354), .ZN(n360) );
  XOR2_X1 U412 ( .A(n356), .B(KEYINPUT12), .Z(n358) );
  NAND2_X1 U413 ( .A1(G231GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U414 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U415 ( .A(n360), .B(n359), .Z(n368) );
  XOR2_X1 U416 ( .A(KEYINPUT83), .B(G64GAT), .Z(n362) );
  XNOR2_X1 U417 ( .A(G8GAT), .B(G71GAT), .ZN(n361) );
  XNOR2_X1 U418 ( .A(n362), .B(n361), .ZN(n366) );
  XOR2_X1 U419 ( .A(KEYINPUT82), .B(KEYINPUT81), .Z(n364) );
  XNOR2_X1 U420 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n363) );
  XNOR2_X1 U421 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U422 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U423 ( .A(n368), .B(n367), .Z(n587) );
  NOR2_X1 U424 ( .A1(n568), .A2(n587), .ZN(n369) );
  AND2_X1 U425 ( .A1(n370), .A2(n369), .ZN(n371) );
  XOR2_X1 U426 ( .A(KEYINPUT47), .B(n371), .Z(n378) );
  INV_X1 U427 ( .A(n587), .ZN(n548) );
  NOR2_X1 U428 ( .A1(n496), .A2(n548), .ZN(n373) );
  XNOR2_X1 U429 ( .A(KEYINPUT66), .B(KEYINPUT45), .ZN(n372) );
  XNOR2_X1 U430 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U431 ( .A(n577), .B(KEYINPUT72), .Z(n571) );
  NAND2_X1 U432 ( .A1(n374), .A2(n571), .ZN(n375) );
  NOR2_X1 U433 ( .A1(n582), .A2(n375), .ZN(n376) );
  XNOR2_X1 U434 ( .A(KEYINPUT114), .B(n376), .ZN(n377) );
  NOR2_X1 U435 ( .A1(n378), .A2(n377), .ZN(n379) );
  XNOR2_X1 U436 ( .A(KEYINPUT48), .B(n379), .ZN(n559) );
  XNOR2_X1 U437 ( .A(n381), .B(n380), .ZN(n394) );
  XOR2_X1 U438 ( .A(KEYINPUT95), .B(KEYINPUT94), .Z(n388) );
  XOR2_X1 U439 ( .A(G183GAT), .B(KEYINPUT17), .Z(n383) );
  XNOR2_X1 U440 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n382) );
  XNOR2_X1 U441 ( .A(n383), .B(n382), .ZN(n444) );
  XOR2_X1 U442 ( .A(KEYINPUT90), .B(G218GAT), .Z(n385) );
  XNOR2_X1 U443 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n384) );
  XNOR2_X1 U444 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U445 ( .A(G197GAT), .B(n386), .Z(n428) );
  XNOR2_X1 U446 ( .A(n444), .B(n428), .ZN(n387) );
  XNOR2_X1 U447 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U448 ( .A(n390), .B(n389), .Z(n392) );
  NAND2_X1 U449 ( .A1(G226GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U450 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U451 ( .A(n394), .B(n393), .Z(n528) );
  XNOR2_X1 U452 ( .A(KEYINPUT120), .B(n528), .ZN(n395) );
  NOR2_X1 U453 ( .A1(n559), .A2(n395), .ZN(n396) );
  XNOR2_X1 U454 ( .A(KEYINPUT54), .B(n396), .ZN(n459) );
  XOR2_X1 U455 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n398) );
  XNOR2_X1 U456 ( .A(KEYINPUT93), .B(KEYINPUT1), .ZN(n397) );
  XNOR2_X1 U457 ( .A(n398), .B(n397), .ZN(n416) );
  XOR2_X1 U458 ( .A(G85GAT), .B(G148GAT), .Z(n400) );
  XNOR2_X1 U459 ( .A(G29GAT), .B(G141GAT), .ZN(n399) );
  XNOR2_X1 U460 ( .A(n400), .B(n399), .ZN(n404) );
  XOR2_X1 U461 ( .A(KEYINPUT6), .B(G57GAT), .Z(n402) );
  XNOR2_X1 U462 ( .A(G1GAT), .B(G120GAT), .ZN(n401) );
  XNOR2_X1 U463 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U464 ( .A(n404), .B(n403), .Z(n414) );
  XOR2_X1 U465 ( .A(KEYINPUT91), .B(G162GAT), .Z(n406) );
  XNOR2_X1 U466 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n405) );
  XNOR2_X1 U467 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U468 ( .A(KEYINPUT3), .B(n407), .Z(n423) );
  XNOR2_X1 U469 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n408) );
  XNOR2_X1 U470 ( .A(n408), .B(G127GAT), .ZN(n445) );
  XOR2_X1 U471 ( .A(n409), .B(n445), .Z(n411) );
  NAND2_X1 U472 ( .A1(G225GAT), .A2(G233GAT), .ZN(n410) );
  XNOR2_X1 U473 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U474 ( .A(n423), .B(n412), .ZN(n413) );
  XNOR2_X1 U475 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U476 ( .A(n416), .B(n415), .ZN(n556) );
  INV_X1 U477 ( .A(n556), .ZN(n526) );
  NAND2_X1 U478 ( .A1(n459), .A2(n526), .ZN(n452) );
  XOR2_X1 U479 ( .A(KEYINPUT89), .B(KEYINPUT22), .Z(n418) );
  XNOR2_X1 U480 ( .A(KEYINPUT24), .B(KEYINPUT88), .ZN(n417) );
  XNOR2_X1 U481 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U482 ( .A(G204GAT), .B(n419), .Z(n421) );
  NAND2_X1 U483 ( .A1(G228GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U484 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U485 ( .A(n422), .B(KEYINPUT92), .Z(n425) );
  XNOR2_X1 U486 ( .A(n423), .B(KEYINPUT23), .ZN(n424) );
  XNOR2_X1 U487 ( .A(n425), .B(n424), .ZN(n427) );
  XOR2_X1 U488 ( .A(n427), .B(n426), .Z(n431) );
  XNOR2_X1 U489 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U490 ( .A(n431), .B(n430), .ZN(n475) );
  XOR2_X1 U491 ( .A(G190GAT), .B(G99GAT), .Z(n433) );
  XNOR2_X1 U492 ( .A(G43GAT), .B(G134GAT), .ZN(n432) );
  XNOR2_X1 U493 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U494 ( .A(n435), .B(n434), .Z(n437) );
  NAND2_X1 U495 ( .A1(G227GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U496 ( .A(n437), .B(n436), .ZN(n449) );
  XOR2_X1 U497 ( .A(KEYINPUT85), .B(G176GAT), .Z(n439) );
  XNOR2_X1 U498 ( .A(KEYINPUT20), .B(KEYINPUT87), .ZN(n438) );
  XNOR2_X1 U499 ( .A(n439), .B(n438), .ZN(n443) );
  XOR2_X1 U500 ( .A(KEYINPUT84), .B(KEYINPUT86), .Z(n441) );
  XNOR2_X1 U501 ( .A(G169GAT), .B(G15GAT), .ZN(n440) );
  XNOR2_X1 U502 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U503 ( .A(n443), .B(n442), .Z(n447) );
  XNOR2_X1 U504 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U505 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U506 ( .A(n449), .B(n448), .ZN(n540) );
  INV_X1 U507 ( .A(n540), .ZN(n531) );
  NAND2_X1 U508 ( .A1(n475), .A2(n531), .ZN(n450) );
  XNOR2_X1 U509 ( .A(n450), .B(KEYINPUT96), .ZN(n451) );
  XNOR2_X1 U510 ( .A(KEYINPUT26), .B(n451), .ZN(n469) );
  INV_X1 U511 ( .A(n586), .ZN(n453) );
  NOR2_X1 U512 ( .A1(n496), .A2(n453), .ZN(n457) );
  XNOR2_X1 U513 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n455) );
  NOR2_X1 U514 ( .A1(n556), .A2(n475), .ZN(n458) );
  AND2_X1 U515 ( .A1(n459), .A2(n458), .ZN(n460) );
  XNOR2_X1 U516 ( .A(n460), .B(KEYINPUT55), .ZN(n461) );
  NAND2_X1 U517 ( .A1(n575), .A2(n564), .ZN(n465) );
  XOR2_X1 U518 ( .A(KEYINPUT122), .B(KEYINPUT56), .Z(n463) );
  XNOR2_X1 U519 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n462) );
  XNOR2_X1 U520 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U521 ( .A(n465), .B(n464), .ZN(G1349GAT) );
  NAND2_X1 U522 ( .A1(n575), .A2(n568), .ZN(n468) );
  XOR2_X1 U523 ( .A(KEYINPUT58), .B(KEYINPUT123), .Z(n466) );
  XOR2_X1 U524 ( .A(n528), .B(KEYINPUT27), .Z(n476) );
  INV_X1 U525 ( .A(n476), .ZN(n470) );
  NOR2_X1 U526 ( .A1(n470), .A2(n469), .ZN(n557) );
  NOR2_X1 U527 ( .A1(n531), .A2(n528), .ZN(n471) );
  NOR2_X1 U528 ( .A1(n475), .A2(n471), .ZN(n472) );
  XOR2_X1 U529 ( .A(KEYINPUT25), .B(n472), .Z(n473) );
  NOR2_X1 U530 ( .A1(n557), .A2(n473), .ZN(n474) );
  NOR2_X1 U531 ( .A1(n474), .A2(n556), .ZN(n479) );
  XOR2_X1 U532 ( .A(n475), .B(KEYINPUT28), .Z(n535) );
  AND2_X1 U533 ( .A1(n556), .A2(n535), .ZN(n477) );
  NAND2_X1 U534 ( .A1(n477), .A2(n476), .ZN(n539) );
  NOR2_X1 U535 ( .A1(n539), .A2(n540), .ZN(n478) );
  NOR2_X1 U536 ( .A1(n479), .A2(n478), .ZN(n495) );
  NOR2_X1 U537 ( .A1(n568), .A2(n548), .ZN(n480) );
  XOR2_X1 U538 ( .A(KEYINPUT16), .B(n480), .Z(n481) );
  NOR2_X1 U539 ( .A1(n495), .A2(n481), .ZN(n510) );
  NOR2_X1 U540 ( .A1(n582), .A2(n571), .ZN(n482) );
  XNOR2_X1 U541 ( .A(n482), .B(KEYINPUT76), .ZN(n499) );
  NAND2_X1 U542 ( .A1(n510), .A2(n499), .ZN(n491) );
  NOR2_X1 U543 ( .A1(n526), .A2(n491), .ZN(n484) );
  XNOR2_X1 U544 ( .A(KEYINPUT34), .B(KEYINPUT97), .ZN(n483) );
  XNOR2_X1 U545 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U546 ( .A(G1GAT), .B(n485), .ZN(G1324GAT) );
  NOR2_X1 U547 ( .A1(n528), .A2(n491), .ZN(n486) );
  XOR2_X1 U548 ( .A(KEYINPUT98), .B(n486), .Z(n487) );
  XNOR2_X1 U549 ( .A(G8GAT), .B(n487), .ZN(G1325GAT) );
  NOR2_X1 U550 ( .A1(n531), .A2(n491), .ZN(n489) );
  XNOR2_X1 U551 ( .A(KEYINPUT35), .B(KEYINPUT99), .ZN(n488) );
  XNOR2_X1 U552 ( .A(n489), .B(n488), .ZN(n490) );
  XOR2_X1 U553 ( .A(G15GAT), .B(n490), .Z(G1326GAT) );
  NOR2_X1 U554 ( .A1(n535), .A2(n491), .ZN(n492) );
  XOR2_X1 U555 ( .A(G22GAT), .B(n492), .Z(G1327GAT) );
  XOR2_X1 U556 ( .A(KEYINPUT102), .B(KEYINPUT39), .Z(n494) );
  XNOR2_X1 U557 ( .A(G29GAT), .B(KEYINPUT100), .ZN(n493) );
  XNOR2_X1 U558 ( .A(n494), .B(n493), .ZN(n502) );
  NOR2_X1 U559 ( .A1(n496), .A2(n495), .ZN(n497) );
  NAND2_X1 U560 ( .A1(n548), .A2(n497), .ZN(n498) );
  XNOR2_X1 U561 ( .A(KEYINPUT37), .B(n498), .ZN(n525) );
  NAND2_X1 U562 ( .A1(n499), .A2(n525), .ZN(n500) );
  XNOR2_X1 U563 ( .A(n500), .B(KEYINPUT38), .ZN(n508) );
  NOR2_X1 U564 ( .A1(n526), .A2(n508), .ZN(n501) );
  XOR2_X1 U565 ( .A(n502), .B(n501), .Z(G1328GAT) );
  NOR2_X1 U566 ( .A1(n508), .A2(n528), .ZN(n503) );
  XOR2_X1 U567 ( .A(G36GAT), .B(n503), .Z(G1329GAT) );
  XOR2_X1 U568 ( .A(KEYINPUT40), .B(KEYINPUT104), .Z(n505) );
  XNOR2_X1 U569 ( .A(G43GAT), .B(KEYINPUT103), .ZN(n504) );
  XNOR2_X1 U570 ( .A(n505), .B(n504), .ZN(n507) );
  NOR2_X1 U571 ( .A1(n531), .A2(n508), .ZN(n506) );
  XOR2_X1 U572 ( .A(n507), .B(n506), .Z(G1330GAT) );
  NOR2_X1 U573 ( .A1(n535), .A2(n508), .ZN(n509) );
  XOR2_X1 U574 ( .A(G50GAT), .B(n509), .Z(G1331GAT) );
  NOR2_X1 U575 ( .A1(n577), .A2(n543), .ZN(n524) );
  NAND2_X1 U576 ( .A1(n524), .A2(n510), .ZN(n511) );
  XOR2_X1 U577 ( .A(KEYINPUT105), .B(n511), .Z(n521) );
  NOR2_X1 U578 ( .A1(n526), .A2(n521), .ZN(n513) );
  XNOR2_X1 U579 ( .A(KEYINPUT42), .B(KEYINPUT106), .ZN(n512) );
  XNOR2_X1 U580 ( .A(n513), .B(n512), .ZN(n514) );
  XOR2_X1 U581 ( .A(G57GAT), .B(n514), .Z(G1332GAT) );
  NOR2_X1 U582 ( .A1(n528), .A2(n521), .ZN(n516) );
  XNOR2_X1 U583 ( .A(KEYINPUT107), .B(KEYINPUT108), .ZN(n515) );
  XNOR2_X1 U584 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U585 ( .A(G64GAT), .B(n517), .ZN(G1333GAT) );
  NOR2_X1 U586 ( .A1(n531), .A2(n521), .ZN(n519) );
  XNOR2_X1 U587 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n518) );
  XNOR2_X1 U588 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U589 ( .A(G71GAT), .B(n520), .ZN(G1334GAT) );
  NOR2_X1 U590 ( .A1(n535), .A2(n521), .ZN(n523) );
  XNOR2_X1 U591 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n522) );
  XNOR2_X1 U592 ( .A(n523), .B(n522), .ZN(G1335GAT) );
  NAND2_X1 U593 ( .A1(n525), .A2(n524), .ZN(n534) );
  NOR2_X1 U594 ( .A1(n526), .A2(n534), .ZN(n527) );
  XOR2_X1 U595 ( .A(G85GAT), .B(n527), .Z(G1336GAT) );
  NOR2_X1 U596 ( .A1(n528), .A2(n534), .ZN(n530) );
  XNOR2_X1 U597 ( .A(G92GAT), .B(KEYINPUT111), .ZN(n529) );
  XNOR2_X1 U598 ( .A(n530), .B(n529), .ZN(G1337GAT) );
  NOR2_X1 U599 ( .A1(n531), .A2(n534), .ZN(n532) );
  XOR2_X1 U600 ( .A(KEYINPUT112), .B(n532), .Z(n533) );
  XNOR2_X1 U601 ( .A(G99GAT), .B(n533), .ZN(G1338GAT) );
  NOR2_X1 U602 ( .A1(n535), .A2(n534), .ZN(n537) );
  XNOR2_X1 U603 ( .A(KEYINPUT44), .B(KEYINPUT113), .ZN(n536) );
  XNOR2_X1 U604 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U605 ( .A(G106GAT), .B(n538), .ZN(G1339GAT) );
  NOR2_X1 U606 ( .A1(n559), .A2(n539), .ZN(n541) );
  NAND2_X1 U607 ( .A1(n541), .A2(n540), .ZN(n551) );
  NOR2_X1 U608 ( .A1(n571), .A2(n551), .ZN(n542) );
  XOR2_X1 U609 ( .A(G113GAT), .B(n542), .Z(G1340GAT) );
  NOR2_X1 U610 ( .A1(n551), .A2(n543), .ZN(n547) );
  XOR2_X1 U611 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n545) );
  XNOR2_X1 U612 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n544) );
  XNOR2_X1 U613 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U614 ( .A(n547), .B(n546), .ZN(G1341GAT) );
  NOR2_X1 U615 ( .A1(n548), .A2(n551), .ZN(n549) );
  XOR2_X1 U616 ( .A(KEYINPUT50), .B(n549), .Z(n550) );
  XNOR2_X1 U617 ( .A(G127GAT), .B(n550), .ZN(G1342GAT) );
  NOR2_X1 U618 ( .A1(n552), .A2(n551), .ZN(n554) );
  XNOR2_X1 U619 ( .A(KEYINPUT51), .B(KEYINPUT117), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n554), .B(n553), .ZN(n555) );
  XOR2_X1 U621 ( .A(G134GAT), .B(n555), .Z(G1343GAT) );
  NAND2_X1 U622 ( .A1(n557), .A2(n556), .ZN(n558) );
  NOR2_X1 U623 ( .A1(n559), .A2(n558), .ZN(n569) );
  NAND2_X1 U624 ( .A1(n569), .A2(n577), .ZN(n560) );
  XNOR2_X1 U625 ( .A(n560), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U626 ( .A(KEYINPUT53), .B(KEYINPUT119), .Z(n562) );
  XNOR2_X1 U627 ( .A(G148GAT), .B(KEYINPUT118), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(n563) );
  XOR2_X1 U629 ( .A(KEYINPUT52), .B(n563), .Z(n566) );
  NAND2_X1 U630 ( .A1(n569), .A2(n564), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n566), .B(n565), .ZN(G1345GAT) );
  NAND2_X1 U632 ( .A1(n587), .A2(n569), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n567), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U635 ( .A(n570), .B(G162GAT), .ZN(G1347GAT) );
  XOR2_X1 U636 ( .A(G169GAT), .B(KEYINPUT121), .Z(n574) );
  INV_X1 U637 ( .A(n571), .ZN(n572) );
  NAND2_X1 U638 ( .A1(n575), .A2(n572), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1348GAT) );
  NAND2_X1 U640 ( .A1(n587), .A2(n575), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n576), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U642 ( .A1(n586), .A2(n577), .ZN(n581) );
  XOR2_X1 U643 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n579) );
  XNOR2_X1 U644 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1352GAT) );
  XOR2_X1 U647 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n584) );
  NAND2_X1 U648 ( .A1(n586), .A2(n582), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(n585) );
  XOR2_X1 U650 ( .A(G204GAT), .B(n585), .Z(G1353GAT) );
  NAND2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U652 ( .A(n588), .B(G211GAT), .ZN(G1354GAT) );
endmodule

