

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U554 ( .A1(n712), .A2(n711), .ZN(n522) );
  INV_X1 U555 ( .A(G168), .ZN(n711) );
  XNOR2_X1 U556 ( .A(KEYINPUT32), .B(KEYINPUT94), .ZN(n733) );
  NAND2_X1 U557 ( .A1(G8), .A2(n719), .ZN(n754) );
  OR2_X1 U558 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U559 ( .A(n664), .B(KEYINPUT15), .ZN(n1018) );
  NOR2_X1 U560 ( .A1(G651), .A2(n603), .ZN(n786) );
  AND2_X1 U561 ( .A1(n546), .A2(n545), .ZN(G160) );
  NOR2_X1 U562 ( .A1(G651), .A2(G543), .ZN(n787) );
  NAND2_X1 U563 ( .A1(n787), .A2(G89), .ZN(n523) );
  XNOR2_X1 U564 ( .A(KEYINPUT4), .B(n523), .ZN(n526) );
  XOR2_X1 U565 ( .A(G543), .B(KEYINPUT0), .Z(n603) );
  XOR2_X1 U566 ( .A(G651), .B(KEYINPUT66), .Z(n528) );
  NOR2_X1 U567 ( .A1(n603), .A2(n528), .ZN(n790) );
  NAND2_X1 U568 ( .A1(G76), .A2(n790), .ZN(n524) );
  XOR2_X1 U569 ( .A(KEYINPUT75), .B(n524), .Z(n525) );
  NAND2_X1 U570 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U571 ( .A(n527), .B(KEYINPUT5), .ZN(n534) );
  NAND2_X1 U572 ( .A1(G51), .A2(n786), .ZN(n531) );
  NOR2_X1 U573 ( .A1(n528), .A2(G543), .ZN(n529) );
  XOR2_X2 U574 ( .A(KEYINPUT1), .B(n529), .Z(n794) );
  NAND2_X1 U575 ( .A1(G63), .A2(n794), .ZN(n530) );
  NAND2_X1 U576 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U577 ( .A(KEYINPUT6), .B(n532), .Z(n533) );
  NAND2_X1 U578 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U579 ( .A(n535), .B(KEYINPUT7), .ZN(G168) );
  AND2_X1 U580 ( .A1(G2105), .A2(G2104), .ZN(n865) );
  NAND2_X1 U581 ( .A1(G113), .A2(n865), .ZN(n538) );
  NOR2_X1 U582 ( .A1(G2105), .A2(G2104), .ZN(n536) );
  XOR2_X2 U583 ( .A(KEYINPUT17), .B(n536), .Z(n870) );
  NAND2_X1 U584 ( .A1(G137), .A2(n870), .ZN(n537) );
  NAND2_X1 U585 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U586 ( .A(KEYINPUT65), .B(n539), .ZN(n546) );
  INV_X1 U587 ( .A(G2105), .ZN(n541) );
  NOR2_X1 U588 ( .A1(G2104), .A2(n541), .ZN(n866) );
  NAND2_X1 U589 ( .A1(G125), .A2(n866), .ZN(n540) );
  XNOR2_X1 U590 ( .A(n540), .B(KEYINPUT64), .ZN(n544) );
  AND2_X1 U591 ( .A1(n541), .A2(G2104), .ZN(n871) );
  NAND2_X1 U592 ( .A1(G101), .A2(n871), .ZN(n542) );
  XOR2_X1 U593 ( .A(KEYINPUT23), .B(n542), .Z(n543) );
  AND2_X1 U594 ( .A1(n544), .A2(n543), .ZN(n545) );
  NAND2_X1 U595 ( .A1(G52), .A2(n786), .ZN(n548) );
  NAND2_X1 U596 ( .A1(G64), .A2(n794), .ZN(n547) );
  NAND2_X1 U597 ( .A1(n548), .A2(n547), .ZN(n553) );
  NAND2_X1 U598 ( .A1(n787), .A2(G90), .ZN(n550) );
  NAND2_X1 U599 ( .A1(G77), .A2(n790), .ZN(n549) );
  NAND2_X1 U600 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U601 ( .A(KEYINPUT9), .B(n551), .Z(n552) );
  NOR2_X1 U602 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U603 ( .A(KEYINPUT69), .B(n554), .Z(G171) );
  INV_X1 U604 ( .A(G171), .ZN(G301) );
  AND2_X1 U605 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U606 ( .A1(G123), .A2(n866), .ZN(n555) );
  XNOR2_X1 U607 ( .A(n555), .B(KEYINPUT18), .ZN(n558) );
  NAND2_X1 U608 ( .A1(G111), .A2(n865), .ZN(n556) );
  XNOR2_X1 U609 ( .A(n556), .B(KEYINPUT76), .ZN(n557) );
  NAND2_X1 U610 ( .A1(n558), .A2(n557), .ZN(n562) );
  NAND2_X1 U611 ( .A1(G135), .A2(n870), .ZN(n560) );
  NAND2_X1 U612 ( .A1(G99), .A2(n871), .ZN(n559) );
  NAND2_X1 U613 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U614 ( .A1(n562), .A2(n561), .ZN(n974) );
  XNOR2_X1 U615 ( .A(n974), .B(G2096), .ZN(n563) );
  XNOR2_X1 U616 ( .A(n563), .B(KEYINPUT77), .ZN(n564) );
  OR2_X1 U617 ( .A1(G2100), .A2(n564), .ZN(G156) );
  INV_X1 U618 ( .A(G57), .ZN(G237) );
  INV_X1 U619 ( .A(G132), .ZN(G219) );
  INV_X1 U620 ( .A(G82), .ZN(G220) );
  NAND2_X1 U621 ( .A1(G138), .A2(n870), .ZN(n566) );
  NAND2_X1 U622 ( .A1(G102), .A2(n871), .ZN(n565) );
  NAND2_X1 U623 ( .A1(n566), .A2(n565), .ZN(n570) );
  NAND2_X1 U624 ( .A1(G114), .A2(n865), .ZN(n568) );
  NAND2_X1 U625 ( .A1(G126), .A2(n866), .ZN(n567) );
  NAND2_X1 U626 ( .A1(n568), .A2(n567), .ZN(n569) );
  NOR2_X1 U627 ( .A1(n570), .A2(n569), .ZN(G164) );
  XOR2_X1 U628 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U629 ( .A1(n794), .A2(G60), .ZN(n571) );
  XNOR2_X1 U630 ( .A(n571), .B(KEYINPUT68), .ZN(n578) );
  NAND2_X1 U631 ( .A1(G47), .A2(n786), .ZN(n573) );
  NAND2_X1 U632 ( .A1(G85), .A2(n787), .ZN(n572) );
  NAND2_X1 U633 ( .A1(n573), .A2(n572), .ZN(n576) );
  NAND2_X1 U634 ( .A1(G72), .A2(n790), .ZN(n574) );
  XNOR2_X1 U635 ( .A(KEYINPUT67), .B(n574), .ZN(n575) );
  NOR2_X1 U636 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U637 ( .A1(n578), .A2(n577), .ZN(G290) );
  NAND2_X1 U638 ( .A1(n787), .A2(G86), .ZN(n580) );
  NAND2_X1 U639 ( .A1(G61), .A2(n794), .ZN(n579) );
  NAND2_X1 U640 ( .A1(n580), .A2(n579), .ZN(n584) );
  NAND2_X1 U641 ( .A1(n790), .A2(G73), .ZN(n581) );
  XNOR2_X1 U642 ( .A(n581), .B(KEYINPUT2), .ZN(n582) );
  XNOR2_X1 U643 ( .A(n582), .B(KEYINPUT79), .ZN(n583) );
  NOR2_X1 U644 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U645 ( .A(n585), .B(KEYINPUT80), .ZN(n587) );
  NAND2_X1 U646 ( .A1(G48), .A2(n786), .ZN(n586) );
  NAND2_X1 U647 ( .A1(n587), .A2(n586), .ZN(G305) );
  NAND2_X1 U648 ( .A1(G65), .A2(n794), .ZN(n594) );
  NAND2_X1 U649 ( .A1(G53), .A2(n786), .ZN(n589) );
  NAND2_X1 U650 ( .A1(G91), .A2(n787), .ZN(n588) );
  NAND2_X1 U651 ( .A1(n589), .A2(n588), .ZN(n592) );
  NAND2_X1 U652 ( .A1(n790), .A2(G78), .ZN(n590) );
  XOR2_X1 U653 ( .A(KEYINPUT70), .B(n590), .Z(n591) );
  NOR2_X1 U654 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U655 ( .A1(n594), .A2(n593), .ZN(n595) );
  XOR2_X1 U656 ( .A(KEYINPUT71), .B(n595), .Z(G299) );
  NAND2_X1 U657 ( .A1(G50), .A2(n786), .ZN(n597) );
  NAND2_X1 U658 ( .A1(G62), .A2(n794), .ZN(n596) );
  NAND2_X1 U659 ( .A1(n597), .A2(n596), .ZN(n601) );
  NAND2_X1 U660 ( .A1(n787), .A2(G88), .ZN(n599) );
  NAND2_X1 U661 ( .A1(G75), .A2(n790), .ZN(n598) );
  NAND2_X1 U662 ( .A1(n599), .A2(n598), .ZN(n600) );
  NOR2_X1 U663 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U664 ( .A(n602), .B(KEYINPUT81), .ZN(G303) );
  NAND2_X1 U665 ( .A1(G87), .A2(n603), .ZN(n605) );
  NAND2_X1 U666 ( .A1(G74), .A2(G651), .ZN(n604) );
  NAND2_X1 U667 ( .A1(n605), .A2(n604), .ZN(n606) );
  NOR2_X1 U668 ( .A1(n794), .A2(n606), .ZN(n608) );
  NAND2_X1 U669 ( .A1(n786), .A2(G49), .ZN(n607) );
  NAND2_X1 U670 ( .A1(n608), .A2(n607), .ZN(G288) );
  INV_X1 U671 ( .A(KEYINPUT40), .ZN(n770) );
  NOR2_X1 U672 ( .A1(G164), .A2(G1384), .ZN(n654) );
  NAND2_X1 U673 ( .A1(G160), .A2(G40), .ZN(n609) );
  NOR2_X1 U674 ( .A1(n654), .A2(n609), .ZN(n650) );
  NAND2_X1 U675 ( .A1(G107), .A2(n865), .ZN(n611) );
  NAND2_X1 U676 ( .A1(G119), .A2(n866), .ZN(n610) );
  NAND2_X1 U677 ( .A1(n611), .A2(n610), .ZN(n615) );
  NAND2_X1 U678 ( .A1(G131), .A2(n870), .ZN(n613) );
  NAND2_X1 U679 ( .A1(G95), .A2(n871), .ZN(n612) );
  NAND2_X1 U680 ( .A1(n613), .A2(n612), .ZN(n614) );
  OR2_X1 U681 ( .A1(n615), .A2(n614), .ZN(n878) );
  NAND2_X1 U682 ( .A1(G1991), .A2(n878), .ZN(n616) );
  XNOR2_X1 U683 ( .A(n616), .B(KEYINPUT86), .ZN(n625) );
  NAND2_X1 U684 ( .A1(G117), .A2(n865), .ZN(n618) );
  NAND2_X1 U685 ( .A1(G129), .A2(n866), .ZN(n617) );
  NAND2_X1 U686 ( .A1(n618), .A2(n617), .ZN(n621) );
  NAND2_X1 U687 ( .A1(n871), .A2(G105), .ZN(n619) );
  XOR2_X1 U688 ( .A(KEYINPUT38), .B(n619), .Z(n620) );
  NOR2_X1 U689 ( .A1(n621), .A2(n620), .ZN(n623) );
  NAND2_X1 U690 ( .A1(n870), .A2(G141), .ZN(n622) );
  NAND2_X1 U691 ( .A1(n623), .A2(n622), .ZN(n886) );
  NAND2_X1 U692 ( .A1(G1996), .A2(n886), .ZN(n624) );
  NAND2_X1 U693 ( .A1(n625), .A2(n624), .ZN(n649) );
  NOR2_X1 U694 ( .A1(G1986), .A2(G290), .ZN(n648) );
  NOR2_X1 U695 ( .A1(G1991), .A2(n878), .ZN(n626) );
  XOR2_X1 U696 ( .A(KEYINPUT99), .B(n626), .Z(n975) );
  NOR2_X1 U697 ( .A1(n648), .A2(n975), .ZN(n627) );
  XNOR2_X1 U698 ( .A(n627), .B(KEYINPUT100), .ZN(n628) );
  NOR2_X1 U699 ( .A1(n649), .A2(n628), .ZN(n630) );
  NOR2_X1 U700 ( .A1(n886), .A2(G1996), .ZN(n629) );
  XNOR2_X1 U701 ( .A(n629), .B(KEYINPUT98), .ZN(n985) );
  NOR2_X1 U702 ( .A1(n630), .A2(n985), .ZN(n631) );
  XNOR2_X1 U703 ( .A(n631), .B(KEYINPUT39), .ZN(n642) );
  XNOR2_X1 U704 ( .A(KEYINPUT37), .B(G2067), .ZN(n643) );
  NAND2_X1 U705 ( .A1(G140), .A2(n870), .ZN(n633) );
  NAND2_X1 U706 ( .A1(G104), .A2(n871), .ZN(n632) );
  NAND2_X1 U707 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U708 ( .A(KEYINPUT34), .B(n634), .ZN(n640) );
  NAND2_X1 U709 ( .A1(n865), .A2(G116), .ZN(n635) );
  XOR2_X1 U710 ( .A(KEYINPUT85), .B(n635), .Z(n637) );
  NAND2_X1 U711 ( .A1(n866), .A2(G128), .ZN(n636) );
  NAND2_X1 U712 ( .A1(n637), .A2(n636), .ZN(n638) );
  XOR2_X1 U713 ( .A(KEYINPUT35), .B(n638), .Z(n639) );
  NOR2_X1 U714 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U715 ( .A(KEYINPUT36), .B(n641), .ZN(n889) );
  NOR2_X1 U716 ( .A1(n643), .A2(n889), .ZN(n980) );
  NAND2_X1 U717 ( .A1(n980), .A2(n650), .ZN(n652) );
  NAND2_X1 U718 ( .A1(n642), .A2(n652), .ZN(n644) );
  NAND2_X1 U719 ( .A1(n643), .A2(n889), .ZN(n991) );
  NAND2_X1 U720 ( .A1(n644), .A2(n991), .ZN(n645) );
  NAND2_X1 U721 ( .A1(n650), .A2(n645), .ZN(n646) );
  XNOR2_X1 U722 ( .A(n646), .B(KEYINPUT101), .ZN(n768) );
  AND2_X1 U723 ( .A1(G290), .A2(G1986), .ZN(n647) );
  NOR2_X1 U724 ( .A1(n648), .A2(n647), .ZN(n1022) );
  INV_X1 U725 ( .A(n649), .ZN(n982) );
  NAND2_X1 U726 ( .A1(n1022), .A2(n982), .ZN(n651) );
  NAND2_X1 U727 ( .A1(n651), .A2(n650), .ZN(n653) );
  NAND2_X1 U728 ( .A1(n653), .A2(n652), .ZN(n766) );
  OR2_X1 U729 ( .A1(G1981), .A2(G305), .ZN(n743) );
  XOR2_X1 U730 ( .A(KEYINPUT24), .B(n743), .Z(n656) );
  AND2_X1 U731 ( .A1(n654), .A2(G40), .ZN(n665) );
  NAND2_X1 U732 ( .A1(G160), .A2(n665), .ZN(n719) );
  INV_X1 U733 ( .A(n754), .ZN(n655) );
  NAND2_X1 U734 ( .A1(n656), .A2(n655), .ZN(n741) );
  NOR2_X1 U735 ( .A1(G2084), .A2(n719), .ZN(n707) );
  NAND2_X1 U736 ( .A1(n707), .A2(G8), .ZN(n718) );
  NOR2_X1 U737 ( .A1(G1966), .A2(n754), .ZN(n716) );
  NAND2_X1 U738 ( .A1(G92), .A2(n787), .ZN(n663) );
  NAND2_X1 U739 ( .A1(n786), .A2(G54), .ZN(n658) );
  NAND2_X1 U740 ( .A1(G79), .A2(n790), .ZN(n657) );
  NAND2_X1 U741 ( .A1(n658), .A2(n657), .ZN(n661) );
  NAND2_X1 U742 ( .A1(n794), .A2(G66), .ZN(n659) );
  XOR2_X1 U743 ( .A(KEYINPUT74), .B(n659), .Z(n660) );
  NOR2_X1 U744 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U745 ( .A1(n663), .A2(n662), .ZN(n664) );
  INV_X1 U746 ( .A(n1018), .ZN(n780) );
  AND2_X1 U747 ( .A1(G160), .A2(n665), .ZN(n701) );
  NOR2_X1 U748 ( .A1(n701), .A2(G1348), .ZN(n667) );
  NOR2_X1 U749 ( .A1(G2067), .A2(n719), .ZN(n666) );
  NOR2_X1 U750 ( .A1(n667), .A2(n666), .ZN(n684) );
  NAND2_X1 U751 ( .A1(n780), .A2(n684), .ZN(n683) );
  NAND2_X1 U752 ( .A1(n787), .A2(G81), .ZN(n668) );
  XNOR2_X1 U753 ( .A(n668), .B(KEYINPUT12), .ZN(n670) );
  NAND2_X1 U754 ( .A1(G68), .A2(n790), .ZN(n669) );
  NAND2_X1 U755 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U756 ( .A(n671), .B(KEYINPUT13), .ZN(n673) );
  NAND2_X1 U757 ( .A1(G43), .A2(n786), .ZN(n672) );
  NAND2_X1 U758 ( .A1(n673), .A2(n672), .ZN(n676) );
  NAND2_X1 U759 ( .A1(n794), .A2(G56), .ZN(n674) );
  XOR2_X1 U760 ( .A(KEYINPUT14), .B(n674), .Z(n675) );
  NOR2_X1 U761 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U762 ( .A(KEYINPUT73), .B(n677), .ZN(n1001) );
  INV_X1 U763 ( .A(G1996), .ZN(n943) );
  NOR2_X1 U764 ( .A1(n719), .A2(n943), .ZN(n678) );
  XOR2_X1 U765 ( .A(n678), .B(KEYINPUT26), .Z(n680) );
  NAND2_X1 U766 ( .A1(n719), .A2(G1341), .ZN(n679) );
  NAND2_X1 U767 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U768 ( .A1(n1001), .A2(n681), .ZN(n682) );
  NAND2_X1 U769 ( .A1(n683), .A2(n682), .ZN(n686) );
  OR2_X1 U770 ( .A1(n684), .A2(n780), .ZN(n685) );
  NAND2_X1 U771 ( .A1(n686), .A2(n685), .ZN(n687) );
  XOR2_X1 U772 ( .A(KEYINPUT90), .B(n687), .Z(n695) );
  INV_X1 U773 ( .A(KEYINPUT88), .ZN(n690) );
  NAND2_X1 U774 ( .A1(G2072), .A2(n701), .ZN(n688) );
  XNOR2_X1 U775 ( .A(KEYINPUT27), .B(n688), .ZN(n689) );
  XNOR2_X1 U776 ( .A(n690), .B(n689), .ZN(n691) );
  XNOR2_X1 U777 ( .A(n691), .B(KEYINPUT87), .ZN(n693) );
  XNOR2_X1 U778 ( .A(G1956), .B(KEYINPUT89), .ZN(n925) );
  NOR2_X1 U779 ( .A1(n925), .A2(n701), .ZN(n692) );
  NOR2_X1 U780 ( .A1(n693), .A2(n692), .ZN(n696) );
  INV_X1 U781 ( .A(G299), .ZN(n1019) );
  NAND2_X1 U782 ( .A1(n696), .A2(n1019), .ZN(n694) );
  NAND2_X1 U783 ( .A1(n695), .A2(n694), .ZN(n699) );
  NOR2_X1 U784 ( .A1(n696), .A2(n1019), .ZN(n697) );
  XOR2_X1 U785 ( .A(n697), .B(KEYINPUT28), .Z(n698) );
  NAND2_X1 U786 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U787 ( .A(n700), .B(KEYINPUT29), .ZN(n705) );
  XOR2_X1 U788 ( .A(G2078), .B(KEYINPUT25), .Z(n944) );
  NOR2_X1 U789 ( .A1(n944), .A2(n719), .ZN(n703) );
  NOR2_X1 U790 ( .A1(n701), .A2(G1961), .ZN(n702) );
  NOR2_X1 U791 ( .A1(n703), .A2(n702), .ZN(n706) );
  NOR2_X1 U792 ( .A1(G301), .A2(n706), .ZN(n704) );
  NOR2_X1 U793 ( .A1(n705), .A2(n704), .ZN(n729) );
  AND2_X1 U794 ( .A1(G301), .A2(n706), .ZN(n713) );
  NOR2_X1 U795 ( .A1(n716), .A2(n707), .ZN(n708) );
  NAND2_X1 U796 ( .A1(G8), .A2(n708), .ZN(n709) );
  XNOR2_X1 U797 ( .A(KEYINPUT91), .B(n709), .ZN(n710) );
  XNOR2_X1 U798 ( .A(n710), .B(KEYINPUT30), .ZN(n712) );
  NOR2_X1 U799 ( .A1(n713), .A2(n522), .ZN(n714) );
  XNOR2_X1 U800 ( .A(n714), .B(KEYINPUT31), .ZN(n727) );
  NOR2_X1 U801 ( .A1(n729), .A2(n727), .ZN(n715) );
  NOR2_X1 U802 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U803 ( .A1(n718), .A2(n717), .ZN(n736) );
  INV_X1 U804 ( .A(G8), .ZN(n726) );
  NOR2_X1 U805 ( .A1(G2090), .A2(n719), .ZN(n720) );
  XNOR2_X1 U806 ( .A(n720), .B(KEYINPUT92), .ZN(n722) );
  NOR2_X1 U807 ( .A1(n754), .A2(G1971), .ZN(n721) );
  NOR2_X1 U808 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U809 ( .A(KEYINPUT93), .B(n723), .Z(n724) );
  NAND2_X1 U810 ( .A1(n724), .A2(G303), .ZN(n725) );
  NOR2_X1 U811 ( .A1(n726), .A2(n725), .ZN(n730) );
  OR2_X1 U812 ( .A1(n727), .A2(n730), .ZN(n728) );
  OR2_X1 U813 ( .A1(n729), .A2(n728), .ZN(n732) );
  OR2_X1 U814 ( .A1(n730), .A2(G286), .ZN(n731) );
  NAND2_X1 U815 ( .A1(n732), .A2(n731), .ZN(n734) );
  XNOR2_X1 U816 ( .A(n734), .B(n733), .ZN(n735) );
  NAND2_X1 U817 ( .A1(n736), .A2(n735), .ZN(n745) );
  NOR2_X1 U818 ( .A1(G2090), .A2(G303), .ZN(n737) );
  NAND2_X1 U819 ( .A1(G8), .A2(n737), .ZN(n738) );
  NAND2_X1 U820 ( .A1(n745), .A2(n738), .ZN(n739) );
  NAND2_X1 U821 ( .A1(n754), .A2(n739), .ZN(n740) );
  NAND2_X1 U822 ( .A1(n741), .A2(n740), .ZN(n764) );
  NAND2_X1 U823 ( .A1(G1981), .A2(G305), .ZN(n742) );
  NAND2_X1 U824 ( .A1(n743), .A2(n742), .ZN(n1012) );
  NOR2_X1 U825 ( .A1(G1976), .A2(G288), .ZN(n744) );
  XNOR2_X1 U826 ( .A(KEYINPUT95), .B(n744), .ZN(n1004) );
  NAND2_X1 U827 ( .A1(n1004), .A2(n745), .ZN(n752) );
  NOR2_X1 U828 ( .A1(G1971), .A2(G303), .ZN(n750) );
  INV_X1 U829 ( .A(KEYINPUT33), .ZN(n748) );
  OR2_X1 U830 ( .A1(n754), .A2(n1004), .ZN(n746) );
  NOR2_X1 U831 ( .A1(n748), .A2(n746), .ZN(n747) );
  XOR2_X1 U832 ( .A(n747), .B(KEYINPUT97), .Z(n756) );
  OR2_X1 U833 ( .A1(n756), .A2(n748), .ZN(n759) );
  INV_X1 U834 ( .A(n759), .ZN(n749) );
  OR2_X1 U835 ( .A1(n750), .A2(n749), .ZN(n751) );
  NOR2_X1 U836 ( .A1(n752), .A2(n751), .ZN(n761) );
  NAND2_X1 U837 ( .A1(G288), .A2(G1976), .ZN(n753) );
  XNOR2_X1 U838 ( .A(n753), .B(KEYINPUT96), .ZN(n1005) );
  INV_X1 U839 ( .A(n1005), .ZN(n755) );
  OR2_X1 U840 ( .A1(n755), .A2(n754), .ZN(n757) );
  OR2_X1 U841 ( .A1(n757), .A2(n756), .ZN(n758) );
  AND2_X1 U842 ( .A1(n759), .A2(n758), .ZN(n760) );
  NOR2_X1 U843 ( .A1(n1012), .A2(n762), .ZN(n763) );
  NOR2_X1 U844 ( .A1(n764), .A2(n763), .ZN(n765) );
  NOR2_X1 U845 ( .A1(n766), .A2(n765), .ZN(n767) );
  NOR2_X1 U846 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U847 ( .A(n770), .B(n769), .ZN(G329) );
  NAND2_X1 U848 ( .A1(G7), .A2(G661), .ZN(n771) );
  XNOR2_X1 U849 ( .A(n771), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U850 ( .A(KEYINPUT11), .B(KEYINPUT72), .Z(n773) );
  INV_X1 U851 ( .A(G223), .ZN(n824) );
  NAND2_X1 U852 ( .A1(G567), .A2(n824), .ZN(n772) );
  XNOR2_X1 U853 ( .A(n773), .B(n772), .ZN(G234) );
  INV_X1 U854 ( .A(G860), .ZN(n785) );
  OR2_X1 U855 ( .A1(n1001), .A2(n785), .ZN(G153) );
  NAND2_X1 U856 ( .A1(G868), .A2(G301), .ZN(n775) );
  INV_X1 U857 ( .A(G868), .ZN(n806) );
  NAND2_X1 U858 ( .A1(n780), .A2(n806), .ZN(n774) );
  NAND2_X1 U859 ( .A1(n775), .A2(n774), .ZN(G284) );
  NAND2_X1 U860 ( .A1(G286), .A2(G868), .ZN(n777) );
  NAND2_X1 U861 ( .A1(G299), .A2(n806), .ZN(n776) );
  NAND2_X1 U862 ( .A1(n777), .A2(n776), .ZN(G297) );
  NAND2_X1 U863 ( .A1(n785), .A2(G559), .ZN(n778) );
  NAND2_X1 U864 ( .A1(n778), .A2(n1018), .ZN(n779) );
  XNOR2_X1 U865 ( .A(n779), .B(KEYINPUT16), .ZN(G148) );
  OR2_X1 U866 ( .A1(G559), .A2(n780), .ZN(n781) );
  NAND2_X1 U867 ( .A1(n781), .A2(G868), .ZN(n783) );
  NAND2_X1 U868 ( .A1(n1001), .A2(n806), .ZN(n782) );
  NAND2_X1 U869 ( .A1(n783), .A2(n782), .ZN(G282) );
  NAND2_X1 U870 ( .A1(G559), .A2(n1018), .ZN(n784) );
  XOR2_X1 U871 ( .A(n1001), .B(n784), .Z(n804) );
  NAND2_X1 U872 ( .A1(n785), .A2(n804), .ZN(n797) );
  NAND2_X1 U873 ( .A1(G55), .A2(n786), .ZN(n789) );
  NAND2_X1 U874 ( .A1(G93), .A2(n787), .ZN(n788) );
  NAND2_X1 U875 ( .A1(n789), .A2(n788), .ZN(n793) );
  NAND2_X1 U876 ( .A1(n790), .A2(G80), .ZN(n791) );
  XOR2_X1 U877 ( .A(KEYINPUT78), .B(n791), .Z(n792) );
  NOR2_X1 U878 ( .A1(n793), .A2(n792), .ZN(n796) );
  NAND2_X1 U879 ( .A1(G67), .A2(n794), .ZN(n795) );
  NAND2_X1 U880 ( .A1(n796), .A2(n795), .ZN(n807) );
  XNOR2_X1 U881 ( .A(n797), .B(n807), .ZN(G145) );
  INV_X1 U882 ( .A(G303), .ZN(G166) );
  XOR2_X1 U883 ( .A(G305), .B(G290), .Z(n799) );
  XNOR2_X1 U884 ( .A(G166), .B(n1019), .ZN(n798) );
  XNOR2_X1 U885 ( .A(n799), .B(n798), .ZN(n800) );
  XNOR2_X1 U886 ( .A(n800), .B(G288), .ZN(n803) );
  XNOR2_X1 U887 ( .A(KEYINPUT19), .B(KEYINPUT82), .ZN(n801) );
  XNOR2_X1 U888 ( .A(n801), .B(n807), .ZN(n802) );
  XNOR2_X1 U889 ( .A(n803), .B(n802), .ZN(n892) );
  XOR2_X1 U890 ( .A(n892), .B(n804), .Z(n805) );
  NOR2_X1 U891 ( .A1(n806), .A2(n805), .ZN(n809) );
  NOR2_X1 U892 ( .A1(G868), .A2(n807), .ZN(n808) );
  NOR2_X1 U893 ( .A1(n809), .A2(n808), .ZN(G295) );
  NAND2_X1 U894 ( .A1(G2078), .A2(G2084), .ZN(n810) );
  XOR2_X1 U895 ( .A(KEYINPUT20), .B(n810), .Z(n811) );
  NAND2_X1 U896 ( .A1(G2090), .A2(n811), .ZN(n812) );
  XNOR2_X1 U897 ( .A(KEYINPUT21), .B(n812), .ZN(n813) );
  NAND2_X1 U898 ( .A1(n813), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U899 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U900 ( .A1(G483), .A2(G661), .ZN(n822) );
  NOR2_X1 U901 ( .A1(G220), .A2(G219), .ZN(n814) );
  XOR2_X1 U902 ( .A(KEYINPUT22), .B(n814), .Z(n815) );
  NOR2_X1 U903 ( .A1(G218), .A2(n815), .ZN(n816) );
  XOR2_X1 U904 ( .A(KEYINPUT83), .B(n816), .Z(n817) );
  NAND2_X1 U905 ( .A1(G96), .A2(n817), .ZN(n828) );
  NAND2_X1 U906 ( .A1(n828), .A2(G2106), .ZN(n821) );
  NAND2_X1 U907 ( .A1(G69), .A2(G120), .ZN(n818) );
  NOR2_X1 U908 ( .A1(G237), .A2(n818), .ZN(n819) );
  NAND2_X1 U909 ( .A1(G108), .A2(n819), .ZN(n829) );
  NAND2_X1 U910 ( .A1(n829), .A2(G567), .ZN(n820) );
  NAND2_X1 U911 ( .A1(n821), .A2(n820), .ZN(n830) );
  NOR2_X1 U912 ( .A1(n822), .A2(n830), .ZN(n823) );
  XNOR2_X1 U913 ( .A(n823), .B(KEYINPUT84), .ZN(n827) );
  NAND2_X1 U914 ( .A1(G36), .A2(n827), .ZN(G176) );
  NAND2_X1 U915 ( .A1(G2106), .A2(n824), .ZN(G217) );
  AND2_X1 U916 ( .A1(G15), .A2(G2), .ZN(n825) );
  NAND2_X1 U917 ( .A1(G661), .A2(n825), .ZN(G259) );
  NAND2_X1 U918 ( .A1(G3), .A2(G1), .ZN(n826) );
  NAND2_X1 U919 ( .A1(n827), .A2(n826), .ZN(G188) );
  INV_X1 U921 ( .A(G120), .ZN(G236) );
  INV_X1 U922 ( .A(G96), .ZN(G221) );
  INV_X1 U923 ( .A(G69), .ZN(G235) );
  NOR2_X1 U924 ( .A1(n829), .A2(n828), .ZN(G325) );
  INV_X1 U925 ( .A(G325), .ZN(G261) );
  INV_X1 U926 ( .A(n830), .ZN(G319) );
  XOR2_X1 U927 ( .A(G2100), .B(G2096), .Z(n832) );
  XNOR2_X1 U928 ( .A(KEYINPUT42), .B(G2678), .ZN(n831) );
  XNOR2_X1 U929 ( .A(n832), .B(n831), .ZN(n836) );
  XOR2_X1 U930 ( .A(KEYINPUT43), .B(G2072), .Z(n834) );
  XNOR2_X1 U931 ( .A(G2067), .B(G2090), .ZN(n833) );
  XNOR2_X1 U932 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U933 ( .A(n836), .B(n835), .Z(n838) );
  XNOR2_X1 U934 ( .A(G2078), .B(G2084), .ZN(n837) );
  XNOR2_X1 U935 ( .A(n838), .B(n837), .ZN(G227) );
  XOR2_X1 U936 ( .A(G1986), .B(G1981), .Z(n840) );
  XNOR2_X1 U937 ( .A(G1961), .B(G1966), .ZN(n839) );
  XNOR2_X1 U938 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U939 ( .A(n841), .B(KEYINPUT41), .Z(n843) );
  XNOR2_X1 U940 ( .A(G1971), .B(G1976), .ZN(n842) );
  XNOR2_X1 U941 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U942 ( .A(G2474), .B(G1991), .Z(n845) );
  XNOR2_X1 U943 ( .A(G1956), .B(G1996), .ZN(n844) );
  XNOR2_X1 U944 ( .A(n845), .B(n844), .ZN(n846) );
  XNOR2_X1 U945 ( .A(n847), .B(n846), .ZN(G229) );
  NAND2_X1 U946 ( .A1(G112), .A2(n865), .ZN(n849) );
  NAND2_X1 U947 ( .A1(G100), .A2(n871), .ZN(n848) );
  NAND2_X1 U948 ( .A1(n849), .A2(n848), .ZN(n857) );
  NAND2_X1 U949 ( .A1(n870), .A2(G136), .ZN(n850) );
  XNOR2_X1 U950 ( .A(KEYINPUT104), .B(n850), .ZN(n854) );
  XOR2_X1 U951 ( .A(KEYINPUT103), .B(KEYINPUT44), .Z(n852) );
  NAND2_X1 U952 ( .A1(G124), .A2(n866), .ZN(n851) );
  XNOR2_X1 U953 ( .A(n852), .B(n851), .ZN(n853) );
  NAND2_X1 U954 ( .A1(n854), .A2(n853), .ZN(n855) );
  XOR2_X1 U955 ( .A(KEYINPUT105), .B(n855), .Z(n856) );
  NOR2_X1 U956 ( .A1(n857), .A2(n856), .ZN(G162) );
  NAND2_X1 U957 ( .A1(G118), .A2(n865), .ZN(n859) );
  NAND2_X1 U958 ( .A1(G130), .A2(n866), .ZN(n858) );
  NAND2_X1 U959 ( .A1(n859), .A2(n858), .ZN(n864) );
  NAND2_X1 U960 ( .A1(G142), .A2(n870), .ZN(n861) );
  NAND2_X1 U961 ( .A1(G106), .A2(n871), .ZN(n860) );
  NAND2_X1 U962 ( .A1(n861), .A2(n860), .ZN(n862) );
  XOR2_X1 U963 ( .A(n862), .B(KEYINPUT45), .Z(n863) );
  NOR2_X1 U964 ( .A1(n864), .A2(n863), .ZN(n877) );
  NAND2_X1 U965 ( .A1(G115), .A2(n865), .ZN(n868) );
  NAND2_X1 U966 ( .A1(G127), .A2(n866), .ZN(n867) );
  NAND2_X1 U967 ( .A1(n868), .A2(n867), .ZN(n869) );
  XNOR2_X1 U968 ( .A(KEYINPUT47), .B(n869), .ZN(n876) );
  NAND2_X1 U969 ( .A1(G139), .A2(n870), .ZN(n873) );
  NAND2_X1 U970 ( .A1(G103), .A2(n871), .ZN(n872) );
  NAND2_X1 U971 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U972 ( .A(KEYINPUT107), .B(n874), .ZN(n875) );
  NAND2_X1 U973 ( .A1(n876), .A2(n875), .ZN(n968) );
  XNOR2_X1 U974 ( .A(n877), .B(n968), .ZN(n885) );
  XNOR2_X1 U975 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n880) );
  XNOR2_X1 U976 ( .A(n878), .B(KEYINPUT106), .ZN(n879) );
  XNOR2_X1 U977 ( .A(n880), .B(n879), .ZN(n881) );
  XOR2_X1 U978 ( .A(n881), .B(n974), .Z(n883) );
  XNOR2_X1 U979 ( .A(G164), .B(G160), .ZN(n882) );
  XNOR2_X1 U980 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U981 ( .A(n885), .B(n884), .ZN(n888) );
  XNOR2_X1 U982 ( .A(n886), .B(G162), .ZN(n887) );
  XNOR2_X1 U983 ( .A(n888), .B(n887), .ZN(n890) );
  XNOR2_X1 U984 ( .A(n890), .B(n889), .ZN(n891) );
  NOR2_X1 U985 ( .A1(G37), .A2(n891), .ZN(G395) );
  XNOR2_X1 U986 ( .A(n1001), .B(n892), .ZN(n894) );
  XNOR2_X1 U987 ( .A(G171), .B(n1018), .ZN(n893) );
  XNOR2_X1 U988 ( .A(n894), .B(n893), .ZN(n895) );
  XOR2_X1 U989 ( .A(G286), .B(n895), .Z(n896) );
  NOR2_X1 U990 ( .A1(G37), .A2(n896), .ZN(n897) );
  XNOR2_X1 U991 ( .A(KEYINPUT108), .B(n897), .ZN(G397) );
  XOR2_X1 U992 ( .A(KEYINPUT102), .B(G2446), .Z(n899) );
  XNOR2_X1 U993 ( .A(G2443), .B(G2454), .ZN(n898) );
  XNOR2_X1 U994 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U995 ( .A(n900), .B(G2451), .Z(n902) );
  XNOR2_X1 U996 ( .A(G1348), .B(G1341), .ZN(n901) );
  XNOR2_X1 U997 ( .A(n902), .B(n901), .ZN(n906) );
  XOR2_X1 U998 ( .A(G2435), .B(G2427), .Z(n904) );
  XNOR2_X1 U999 ( .A(G2430), .B(G2438), .ZN(n903) );
  XNOR2_X1 U1000 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U1001 ( .A(n906), .B(n905), .Z(n907) );
  NAND2_X1 U1002 ( .A1(G14), .A2(n907), .ZN(n914) );
  NAND2_X1 U1003 ( .A1(G319), .A2(n914), .ZN(n911) );
  NOR2_X1 U1004 ( .A1(G227), .A2(G229), .ZN(n908) );
  XOR2_X1 U1005 ( .A(KEYINPUT49), .B(n908), .Z(n909) );
  XNOR2_X1 U1006 ( .A(n909), .B(KEYINPUT109), .ZN(n910) );
  NOR2_X1 U1007 ( .A1(n911), .A2(n910), .ZN(n913) );
  NOR2_X1 U1008 ( .A1(G395), .A2(G397), .ZN(n912) );
  NAND2_X1 U1009 ( .A1(n913), .A2(n912), .ZN(G225) );
  INV_X1 U1010 ( .A(G225), .ZN(G308) );
  INV_X1 U1011 ( .A(G108), .ZN(G238) );
  INV_X1 U1012 ( .A(n914), .ZN(G401) );
  XOR2_X1 U1013 ( .A(G1961), .B(KEYINPUT124), .Z(n915) );
  XNOR2_X1 U1014 ( .A(G5), .B(n915), .ZN(n923) );
  XOR2_X1 U1015 ( .A(G1971), .B(KEYINPUT127), .Z(n916) );
  XNOR2_X1 U1016 ( .A(G22), .B(n916), .ZN(n920) );
  XOR2_X1 U1017 ( .A(G1976), .B(G23), .Z(n918) );
  XOR2_X1 U1018 ( .A(G1986), .B(G24), .Z(n917) );
  NAND2_X1 U1019 ( .A1(n918), .A2(n917), .ZN(n919) );
  NOR2_X1 U1020 ( .A1(n920), .A2(n919), .ZN(n921) );
  XNOR2_X1 U1021 ( .A(n921), .B(KEYINPUT58), .ZN(n922) );
  NAND2_X1 U1022 ( .A1(n923), .A2(n922), .ZN(n938) );
  XNOR2_X1 U1023 ( .A(G1348), .B(KEYINPUT59), .ZN(n924) );
  XNOR2_X1 U1024 ( .A(n924), .B(G4), .ZN(n929) );
  XOR2_X1 U1025 ( .A(n925), .B(G20), .Z(n927) );
  XNOR2_X1 U1026 ( .A(G6), .B(G1981), .ZN(n926) );
  NOR2_X1 U1027 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1028 ( .A1(n929), .A2(n928), .ZN(n932) );
  XOR2_X1 U1029 ( .A(KEYINPUT125), .B(G1341), .Z(n930) );
  XNOR2_X1 U1030 ( .A(G19), .B(n930), .ZN(n931) );
  NOR2_X1 U1031 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1032 ( .A(KEYINPUT60), .B(n933), .Z(n935) );
  XNOR2_X1 U1033 ( .A(G1966), .B(G21), .ZN(n934) );
  NOR2_X1 U1034 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1035 ( .A(KEYINPUT126), .B(n936), .Z(n937) );
  NOR2_X1 U1036 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1037 ( .A(KEYINPUT61), .B(n939), .Z(n940) );
  NOR2_X1 U1038 ( .A1(G16), .A2(n940), .ZN(n967) );
  XNOR2_X1 U1039 ( .A(G2090), .B(G35), .ZN(n957) );
  XNOR2_X1 U1040 ( .A(G1991), .B(G25), .ZN(n941) );
  XNOR2_X1 U1041 ( .A(n941), .B(KEYINPUT117), .ZN(n942) );
  NAND2_X1 U1042 ( .A1(n942), .A2(G28), .ZN(n954) );
  XNOR2_X1 U1043 ( .A(G32), .B(n943), .ZN(n948) );
  XNOR2_X1 U1044 ( .A(n944), .B(G27), .ZN(n946) );
  XNOR2_X1 U1045 ( .A(G2072), .B(G33), .ZN(n945) );
  NOR2_X1 U1046 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1047 ( .A1(n948), .A2(n947), .ZN(n951) );
  XNOR2_X1 U1048 ( .A(KEYINPUT118), .B(G2067), .ZN(n949) );
  XNOR2_X1 U1049 ( .A(G26), .B(n949), .ZN(n950) );
  NOR2_X1 U1050 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1051 ( .A(n952), .B(KEYINPUT119), .ZN(n953) );
  NOR2_X1 U1052 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1053 ( .A(KEYINPUT53), .B(n955), .ZN(n956) );
  NOR2_X1 U1054 ( .A1(n957), .A2(n956), .ZN(n960) );
  XOR2_X1 U1055 ( .A(G2084), .B(G34), .Z(n958) );
  XNOR2_X1 U1056 ( .A(KEYINPUT54), .B(n958), .ZN(n959) );
  NAND2_X1 U1057 ( .A1(n960), .A2(n959), .ZN(n961) );
  XOR2_X1 U1058 ( .A(KEYINPUT55), .B(KEYINPUT116), .Z(n996) );
  XNOR2_X1 U1059 ( .A(n961), .B(n996), .ZN(n963) );
  INV_X1 U1060 ( .A(G29), .ZN(n962) );
  NAND2_X1 U1061 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1062 ( .A1(G11), .A2(n964), .ZN(n965) );
  XNOR2_X1 U1063 ( .A(KEYINPUT120), .B(n965), .ZN(n966) );
  NOR2_X1 U1064 ( .A1(n967), .A2(n966), .ZN(n1000) );
  XNOR2_X1 U1065 ( .A(G164), .B(G2078), .ZN(n971) );
  XNOR2_X1 U1066 ( .A(G2072), .B(KEYINPUT115), .ZN(n969) );
  XNOR2_X1 U1067 ( .A(n969), .B(n968), .ZN(n970) );
  NAND2_X1 U1068 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1069 ( .A(n972), .B(KEYINPUT50), .ZN(n994) );
  XNOR2_X1 U1070 ( .A(G2084), .B(G160), .ZN(n973) );
  XNOR2_X1 U1071 ( .A(n973), .B(KEYINPUT110), .ZN(n978) );
  NOR2_X1 U1072 ( .A1(n975), .A2(n974), .ZN(n976) );
  XOR2_X1 U1073 ( .A(KEYINPUT111), .B(n976), .Z(n977) );
  NAND2_X1 U1074 ( .A1(n978), .A2(n977), .ZN(n979) );
  NOR2_X1 U1075 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1076 ( .A(KEYINPUT112), .B(n981), .ZN(n983) );
  NAND2_X1 U1077 ( .A1(n983), .A2(n982), .ZN(n989) );
  XNOR2_X1 U1078 ( .A(G2090), .B(G162), .ZN(n984) );
  XNOR2_X1 U1079 ( .A(n984), .B(KEYINPUT113), .ZN(n986) );
  NOR2_X1 U1080 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1081 ( .A(KEYINPUT51), .B(n987), .ZN(n988) );
  NOR2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1083 ( .A(n990), .B(KEYINPUT114), .ZN(n992) );
  NAND2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n993) );
  NOR2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1086 ( .A(KEYINPUT52), .B(n995), .ZN(n997) );
  NAND2_X1 U1087 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1088 ( .A1(n998), .A2(G29), .ZN(n999) );
  NAND2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1029) );
  XOR2_X1 U1090 ( .A(KEYINPUT56), .B(G16), .Z(n1027) );
  XNOR2_X1 U1091 ( .A(G301), .B(G1961), .ZN(n1003) );
  XNOR2_X1 U1092 ( .A(n1001), .B(G1341), .ZN(n1002) );
  NOR2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1017) );
  XOR2_X1 U1094 ( .A(n1004), .B(KEYINPUT121), .Z(n1006) );
  NAND2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1096 ( .A(KEYINPUT122), .B(n1007), .ZN(n1009) );
  XNOR2_X1 U1097 ( .A(G1971), .B(G303), .ZN(n1008) );
  NOR2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1099 ( .A(KEYINPUT123), .B(n1010), .ZN(n1015) );
  XOR2_X1 U1100 ( .A(G168), .B(G1966), .Z(n1011) );
  NOR2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1102 ( .A(KEYINPUT57), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1025) );
  XOR2_X1 U1105 ( .A(G1348), .B(n1018), .Z(n1021) );
  XOR2_X1 U1106 ( .A(n1019), .B(G1956), .Z(n1020) );
  NOR2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1023) );
  NAND2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1109 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NOR2_X1 U1110 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NOR2_X1 U1111 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XNOR2_X1 U1112 ( .A(n1030), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1113 ( .A(G311), .ZN(G150) );
endmodule

