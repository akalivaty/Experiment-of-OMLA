//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 0 0 0 0 1 1 0 0 1 0 0 1 1 0 1 1 1 0 1 1 0 1 0 1 0 1 0 0 0 1 0 0 1 0 1 1 1 1 1 0 1 0 0 1 0 1 0 0 1 0 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:01 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n597, new_n598, new_n599, new_n600, new_n601, new_n602, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n621, new_n622, new_n623, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n632, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n860, new_n861, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G143), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  NAND4_X1  g004(.A1(new_n188), .A2(new_n190), .A3(KEYINPUT0), .A4(G128), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT0), .ZN(new_n192));
  INV_X1    g006(.A(G128), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(new_n193), .A3(KEYINPUT65), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT65), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n195), .B1(KEYINPUT0), .B2(G128), .ZN(new_n196));
  NAND2_X1  g010(.A1(KEYINPUT0), .A2(G128), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n194), .A2(new_n196), .A3(new_n197), .ZN(new_n198));
  XNOR2_X1  g012(.A(G143), .B(G146), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n191), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G104), .ZN(new_n202));
  OAI21_X1  g016(.A(KEYINPUT3), .B1(new_n202), .B2(G107), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT3), .ZN(new_n204));
  INV_X1    g018(.A(G107), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n204), .A2(new_n205), .A3(G104), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n202), .A2(G107), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n203), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT4), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(new_n209), .A3(G101), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT75), .ZN(new_n211));
  INV_X1    g025(.A(G101), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n203), .A2(new_n206), .A3(new_n212), .A4(new_n207), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(KEYINPUT74), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n208), .A2(G101), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n208), .A2(KEYINPUT74), .A3(G101), .ZN(new_n217));
  AND4_X1   g031(.A1(new_n211), .A2(new_n216), .A3(KEYINPUT4), .A4(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n209), .B1(new_n214), .B2(new_n215), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n211), .B1(new_n219), .B2(new_n217), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n201), .B(new_n210), .C1(new_n218), .C2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT11), .ZN(new_n222));
  INV_X1    g036(.A(G134), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n222), .B1(new_n223), .B2(G137), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(G137), .ZN(new_n225));
  INV_X1    g039(.A(G137), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n226), .A2(KEYINPUT11), .A3(G134), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n224), .A2(new_n225), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G131), .ZN(new_n229));
  INV_X1    g043(.A(G131), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n224), .A2(new_n227), .A3(new_n230), .A4(new_n225), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT10), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n193), .A2(KEYINPUT1), .ZN(new_n235));
  AND3_X1   g049(.A1(new_n235), .A2(new_n188), .A3(new_n190), .ZN(new_n236));
  AOI21_X1  g050(.A(G128), .B1(new_n188), .B2(new_n190), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n189), .A2(KEYINPUT1), .A3(G146), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  NOR3_X1   g053(.A1(new_n236), .A2(new_n237), .A3(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n205), .A2(KEYINPUT76), .A3(G104), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT76), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n242), .B1(new_n202), .B2(G107), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n205), .A2(G104), .ZN(new_n244));
  OAI211_X1 g058(.A(G101), .B(new_n241), .C1(new_n243), .C2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(new_n213), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n234), .B1(new_n240), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT77), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n235), .A2(new_n188), .A3(new_n190), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n250), .B(new_n238), .C1(G128), .C2(new_n199), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n251), .A2(new_n213), .A3(new_n245), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n252), .A2(KEYINPUT77), .A3(new_n234), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n246), .A2(KEYINPUT78), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT78), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n255), .B1(new_n245), .B2(new_n213), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n240), .A2(new_n234), .ZN(new_n258));
  AOI22_X1  g072(.A1(new_n249), .A2(new_n253), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n221), .A2(new_n233), .A3(new_n259), .ZN(new_n260));
  XNOR2_X1  g074(.A(G110), .B(G140), .ZN(new_n261));
  INV_X1    g075(.A(G953), .ZN(new_n262));
  AND2_X1   g076(.A1(new_n262), .A2(G227), .ZN(new_n263));
  XOR2_X1   g077(.A(new_n261), .B(new_n263), .Z(new_n264));
  NAND2_X1  g078(.A1(new_n240), .A2(new_n246), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(new_n252), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n233), .B1(new_n266), .B2(KEYINPUT80), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT80), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n265), .A2(new_n268), .A3(new_n252), .ZN(new_n269));
  AOI21_X1  g083(.A(KEYINPUT12), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n266), .A2(KEYINPUT12), .A3(new_n232), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(KEYINPUT79), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT79), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n266), .A2(new_n273), .A3(KEYINPUT12), .A4(new_n232), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n260), .B(new_n264), .C1(new_n270), .C2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT81), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n264), .ZN(new_n279));
  INV_X1    g093(.A(new_n260), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n233), .B1(new_n221), .B2(new_n259), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n266), .A2(KEYINPUT80), .ZN(new_n283));
  AND3_X1   g097(.A1(new_n283), .A2(new_n232), .A3(new_n269), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n272), .B(new_n274), .C1(new_n284), .C2(KEYINPUT12), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n285), .A2(KEYINPUT81), .A3(new_n260), .A4(new_n264), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n278), .A2(new_n282), .A3(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(G469), .ZN(new_n288));
  INV_X1    g102(.A(G902), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(G469), .A2(G902), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n264), .B1(new_n280), .B2(new_n281), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n285), .A2(new_n260), .A3(new_n279), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(G469), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n290), .A2(new_n291), .A3(new_n295), .ZN(new_n296));
  XOR2_X1   g110(.A(KEYINPUT9), .B(G234), .Z(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(G221), .B1(new_n298), .B2(G902), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT82), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n296), .A2(KEYINPUT82), .A3(new_n299), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n200), .A2(KEYINPUT66), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT66), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n306), .B(new_n191), .C1(new_n198), .C2(new_n199), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n305), .A2(new_n232), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(KEYINPUT67), .ZN(new_n309));
  INV_X1    g123(.A(new_n225), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n223), .A2(G137), .ZN(new_n311));
  OAI21_X1  g125(.A(G131), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n251), .A2(new_n231), .A3(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT67), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n305), .A2(new_n314), .A3(new_n232), .A4(new_n307), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n309), .A2(new_n313), .A3(new_n315), .ZN(new_n316));
  XNOR2_X1  g130(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NOR2_X1   g132(.A1(KEYINPUT2), .A2(G113), .ZN(new_n319));
  AND2_X1   g133(.A1(KEYINPUT2), .A2(G113), .ZN(new_n320));
  OR2_X1    g134(.A1(new_n320), .A2(KEYINPUT68), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(KEYINPUT68), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n319), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G119), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G116), .ZN(new_n325));
  INV_X1    g139(.A(G116), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G119), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n323), .B(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n201), .A2(new_n232), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(KEYINPUT30), .A3(new_n313), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n318), .A2(new_n330), .A3(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT31), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n323), .B(new_n328), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n335), .A2(new_n331), .A3(new_n313), .ZN(new_n336));
  XNOR2_X1  g150(.A(KEYINPUT26), .B(G101), .ZN(new_n337));
  NOR2_X1   g151(.A1(G237), .A2(G953), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G210), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n337), .B(new_n339), .ZN(new_n340));
  XNOR2_X1  g154(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n340), .B(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n333), .A2(new_n334), .A3(new_n336), .A4(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT70), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n333), .A2(new_n336), .A3(new_n343), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(KEYINPUT31), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n347), .A2(new_n345), .A3(KEYINPUT31), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n316), .A2(new_n330), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n336), .A2(KEYINPUT28), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT28), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n335), .A2(new_n353), .A3(new_n331), .A4(new_n313), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n343), .B1(new_n351), .B2(new_n355), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n356), .B(KEYINPUT71), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n349), .A2(new_n350), .A3(new_n357), .ZN(new_n358));
  NOR2_X1   g172(.A1(G472), .A2(G902), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT32), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n358), .A2(KEYINPUT32), .A3(new_n359), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n331), .A2(new_n313), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n330), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n355), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n343), .A2(KEYINPUT29), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT29), .ZN(new_n368));
  AND2_X1   g182(.A1(new_n333), .A2(new_n336), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n368), .B1(new_n369), .B2(new_n343), .ZN(new_n370));
  AND3_X1   g184(.A1(new_n351), .A2(new_n343), .A3(new_n355), .ZN(new_n371));
  OAI221_X1 g185(.A(new_n289), .B1(new_n366), .B2(new_n367), .C1(new_n370), .C2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(G472), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n362), .A2(new_n363), .A3(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT73), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT25), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(KEYINPUT73), .A2(KEYINPUT25), .ZN(new_n378));
  XNOR2_X1  g192(.A(G125), .B(G140), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(KEYINPUT16), .ZN(new_n380));
  INV_X1    g194(.A(G140), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G125), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n380), .B1(KEYINPUT16), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n187), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n380), .B(G146), .C1(KEYINPUT16), .C2(new_n382), .ZN(new_n385));
  XNOR2_X1  g199(.A(G119), .B(G128), .ZN(new_n386));
  XOR2_X1   g200(.A(KEYINPUT24), .B(G110), .Z(new_n387));
  AOI22_X1  g201(.A1(new_n384), .A2(new_n385), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n324), .A2(G128), .ZN(new_n389));
  OR2_X1    g203(.A1(new_n389), .A2(KEYINPUT23), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(KEYINPUT23), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n390), .B(new_n391), .C1(G119), .C2(new_n193), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G110), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n388), .A2(new_n393), .ZN(new_n394));
  OAI22_X1  g208(.A1(new_n392), .A2(G110), .B1(new_n386), .B2(new_n387), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n379), .A2(new_n187), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n395), .A2(new_n385), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n262), .A2(G221), .A3(G234), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n399), .B(KEYINPUT22), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n400), .B(G137), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n398), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n394), .A2(new_n397), .A3(new_n401), .ZN(new_n404));
  AND2_X1   g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n377), .B(new_n378), .C1(new_n406), .C2(G902), .ZN(new_n407));
  INV_X1    g221(.A(G234), .ZN(new_n408));
  OAI21_X1  g222(.A(G217), .B1(new_n408), .B2(G902), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n409), .B(KEYINPUT72), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n405), .A2(new_n375), .A3(new_n376), .A4(new_n289), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n407), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(G902), .B1(new_n408), .B2(G217), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n405), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n297), .A2(G217), .A3(new_n262), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT87), .ZN(new_n419));
  AOI21_X1  g233(.A(KEYINPUT13), .B1(new_n189), .B2(G128), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n189), .A2(G128), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n419), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n189), .A2(KEYINPUT13), .A3(G128), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT13), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n424), .B1(new_n193), .B2(G143), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n193), .A2(G143), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n425), .A2(KEYINPUT87), .A3(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n422), .A2(new_n423), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(G134), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT88), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  XNOR2_X1  g245(.A(G116), .B(G122), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n432), .B(new_n205), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n428), .A2(KEYINPUT88), .A3(G134), .ZN(new_n434));
  XNOR2_X1  g248(.A(G128), .B(G143), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(new_n223), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n431), .A2(new_n433), .A3(new_n434), .A4(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(KEYINPUT89), .ZN(new_n438));
  INV_X1    g252(.A(new_n436), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n439), .B1(new_n429), .B2(new_n430), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT89), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n440), .A2(new_n441), .A3(new_n433), .A4(new_n434), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n438), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n432), .A2(new_n205), .ZN(new_n444));
  OAI21_X1  g258(.A(KEYINPUT14), .B1(new_n326), .B2(G122), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n432), .B1(KEYINPUT14), .B2(new_n205), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n435), .B(G134), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n418), .B1(new_n443), .B2(new_n451), .ZN(new_n452));
  AOI211_X1 g266(.A(new_n450), .B(new_n417), .C1(new_n438), .C2(new_n442), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n289), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT15), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n454), .A2(new_n455), .A3(G478), .ZN(new_n456));
  INV_X1    g270(.A(G475), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n338), .A2(G214), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n189), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n338), .A2(G143), .A3(G214), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(G131), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT17), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n459), .A2(new_n230), .A3(new_n460), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n461), .A2(KEYINPUT17), .A3(G131), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n465), .A2(new_n384), .A3(new_n466), .A4(new_n385), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n379), .B(new_n187), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT18), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n469), .A2(new_n230), .ZN(new_n470));
  OAI221_X1 g284(.A(new_n468), .B1(new_n461), .B2(new_n470), .C1(new_n462), .C2(new_n469), .ZN(new_n471));
  XNOR2_X1  g285(.A(G113), .B(G122), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n472), .B(new_n202), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n467), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n462), .A2(new_n464), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n379), .B(KEYINPUT19), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(new_n187), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n476), .A2(new_n478), .A3(new_n385), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n473), .B1(new_n479), .B2(new_n471), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n457), .B(new_n289), .C1(new_n475), .C2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(KEYINPUT20), .ZN(new_n482));
  INV_X1    g296(.A(new_n480), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(new_n474), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT20), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n484), .A2(new_n485), .A3(new_n457), .A4(new_n289), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n473), .B1(new_n467), .B2(new_n471), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n289), .B1(new_n475), .B2(new_n487), .ZN(new_n488));
  XNOR2_X1  g302(.A(KEYINPUT86), .B(G475), .ZN(new_n489));
  AOI22_X1  g303(.A1(new_n482), .A2(new_n486), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  AND2_X1   g304(.A1(new_n262), .A2(G952), .ZN(new_n491));
  NAND2_X1  g305(.A1(G234), .A2(G237), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  XOR2_X1   g307(.A(KEYINPUT21), .B(G898), .Z(new_n494));
  NAND3_X1  g308(.A1(new_n492), .A2(G902), .A3(G953), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n455), .A2(G478), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n289), .B(new_n497), .C1(new_n452), .C2(new_n453), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n456), .A2(new_n490), .A3(new_n496), .A4(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT90), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n499), .B(new_n500), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n330), .B(new_n210), .C1(new_n218), .C2(new_n220), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n323), .A2(new_n329), .ZN(new_n503));
  OAI21_X1  g317(.A(G113), .B1(new_n325), .B2(KEYINPUT5), .ZN(new_n504));
  AND2_X1   g318(.A1(new_n329), .A2(KEYINPUT5), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n257), .B(new_n503), .C1(new_n504), .C2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  XOR2_X1   g321(.A(G110), .B(G122), .Z(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n508), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n502), .A2(new_n510), .A3(new_n506), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n509), .A2(KEYINPUT6), .A3(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT6), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n507), .A2(new_n513), .A3(new_n508), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n200), .A2(G125), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n515), .B1(G125), .B2(new_n251), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n262), .A2(G224), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n517), .B(KEYINPUT83), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n516), .B(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n512), .A2(new_n514), .A3(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n503), .B1(new_n505), .B2(new_n504), .ZN(new_n521));
  INV_X1    g335(.A(new_n246), .ZN(new_n522));
  OAI22_X1  g336(.A1(new_n521), .A2(new_n522), .B1(KEYINPUT8), .B2(new_n508), .ZN(new_n523));
  OR2_X1    g337(.A1(new_n505), .A2(KEYINPUT84), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n505), .A2(KEYINPUT84), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n503), .B1(new_n526), .B2(new_n504), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n523), .B1(new_n527), .B2(new_n522), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n508), .A2(KEYINPUT8), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n517), .A2(KEYINPUT7), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n251), .A2(G125), .ZN(new_n531));
  OR2_X1    g345(.A1(new_n531), .A2(KEYINPUT85), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(KEYINPUT85), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n532), .A2(new_n515), .A3(new_n533), .ZN(new_n534));
  AOI22_X1  g348(.A1(new_n528), .A2(new_n529), .B1(new_n530), .B2(new_n534), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n535), .B(new_n511), .C1(new_n530), .C2(new_n516), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n520), .A2(new_n536), .A3(new_n289), .ZN(new_n537));
  OAI21_X1  g351(.A(G210), .B1(G237), .B2(G902), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n520), .A2(new_n536), .A3(new_n289), .A4(new_n538), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(G214), .B1(G237), .B2(G902), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n501), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n304), .A2(new_n374), .A3(new_n416), .A4(new_n545), .ZN(new_n546));
  XNOR2_X1  g360(.A(KEYINPUT91), .B(G101), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n546), .B(new_n547), .ZN(G3));
  INV_X1    g362(.A(new_n543), .ZN(new_n549));
  AND4_X1   g363(.A1(new_n289), .A2(new_n520), .A3(new_n536), .A4(new_n538), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT93), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n452), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n443), .A2(new_n451), .A3(new_n418), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n553), .A2(KEYINPUT33), .A3(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT33), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n556), .B1(new_n452), .B2(new_n453), .ZN(new_n557));
  INV_X1    g371(.A(G478), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n558), .A2(G902), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n555), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n454), .A2(new_n558), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n490), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n540), .A2(KEYINPUT93), .A3(new_n541), .ZN(new_n566));
  AND4_X1   g380(.A1(new_n496), .A2(new_n552), .A3(new_n565), .A4(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(G472), .ZN(new_n568));
  OR2_X1    g382(.A1(new_n568), .A2(KEYINPUT92), .ZN(new_n569));
  AND3_X1   g383(.A1(new_n358), .A2(new_n289), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n569), .B1(new_n358), .B2(new_n289), .ZN(new_n571));
  NOR3_X1   g385(.A1(new_n570), .A2(new_n571), .A3(new_n415), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n304), .A2(new_n567), .A3(new_n572), .ZN(new_n573));
  XOR2_X1   g387(.A(KEYINPUT34), .B(G104), .Z(new_n574));
  XNOR2_X1  g388(.A(new_n573), .B(new_n574), .ZN(G6));
  NOR2_X1   g389(.A1(new_n558), .A2(KEYINPUT15), .ZN(new_n576));
  AND2_X1   g390(.A1(new_n454), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n498), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n490), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  AND4_X1   g394(.A1(new_n496), .A2(new_n552), .A3(new_n566), .A4(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n304), .A2(new_n572), .A3(new_n581), .ZN(new_n582));
  XOR2_X1   g396(.A(KEYINPUT35), .B(G107), .Z(new_n583));
  XNOR2_X1  g397(.A(new_n582), .B(new_n583), .ZN(G9));
  NOR2_X1   g398(.A1(new_n402), .A2(KEYINPUT36), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n398), .B(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n413), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT94), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n587), .B(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n412), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NOR3_X1   g405(.A1(new_n570), .A2(new_n571), .A3(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n304), .A2(new_n545), .A3(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(KEYINPUT95), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(KEYINPUT37), .ZN(new_n595));
  XOR2_X1   g409(.A(new_n595), .B(G110), .Z(G12));
  OR2_X1    g410(.A1(new_n495), .A2(G900), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n493), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n579), .A2(new_n599), .ZN(new_n600));
  AND4_X1   g414(.A1(new_n566), .A2(new_n552), .A3(new_n600), .A4(new_n590), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n304), .A2(new_n374), .A3(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(G128), .ZN(G30));
  XOR2_X1   g417(.A(new_n598), .B(KEYINPUT39), .Z(new_n604));
  AOI21_X1  g418(.A(new_n604), .B1(new_n302), .B2(new_n303), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT40), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OR2_X1    g421(.A1(new_n605), .A2(new_n606), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n542), .B(KEYINPUT38), .ZN(new_n609));
  AND2_X1   g423(.A1(new_n365), .A2(new_n336), .ZN(new_n610));
  OAI211_X1 g424(.A(new_n347), .B(G472), .C1(new_n343), .C2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(G472), .A2(G902), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(KEYINPUT96), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n362), .A2(new_n363), .A3(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n577), .A2(new_n578), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n616), .A2(new_n490), .ZN(new_n617));
  AND4_X1   g431(.A1(new_n543), .A2(new_n615), .A3(new_n591), .A4(new_n617), .ZN(new_n618));
  AND4_X1   g432(.A1(new_n607), .A2(new_n608), .A3(new_n609), .A4(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(new_n189), .ZN(G45));
  AND3_X1   g434(.A1(new_n552), .A2(new_n566), .A3(new_n590), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n564), .A2(new_n599), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n304), .A2(new_n374), .A3(new_n621), .A4(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(G146), .ZN(G48));
  AND3_X1   g438(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n288), .B1(new_n287), .B2(new_n289), .ZN(new_n626));
  INV_X1    g440(.A(new_n299), .ZN(new_n627));
  NOR3_X1   g441(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n567), .A2(new_n374), .A3(new_n416), .A4(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(KEYINPUT41), .B(G113), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G15));
  NAND4_X1  g445(.A1(new_n581), .A2(new_n374), .A3(new_n416), .A4(new_n628), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(G116), .ZN(G18));
  XNOR2_X1  g447(.A(new_n499), .B(KEYINPUT90), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n621), .A2(new_n374), .A3(new_n634), .A4(new_n628), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G119), .ZN(G21));
  AND3_X1   g450(.A1(new_n552), .A2(new_n566), .A3(new_n617), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n568), .B1(new_n358), .B2(new_n289), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n366), .B(KEYINPUT97), .ZN(new_n639));
  OAI211_X1 g453(.A(new_n348), .B(new_n344), .C1(new_n639), .C2(new_n343), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n359), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n638), .A2(new_n642), .A3(new_n415), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n637), .A2(new_n643), .A3(new_n496), .A4(new_n628), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(G122), .ZN(G24));
  NOR2_X1   g459(.A1(new_n638), .A2(new_n642), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n621), .A2(new_n646), .A3(new_n622), .A4(new_n628), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G125), .ZN(G27));
  XNOR2_X1  g462(.A(new_n291), .B(KEYINPUT98), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n290), .A2(new_n295), .A3(new_n650), .ZN(new_n651));
  AND2_X1   g465(.A1(new_n651), .A2(new_n299), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n542), .A2(new_n549), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n374), .A2(new_n416), .A3(new_n652), .A4(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n622), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT42), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(KEYINPUT99), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  OR3_X1    g472(.A1(new_n654), .A2(new_n655), .A3(new_n658), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n658), .B1(new_n654), .B2(new_n655), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G131), .ZN(G33));
  AND2_X1   g476(.A1(new_n600), .A2(KEYINPUT100), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n600), .A2(KEYINPUT100), .ZN(new_n664));
  NOR3_X1   g478(.A1(new_n654), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(new_n223), .ZN(G36));
  XOR2_X1   g480(.A(new_n294), .B(KEYINPUT45), .Z(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(G469), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT101), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n667), .A2(KEYINPUT101), .A3(G469), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n649), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT46), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n625), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n672), .A2(KEYINPUT46), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n627), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n604), .ZN(new_n678));
  INV_X1    g492(.A(new_n653), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n562), .A2(new_n490), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(KEYINPUT43), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n570), .A2(new_n571), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n681), .A2(new_n682), .A3(new_n591), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n679), .B1(new_n683), .B2(KEYINPUT44), .ZN(new_n684));
  OR2_X1    g498(.A1(new_n683), .A2(KEYINPUT44), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n677), .A2(new_n678), .A3(new_n684), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G137), .ZN(G39));
  NAND2_X1  g501(.A1(new_n675), .A2(new_n676), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(new_n299), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(KEYINPUT47), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n374), .A2(new_n416), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT47), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n677), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n679), .A2(new_n655), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n690), .A2(new_n691), .A3(new_n693), .A4(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT102), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G140), .ZN(G42));
  INV_X1    g511(.A(new_n681), .ZN(new_n698));
  AND4_X1   g512(.A1(new_n492), .A2(new_n698), .A3(new_n491), .A4(new_n643), .ZN(new_n699));
  INV_X1    g513(.A(new_n628), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n700), .A2(new_n543), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n699), .B1(KEYINPUT111), .B2(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(KEYINPUT112), .A2(KEYINPUT50), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n609), .B1(new_n701), .B2(KEYINPUT111), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  OR3_X1    g519(.A1(new_n702), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n703), .B1(new_n702), .B2(new_n705), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n679), .A2(new_n700), .A3(new_n493), .ZN(new_n709));
  INV_X1    g523(.A(new_n615), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n709), .A2(new_n416), .A3(new_n710), .ZN(new_n711));
  XOR2_X1   g525(.A(new_n711), .B(KEYINPUT115), .Z(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n490), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n708), .B1(new_n713), .B2(new_n562), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n690), .A2(new_n693), .ZN(new_n715));
  NOR3_X1   g529(.A1(new_n625), .A2(new_n626), .A3(new_n299), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n679), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n714), .B1(new_n718), .B2(new_n699), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n709), .A2(new_n698), .ZN(new_n720));
  XOR2_X1   g534(.A(new_n720), .B(KEYINPUT113), .Z(new_n721));
  NAND3_X1  g535(.A1(new_n721), .A2(new_n590), .A3(new_n646), .ZN(new_n722));
  XOR2_X1   g536(.A(new_n722), .B(KEYINPUT114), .Z(new_n723));
  AND3_X1   g537(.A1(new_n719), .A2(KEYINPUT51), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g538(.A(KEYINPUT51), .B1(new_n719), .B2(new_n723), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT53), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n632), .A2(new_n635), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n358), .A2(new_n289), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(G472), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n628), .A2(new_n730), .A3(new_n416), .A4(new_n641), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n552), .A2(new_n566), .A3(new_n496), .A4(new_n617), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n374), .A2(new_n416), .A3(new_n628), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n733), .B1(new_n734), .B2(new_n567), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT104), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n728), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n629), .A2(new_n632), .A3(new_n635), .A4(new_n644), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(KEYINPUT104), .ZN(new_n739));
  AND2_X1   g553(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n616), .A2(new_n490), .A3(new_n598), .ZN(new_n741));
  XOR2_X1   g555(.A(new_n741), .B(KEYINPUT106), .Z(new_n742));
  NAND3_X1  g556(.A1(new_n742), .A2(new_n304), .A3(new_n374), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n646), .A2(new_n652), .A3(new_n622), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n679), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(new_n590), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n665), .B1(new_n659), .B2(new_n660), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n564), .A2(new_n579), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n549), .B1(new_n540), .B2(new_n541), .ZN(new_n749));
  AND3_X1   g563(.A1(new_n748), .A2(new_n749), .A3(new_n496), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n304), .A2(new_n572), .A3(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n546), .A2(new_n593), .A3(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT105), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n546), .A2(new_n593), .A3(new_n751), .A4(KEYINPUT105), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n740), .A2(new_n746), .A3(new_n747), .A4(new_n756), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n628), .A2(new_n566), .A3(new_n552), .A4(new_n590), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n730), .A2(new_n622), .A3(new_n641), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n363), .ZN(new_n761));
  AOI21_X1  g575(.A(KEYINPUT32), .B1(new_n358), .B2(new_n359), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  AOI22_X1  g577(.A1(new_n763), .A2(new_n373), .B1(new_n302), .B2(new_n303), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n760), .B1(new_n764), .B2(new_n601), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT108), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT107), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n767), .B1(new_n590), .B2(new_n599), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n412), .A2(new_n589), .A3(KEYINPUT107), .A4(new_n598), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n637), .A2(new_n615), .A3(new_n770), .A4(new_n652), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n765), .A2(new_n766), .A3(new_n623), .A4(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n623), .A2(new_n602), .A3(new_n647), .A4(new_n771), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(KEYINPUT108), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(KEYINPUT52), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT52), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n772), .A2(new_n774), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n727), .B1(new_n757), .B2(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n727), .B1(new_n745), .B2(new_n590), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n756), .A2(new_n747), .A3(new_n781), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n782), .A2(new_n738), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT109), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n773), .A2(KEYINPUT52), .ZN(new_n785));
  AND3_X1   g599(.A1(new_n778), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n784), .B1(new_n778), .B2(new_n785), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n783), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT54), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n780), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n415), .B1(new_n763), .B2(new_n373), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n304), .B(new_n545), .C1(new_n791), .C2(new_n592), .ZN(new_n792));
  AOI21_X1  g606(.A(KEYINPUT105), .B1(new_n792), .B2(new_n751), .ZN(new_n793));
  AND4_X1   g607(.A1(KEYINPUT105), .A2(new_n546), .A3(new_n593), .A4(new_n751), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n737), .B(new_n739), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n746), .ZN(new_n796));
  INV_X1    g610(.A(new_n747), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n798), .B1(new_n786), .B2(new_n787), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(new_n727), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n772), .A2(new_n774), .A3(new_n777), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n777), .B1(new_n772), .B2(new_n774), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AND4_X1   g617(.A1(new_n747), .A2(new_n756), .A3(new_n737), .A4(new_n739), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n803), .A2(new_n804), .A3(KEYINPUT53), .A4(new_n746), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT110), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n798), .A2(new_n803), .A3(KEYINPUT110), .A4(KEYINPUT53), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n800), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n790), .B1(new_n809), .B2(KEYINPUT54), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT116), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n712), .A2(new_n565), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n721), .A2(new_n791), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n813), .A2(KEYINPUT48), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n813), .A2(KEYINPUT48), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n491), .B(new_n812), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n699), .A2(new_n566), .A3(new_n552), .A4(new_n628), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n811), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  OR3_X1    g633(.A1(new_n816), .A2(new_n811), .A3(new_n818), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n726), .A2(new_n810), .A3(new_n819), .A4(new_n820), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n821), .B1(G952), .B2(G953), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n415), .A2(new_n627), .A3(new_n549), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n823), .A2(KEYINPUT103), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n609), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n680), .B1(new_n823), .B2(KEYINPUT103), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n625), .A2(new_n626), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(KEYINPUT49), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n825), .A2(new_n710), .A3(new_n826), .A4(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n822), .A2(new_n829), .ZN(G75));
  NAND2_X1  g644(.A1(new_n512), .A2(new_n514), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(KEYINPUT117), .ZN(new_n832));
  XOR2_X1   g646(.A(new_n832), .B(KEYINPUT118), .Z(new_n833));
  XOR2_X1   g647(.A(new_n519), .B(KEYINPUT55), .Z(new_n834));
  AOI21_X1  g648(.A(new_n289), .B1(new_n780), .B2(new_n788), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(G210), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT56), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n834), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(new_n834), .ZN(new_n840));
  AOI211_X1 g654(.A(KEYINPUT56), .B(new_n840), .C1(new_n835), .C2(G210), .ZN(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n833), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n833), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n838), .A2(new_n841), .A3(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n262), .A2(G952), .ZN(new_n846));
  XOR2_X1   g660(.A(new_n846), .B(KEYINPUT119), .Z(new_n847));
  NOR3_X1   g661(.A1(new_n843), .A2(new_n845), .A3(new_n847), .ZN(G51));
  INV_X1    g662(.A(new_n790), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n780), .A2(new_n788), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(KEYINPUT54), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n649), .B(KEYINPUT120), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(KEYINPUT57), .ZN(new_n854));
  OR2_X1    g668(.A1(new_n853), .A2(KEYINPUT57), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n852), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(new_n287), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n835), .A2(new_n670), .A3(new_n671), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n846), .B1(new_n857), .B2(new_n858), .ZN(G54));
  NAND3_X1  g673(.A1(new_n835), .A2(KEYINPUT58), .A3(G475), .ZN(new_n860));
  XOR2_X1   g674(.A(new_n860), .B(new_n484), .Z(new_n861));
  NOR2_X1   g675(.A1(new_n861), .A2(new_n846), .ZN(G60));
  AND2_X1   g676(.A1(new_n555), .A2(new_n557), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  XNOR2_X1  g678(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n865));
  NAND2_X1  g679(.A1(G478), .A2(G902), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n865), .B(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n864), .B1(new_n810), .B2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT122), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n867), .B1(new_n849), .B2(new_n851), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n847), .B1(new_n871), .B2(new_n863), .ZN(new_n872));
  OAI211_X1 g686(.A(KEYINPUT122), .B(new_n864), .C1(new_n810), .C2(new_n867), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n870), .A2(new_n872), .A3(new_n873), .ZN(G63));
  NAND2_X1  g688(.A1(G217), .A2(G902), .ZN(new_n875));
  XOR2_X1   g689(.A(new_n875), .B(KEYINPUT60), .Z(new_n876));
  NAND2_X1  g690(.A1(new_n850), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n847), .B1(new_n877), .B2(new_n406), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n850), .A2(new_n586), .A3(new_n876), .ZN(new_n879));
  AOI22_X1  g693(.A1(new_n878), .A2(new_n879), .B1(KEYINPUT123), .B2(KEYINPUT61), .ZN(new_n880));
  NOR2_X1   g694(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n880), .B(new_n881), .ZN(G66));
  NAND2_X1  g696(.A1(new_n795), .A2(new_n262), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n494), .A2(G224), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n883), .B(KEYINPUT124), .C1(new_n262), .C2(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n885), .B1(KEYINPUT124), .B2(new_n883), .ZN(new_n886));
  INV_X1    g700(.A(G898), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n832), .B1(new_n887), .B2(G953), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n886), .B(new_n888), .ZN(G69));
  AOI21_X1  g703(.A(new_n262), .B1(G227), .B2(G900), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  OR2_X1    g705(.A1(new_n262), .A2(G900), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n318), .A2(new_n332), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n477), .B(KEYINPUT125), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n893), .B(new_n894), .Z(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n695), .A2(new_n686), .A3(new_n747), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n677), .A2(new_n678), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n791), .A2(new_n637), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n623), .B(new_n765), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  OAI211_X1 g715(.A(new_n892), .B(new_n896), .C1(new_n901), .C2(G953), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n765), .A2(new_n623), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n619), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT62), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n791), .A2(new_n605), .A3(new_n653), .A4(new_n748), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n905), .A2(new_n686), .A3(new_n695), .A4(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n907), .A2(new_n262), .A3(new_n895), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n891), .B1(new_n902), .B2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  XNOR2_X1  g724(.A(KEYINPUT126), .B(KEYINPUT127), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n902), .A2(new_n908), .A3(new_n891), .ZN(new_n912));
  AND3_X1   g726(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n911), .B1(new_n910), .B2(new_n912), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n913), .A2(new_n914), .ZN(G72));
  XOR2_X1   g729(.A(new_n612), .B(KEYINPUT63), .Z(new_n916));
  OR2_X1    g730(.A1(new_n369), .A2(new_n342), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n369), .A2(new_n342), .ZN(new_n918));
  AND4_X1   g732(.A1(new_n809), .A2(new_n916), .A3(new_n917), .A4(new_n918), .ZN(new_n919));
  OR2_X1    g733(.A1(new_n907), .A2(new_n795), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n917), .B1(new_n920), .B2(new_n916), .ZN(new_n921));
  INV_X1    g735(.A(new_n795), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n901), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n918), .B1(new_n923), .B2(new_n916), .ZN(new_n924));
  NOR4_X1   g738(.A1(new_n919), .A2(new_n921), .A3(new_n924), .A4(new_n846), .ZN(G57));
endmodule


