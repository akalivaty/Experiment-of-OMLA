//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 0 0 1 0 0 0 0 1 0 1 1 1 0 1 0 0 0 1 0 0 0 0 1 0 0 1 1 1 1 0 0 0 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:02 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n771,
    new_n772, new_n773, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n794,
    new_n795, new_n796, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT65), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT65), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n188), .A2(new_n190), .A3(G143), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT64), .ZN(new_n192));
  INV_X1    g006(.A(G143), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(KEYINPUT64), .A2(G143), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n194), .A2(G146), .A3(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT1), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n191), .A2(new_n196), .A3(new_n197), .A4(G128), .ZN(new_n198));
  AND2_X1   g012(.A1(new_n191), .A2(new_n196), .ZN(new_n199));
  INV_X1    g013(.A(G128), .ZN(new_n200));
  AND2_X1   g014(.A1(KEYINPUT64), .A2(G143), .ZN(new_n201));
  NOR2_X1   g015(.A1(KEYINPUT64), .A2(G143), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n187), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n200), .B1(new_n203), .B2(KEYINPUT1), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n198), .B1(new_n199), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT3), .ZN(new_n206));
  INV_X1    g020(.A(G104), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n206), .B1(new_n207), .B2(G107), .ZN(new_n208));
  INV_X1    g022(.A(G107), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n209), .A2(KEYINPUT3), .A3(G104), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G101), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT80), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n213), .B1(new_n209), .B2(G104), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n207), .A2(KEYINPUT80), .A3(G107), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n211), .A2(new_n212), .A3(new_n214), .A4(new_n215), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n207), .A2(G107), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n209), .A2(G104), .ZN(new_n218));
  OAI21_X1  g032(.A(G101), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  AND2_X1   g033(.A1(new_n216), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT10), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n205), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n216), .A2(new_n219), .ZN(new_n223));
  XNOR2_X1  g037(.A(KEYINPUT65), .B(G146), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n197), .B1(new_n224), .B2(G143), .ZN(new_n225));
  AOI21_X1  g039(.A(G146), .B1(new_n194), .B2(new_n195), .ZN(new_n226));
  AOI21_X1  g040(.A(G143), .B1(new_n188), .B2(new_n190), .ZN(new_n227));
  OAI22_X1  g041(.A1(new_n225), .A2(new_n200), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n223), .B1(new_n228), .B2(new_n198), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n222), .B1(new_n229), .B2(new_n221), .ZN(new_n230));
  AND3_X1   g044(.A1(new_n209), .A2(KEYINPUT3), .A3(G104), .ZN(new_n231));
  AOI21_X1  g045(.A(KEYINPUT3), .B1(new_n209), .B2(G104), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n214), .B(new_n215), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT81), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n211), .A2(KEYINPUT81), .A3(new_n214), .A4(new_n215), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n235), .A2(G101), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n216), .A2(KEYINPUT4), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  AND2_X1   g054(.A1(KEYINPUT0), .A2(G128), .ZN(new_n241));
  NOR2_X1   g055(.A1(KEYINPUT0), .A2(G128), .ZN(new_n242));
  OR2_X1    g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n189), .A2(G146), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n187), .A2(KEYINPUT65), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n193), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n243), .B1(new_n246), .B2(new_n203), .ZN(new_n247));
  AND3_X1   g061(.A1(new_n191), .A2(new_n196), .A3(new_n241), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XOR2_X1   g063(.A(KEYINPUT82), .B(KEYINPUT4), .Z(new_n250));
  NAND4_X1  g064(.A1(new_n235), .A2(G101), .A3(new_n236), .A4(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n240), .A2(new_n249), .A3(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT11), .ZN(new_n253));
  INV_X1    g067(.A(G134), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n253), .B1(new_n254), .B2(G137), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(G137), .ZN(new_n256));
  INV_X1    g070(.A(G137), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n257), .A2(KEYINPUT11), .A3(G134), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n255), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G131), .ZN(new_n260));
  INV_X1    g074(.A(G131), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n255), .A2(new_n258), .A3(new_n261), .A4(new_n256), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n230), .A2(new_n252), .A3(new_n264), .ZN(new_n265));
  XNOR2_X1  g079(.A(G110), .B(G140), .ZN(new_n266));
  INV_X1    g080(.A(G953), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G227), .ZN(new_n268));
  XOR2_X1   g082(.A(new_n266), .B(new_n268), .Z(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT83), .ZN(new_n271));
  AOI211_X1 g085(.A(new_n271), .B(new_n264), .C1(new_n230), .C2(new_n252), .ZN(new_n272));
  AND3_X1   g086(.A1(new_n205), .A2(new_n220), .A3(new_n221), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n227), .A2(new_n226), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n200), .B1(new_n191), .B2(KEYINPUT1), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n198), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n221), .B1(new_n276), .B2(new_n220), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n251), .A2(new_n249), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n212), .B1(new_n233), .B2(new_n234), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n238), .B1(new_n236), .B2(new_n279), .ZN(new_n280));
  OAI22_X1  g094(.A1(new_n273), .A2(new_n277), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(KEYINPUT83), .B1(new_n281), .B2(new_n263), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n265), .B(new_n270), .C1(new_n272), .C2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n205), .A2(new_n220), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n228), .A2(new_n223), .A3(new_n198), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n264), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT12), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n286), .B(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n265), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n269), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(G902), .B1(new_n283), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G469), .ZN(new_n292));
  OAI21_X1  g106(.A(KEYINPUT84), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(G902), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n265), .A2(new_n270), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n281), .A2(new_n263), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(new_n271), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n281), .A2(KEYINPUT83), .A3(new_n263), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n295), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  XNOR2_X1  g113(.A(new_n286), .B(KEYINPUT12), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n270), .B1(new_n300), .B2(new_n265), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n294), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT84), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n302), .A2(new_n303), .A3(G469), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n297), .A2(new_n298), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n270), .B1(new_n305), .B2(new_n265), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n288), .A2(new_n295), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n292), .B(new_n294), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n293), .A2(new_n304), .A3(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT89), .ZN(new_n310));
  INV_X1    g124(.A(G140), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G125), .ZN(new_n312));
  INV_X1    g126(.A(G125), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G140), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT76), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n312), .A2(new_n314), .A3(new_n315), .A4(KEYINPUT16), .ZN(new_n316));
  AND3_X1   g130(.A1(new_n312), .A2(new_n314), .A3(KEYINPUT16), .ZN(new_n317));
  OAI21_X1  g131(.A(KEYINPUT76), .B1(new_n312), .B2(KEYINPUT16), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G146), .ZN(new_n320));
  XNOR2_X1  g134(.A(G125), .B(G140), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n321), .A2(KEYINPUT19), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n321), .A2(KEYINPUT19), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n224), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G237), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n325), .A2(new_n267), .A3(G214), .ZN(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT64), .B(G143), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n326), .B1(new_n327), .B2(KEYINPUT88), .ZN(new_n328));
  INV_X1    g142(.A(G214), .ZN(new_n329));
  NOR3_X1   g143(.A1(new_n329), .A2(G237), .A3(G953), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT88), .ZN(new_n331));
  OAI211_X1 g145(.A(new_n330), .B(new_n193), .C1(new_n192), .C2(new_n331), .ZN(new_n332));
  AND3_X1   g146(.A1(new_n328), .A2(G131), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(G131), .B1(new_n328), .B2(new_n332), .ZN(new_n334));
  OAI211_X1 g148(.A(new_n320), .B(new_n324), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n328), .A2(new_n332), .ZN(new_n336));
  NAND2_X1  g150(.A1(KEYINPUT18), .A2(G131), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n328), .A2(new_n332), .A3(KEYINPUT18), .A4(G131), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n224), .A2(new_n321), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n312), .A2(new_n314), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G146), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n338), .A2(new_n339), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n335), .A2(new_n344), .ZN(new_n345));
  XNOR2_X1  g159(.A(G113), .B(G122), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n346), .B(new_n207), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  NOR3_X1   g163(.A1(new_n333), .A2(new_n334), .A3(KEYINPUT17), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n187), .B(new_n316), .C1(new_n317), .C2(new_n318), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n328), .A2(new_n332), .A3(KEYINPUT17), .A4(G131), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n320), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n347), .B(new_n344), .C1(new_n350), .C2(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n310), .B1(new_n349), .B2(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n347), .B1(new_n335), .B2(new_n344), .ZN(new_n356));
  AND3_X1   g170(.A1(new_n320), .A2(new_n351), .A3(new_n352), .ZN(new_n357));
  INV_X1    g171(.A(new_n334), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT17), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n328), .A2(new_n332), .A3(G131), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  AOI22_X1  g175(.A1(new_n336), .A2(new_n337), .B1(new_n340), .B2(new_n342), .ZN(new_n362));
  AOI22_X1  g176(.A1(new_n357), .A2(new_n361), .B1(new_n339), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n356), .B1(new_n363), .B2(new_n347), .ZN(new_n364));
  NOR2_X1   g178(.A1(G475), .A2(G902), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  OAI22_X1  g180(.A1(new_n355), .A2(KEYINPUT20), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n349), .A2(new_n354), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT20), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n368), .A2(new_n310), .A3(new_n369), .A4(new_n365), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  XNOR2_X1  g185(.A(G116), .B(G122), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n372), .B(new_n209), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n194), .A2(G128), .A3(new_n195), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n200), .A2(G143), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n374), .A2(new_n254), .A3(new_n375), .ZN(new_n376));
  AND3_X1   g190(.A1(new_n374), .A2(KEYINPUT13), .A3(new_n375), .ZN(new_n377));
  OAI21_X1  g191(.A(G134), .B1(new_n374), .B2(KEYINPUT13), .ZN(new_n378));
  OAI211_X1 g192(.A(new_n373), .B(new_n376), .C1(new_n377), .C2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G122), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G116), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n209), .B1(new_n381), .B2(KEYINPUT14), .ZN(new_n382));
  INV_X1    g196(.A(G116), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G122), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  OR2_X1    g199(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n382), .A2(new_n385), .ZN(new_n387));
  INV_X1    g201(.A(new_n376), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n254), .B1(new_n374), .B2(new_n375), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n386), .B(new_n387), .C1(new_n388), .C2(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(KEYINPUT9), .B(G234), .ZN(new_n391));
  INV_X1    g205(.A(G217), .ZN(new_n392));
  NOR3_X1   g206(.A1(new_n391), .A2(new_n392), .A3(G953), .ZN(new_n393));
  AND3_X1   g207(.A1(new_n379), .A2(new_n390), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n393), .B1(new_n379), .B2(new_n390), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n294), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT15), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n396), .A2(new_n397), .A3(G478), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(G478), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n294), .B(new_n399), .C1(new_n394), .C2(new_n395), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  NOR2_X1   g215(.A1(KEYINPUT90), .A2(G952), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(KEYINPUT90), .A2(G952), .ZN(new_n404));
  AOI21_X1  g218(.A(G953), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(G234), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n405), .B1(new_n406), .B2(new_n325), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(KEYINPUT21), .B(G898), .ZN(new_n409));
  AOI211_X1 g223(.A(new_n294), .B(new_n267), .C1(G234), .C2(G237), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n408), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n401), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(G475), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n344), .B1(new_n350), .B2(new_n353), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n348), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(new_n354), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n413), .B1(new_n416), .B2(new_n294), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n371), .A2(new_n412), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(KEYINPUT91), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n417), .B1(new_n367), .B2(new_n370), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT91), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n421), .A2(new_n422), .A3(new_n412), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(G221), .B1(new_n391), .B2(G902), .ZN(new_n425));
  XOR2_X1   g239(.A(new_n425), .B(KEYINPUT79), .Z(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(G214), .B1(G237), .B2(G902), .ZN(new_n428));
  XOR2_X1   g242(.A(new_n428), .B(KEYINPUT85), .Z(new_n429));
  INV_X1    g243(.A(G119), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(G116), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n383), .A2(G119), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n431), .A2(new_n432), .A3(KEYINPUT5), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT5), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n434), .A2(new_n430), .A3(G116), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n433), .A2(G113), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(KEYINPUT2), .A2(G113), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(KEYINPUT67), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT67), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n439), .A2(KEYINPUT2), .A3(G113), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  OR2_X1    g255(.A1(KEYINPUT2), .A2(G113), .ZN(new_n442));
  XNOR2_X1  g256(.A(G116), .B(G119), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n436), .A2(new_n444), .ZN(new_n445));
  OR2_X1    g259(.A1(new_n223), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n441), .A2(new_n442), .ZN(new_n447));
  INV_X1    g261(.A(new_n443), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n444), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n251), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n446), .B1(new_n451), .B2(new_n280), .ZN(new_n452));
  XNOR2_X1  g266(.A(G110), .B(G122), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n453), .B(new_n446), .C1(new_n451), .C2(new_n280), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n455), .A2(KEYINPUT6), .A3(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT6), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n452), .A2(new_n458), .A3(new_n454), .ZN(new_n459));
  OAI21_X1  g273(.A(G125), .B1(new_n247), .B2(new_n248), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n313), .B(new_n198), .C1(new_n274), .C2(new_n275), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(G224), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n463), .A2(G953), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n462), .B(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n457), .A2(new_n459), .A3(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT7), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n460), .A2(new_n461), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n468), .B1(new_n460), .B2(new_n461), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n453), .B(KEYINPUT8), .ZN(new_n472));
  NOR3_X1   g286(.A1(new_n383), .A2(KEYINPUT5), .A3(G119), .ZN(new_n473));
  INV_X1    g287(.A(G113), .ZN(new_n474));
  OAI21_X1  g288(.A(KEYINPUT86), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT86), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n435), .A2(new_n476), .A3(G113), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n475), .A2(new_n433), .A3(new_n477), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n478), .A2(new_n444), .A3(new_n216), .A4(new_n219), .ZN(new_n479));
  AOI22_X1  g293(.A1(new_n216), .A2(new_n219), .B1(new_n436), .B2(new_n444), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n479), .B1(new_n480), .B2(KEYINPUT87), .ZN(new_n481));
  AND3_X1   g295(.A1(new_n223), .A2(KEYINPUT87), .A3(new_n445), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n472), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n471), .A2(new_n456), .A3(new_n483), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n484), .A2(new_n294), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n466), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(G210), .B1(G237), .B2(G902), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n466), .A2(new_n485), .A3(new_n487), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n429), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n309), .A2(new_n424), .A3(new_n427), .A4(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT92), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n489), .A2(new_n490), .ZN(new_n495));
  INV_X1    g309(.A(new_n429), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n497), .B1(new_n423), .B2(new_n420), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n498), .A2(KEYINPUT92), .A3(new_n427), .A4(new_n309), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n494), .A2(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(G472), .A2(G902), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT32), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT31), .ZN(new_n505));
  XNOR2_X1  g319(.A(KEYINPUT26), .B(G101), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n325), .A2(new_n267), .A3(G210), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n506), .B(new_n507), .ZN(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n509));
  XOR2_X1   g323(.A(new_n508), .B(new_n509), .Z(new_n510));
  INV_X1    g324(.A(new_n256), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n254), .A2(G137), .ZN(new_n512));
  OAI21_X1  g326(.A(G131), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n262), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n191), .A2(KEYINPUT1), .ZN(new_n516));
  AOI22_X1  g330(.A1(new_n516), .A2(G128), .B1(new_n246), .B2(new_n203), .ZN(new_n517));
  AND4_X1   g331(.A1(new_n197), .A2(new_n191), .A3(new_n196), .A4(G128), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n515), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n241), .A2(new_n242), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n520), .B1(new_n227), .B2(new_n226), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n191), .A2(new_n196), .A3(new_n241), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n263), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n450), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n519), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT70), .ZN(new_n526));
  AND3_X1   g340(.A1(new_n510), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n526), .B1(new_n510), .B2(new_n525), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT66), .ZN(new_n531));
  AOI22_X1  g345(.A1(new_n263), .A2(new_n249), .B1(new_n276), .B2(new_n515), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n531), .B1(new_n532), .B2(KEYINPUT30), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n519), .A2(new_n523), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT30), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n534), .A2(KEYINPUT66), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n524), .B1(new_n532), .B2(KEYINPUT30), .ZN(new_n538));
  AOI21_X1  g352(.A(KEYINPUT68), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(KEYINPUT66), .B1(new_n534), .B2(new_n535), .ZN(new_n540));
  AOI211_X1 g354(.A(new_n531), .B(KEYINPUT30), .C1(new_n519), .C2(new_n523), .ZN(new_n541));
  OAI211_X1 g355(.A(KEYINPUT68), .B(new_n538), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n505), .B(new_n530), .C1(new_n539), .C2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT73), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n450), .B1(new_n534), .B2(KEYINPUT72), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT72), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n519), .A2(new_n547), .A3(new_n523), .ZN(new_n548));
  AOI21_X1  g362(.A(KEYINPUT28), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT28), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n524), .B1(new_n519), .B2(new_n523), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n550), .B1(new_n552), .B2(new_n525), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n508), .B(new_n509), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n555), .B(KEYINPUT71), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n545), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n514), .B1(new_n228), .B2(new_n198), .ZN(new_n558));
  AND3_X1   g372(.A1(new_n263), .A2(new_n521), .A3(new_n522), .ZN(new_n559));
  OAI21_X1  g373(.A(KEYINPUT72), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n560), .A2(new_n524), .A3(new_n548), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(new_n550), .ZN(new_n562));
  INV_X1    g376(.A(new_n525), .ZN(new_n563));
  OAI21_X1  g377(.A(KEYINPUT28), .B1(new_n563), .B2(new_n551), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n556), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n565), .A2(KEYINPUT73), .A3(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n544), .A2(new_n557), .A3(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n538), .B1(new_n540), .B2(new_n541), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT68), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n529), .B1(new_n571), .B2(new_n542), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n572), .A2(new_n505), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n504), .B1(new_n568), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT29), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n575), .B1(new_n565), .B2(new_n566), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n525), .B1(new_n539), .B2(new_n543), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n576), .B1(new_n577), .B2(new_n555), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n510), .A2(KEYINPUT29), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n294), .B1(new_n565), .B2(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(G472), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n574), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n530), .B1(new_n539), .B2(new_n543), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(KEYINPUT31), .ZN(new_n584));
  AOI21_X1  g398(.A(KEYINPUT73), .B1(new_n565), .B2(new_n566), .ZN(new_n585));
  AOI211_X1 g399(.A(new_n545), .B(new_n556), .C1(new_n562), .C2(new_n564), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n584), .A2(new_n587), .A3(new_n544), .ZN(new_n588));
  AOI21_X1  g402(.A(KEYINPUT32), .B1(new_n588), .B2(new_n501), .ZN(new_n589));
  OAI21_X1  g403(.A(KEYINPUT74), .B1(new_n582), .B2(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n501), .B1(new_n568), .B2(new_n573), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n503), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT74), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n592), .A2(new_n593), .A3(new_n574), .A4(new_n581), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n392), .B1(G234), .B2(new_n294), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NOR2_X1   g410(.A1(KEYINPUT78), .A2(KEYINPUT25), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n320), .A2(new_n351), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n200), .A2(KEYINPUT23), .A3(G119), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n430), .A2(G128), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n430), .A2(G128), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n599), .B(new_n600), .C1(new_n601), .C2(KEYINPUT23), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(G110), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT75), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n602), .A2(KEYINPUT75), .A3(G110), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  XOR2_X1   g421(.A(KEYINPUT24), .B(G110), .Z(new_n608));
  XNOR2_X1  g422(.A(G119), .B(G128), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n598), .A2(new_n607), .A3(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT77), .B(G110), .Z(new_n612));
  OAI22_X1  g426(.A1(new_n602), .A2(new_n612), .B1(new_n608), .B2(new_n609), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n320), .A2(new_n613), .A3(new_n340), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(KEYINPUT22), .B(G137), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n267), .A2(G221), .A3(G234), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n611), .A2(new_n614), .A3(new_n618), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n597), .B1(new_n622), .B2(G902), .ZN(new_n623));
  AND3_X1   g437(.A1(new_n611), .A2(new_n614), .A3(new_n618), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n618), .B1(new_n611), .B2(new_n614), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n597), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n626), .A2(new_n294), .A3(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n596), .B1(new_n623), .B2(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n595), .A2(G902), .ZN(new_n630));
  AND2_X1   g444(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n590), .A2(new_n594), .A3(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n500), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(new_n212), .ZN(G3));
  INV_X1    g449(.A(G472), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n636), .B1(new_n588), .B2(new_n294), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n544), .A2(new_n557), .A3(new_n567), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n502), .B1(new_n638), .B2(new_n584), .ZN(new_n639));
  OR2_X1    g453(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n309), .A2(new_n632), .A3(new_n427), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n487), .B1(new_n466), .B2(new_n485), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n490), .B1(new_n643), .B2(KEYINPUT93), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT93), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n466), .A2(new_n485), .A3(new_n645), .A4(new_n487), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n379), .A2(new_n390), .ZN(new_n648));
  INV_X1    g462(.A(new_n393), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n379), .A2(new_n390), .A3(new_n393), .ZN(new_n651));
  AOI21_X1  g465(.A(G902), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT96), .B(G478), .Z(new_n653));
  NOR2_X1   g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g468(.A(KEYINPUT33), .B1(new_n650), .B2(new_n651), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT94), .ZN(new_n656));
  OAI211_X1 g470(.A(KEYINPUT33), .B(new_n651), .C1(new_n395), .C2(new_n656), .ZN(new_n657));
  AND2_X1   g471(.A1(new_n395), .A2(new_n656), .ZN(new_n658));
  OAI21_X1  g472(.A(KEYINPUT95), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n650), .A2(KEYINPUT94), .ZN(new_n660));
  AND2_X1   g474(.A1(new_n651), .A2(KEYINPUT33), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT95), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n395), .A2(new_n656), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n660), .A2(new_n661), .A3(new_n662), .A4(new_n663), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n655), .B1(new_n659), .B2(new_n664), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n294), .A2(G478), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n654), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n667), .A2(new_n421), .A3(new_n411), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n647), .A2(new_n496), .A3(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT97), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n429), .B1(new_n644), .B2(new_n646), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n672), .A2(KEYINPUT97), .A3(new_n668), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n642), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT34), .B(G104), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G6));
  INV_X1    g491(.A(new_n411), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n366), .B1(new_n349), .B2(new_n354), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(new_n369), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n680), .A2(new_n418), .ZN(new_n681));
  AND4_X1   g495(.A1(new_n678), .A2(new_n672), .A3(new_n401), .A4(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n642), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT99), .B(G107), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT98), .B(KEYINPUT35), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G9));
  INV_X1    g501(.A(KEYINPUT100), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n619), .A2(KEYINPUT36), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n615), .B(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n630), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n688), .B1(new_n629), .B2(new_n692), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n627), .B1(new_n626), .B2(new_n294), .ZN(new_n694));
  NOR4_X1   g508(.A1(new_n624), .A2(new_n625), .A3(G902), .A4(new_n597), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n595), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n696), .A2(KEYINPUT100), .A3(new_n691), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n693), .A2(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n637), .A2(new_n639), .A3(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n494), .A2(new_n499), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(KEYINPUT37), .B(G110), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(KEYINPUT101), .B(KEYINPUT102), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G12));
  NAND3_X1  g519(.A1(new_n309), .A2(new_n427), .A3(new_n672), .ZN(new_n706));
  INV_X1    g520(.A(G900), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n408), .B1(new_n707), .B2(new_n410), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n681), .A2(new_n401), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n698), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n706), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n712), .A2(new_n590), .A3(new_n594), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G128), .ZN(G30));
  AND2_X1   g528(.A1(new_n309), .A2(new_n427), .ZN(new_n715));
  XNOR2_X1  g529(.A(KEYINPUT103), .B(KEYINPUT39), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n708), .B(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  OR2_X1    g532(.A1(new_n718), .A2(KEYINPUT40), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(KEYINPUT40), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n556), .B1(new_n525), .B2(new_n552), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n294), .B1(new_n572), .B2(new_n721), .ZN(new_n722));
  AOI22_X1  g536(.A1(new_n588), .A2(new_n504), .B1(G472), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n592), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n495), .B(KEYINPUT38), .ZN(new_n725));
  INV_X1    g539(.A(new_n401), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n421), .A2(new_n726), .ZN(new_n727));
  AND4_X1   g541(.A1(new_n496), .A2(new_n725), .A3(new_n699), .A4(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n719), .A2(new_n720), .A3(new_n724), .A4(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(new_n327), .ZN(G45));
  OR2_X1    g544(.A1(new_n667), .A2(new_n421), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n731), .A2(new_n708), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n698), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n706), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n734), .A2(new_n590), .A3(new_n594), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G146), .ZN(G48));
  INV_X1    g550(.A(new_n632), .ZN(new_n737));
  INV_X1    g551(.A(new_n425), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n265), .B1(new_n272), .B2(new_n282), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n307), .B1(new_n739), .B2(new_n269), .ZN(new_n740));
  OAI21_X1  g554(.A(G469), .B1(new_n740), .B2(G902), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT104), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n308), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  OAI211_X1 g557(.A(KEYINPUT104), .B(G469), .C1(new_n740), .C2(G902), .ZN(new_n744));
  AOI211_X1 g558(.A(new_n737), .B(new_n738), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n674), .A2(new_n745), .A3(new_n590), .A4(new_n594), .ZN(new_n746));
  XNOR2_X1  g560(.A(KEYINPUT41), .B(G113), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(G15));
  NAND4_X1  g562(.A1(new_n745), .A2(new_n590), .A3(new_n594), .A4(new_n682), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G116), .ZN(G18));
  NAND2_X1  g564(.A1(new_n743), .A2(new_n744), .ZN(new_n751));
  AND3_X1   g565(.A1(new_n751), .A2(new_n425), .A3(new_n672), .ZN(new_n752));
  AND2_X1   g566(.A1(new_n424), .A2(new_n698), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n752), .A2(new_n590), .A3(new_n594), .A4(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G119), .ZN(G21));
  AOI21_X1  g569(.A(new_n738), .B1(new_n743), .B2(new_n744), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n756), .A2(new_n678), .ZN(new_n757));
  OR3_X1    g571(.A1(new_n421), .A2(KEYINPUT106), .A3(new_n726), .ZN(new_n758));
  OAI21_X1  g572(.A(KEYINPUT106), .B1(new_n421), .B2(new_n726), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n760), .A2(new_n672), .ZN(new_n761));
  AOI22_X1  g575(.A1(new_n572), .A2(new_n505), .B1(new_n566), .B2(new_n565), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n502), .B1(new_n762), .B2(new_n584), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n588), .A2(new_n294), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n763), .B1(new_n764), .B2(G472), .ZN(new_n765));
  AOI21_X1  g579(.A(KEYINPUT105), .B1(new_n765), .B2(new_n632), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT105), .ZN(new_n767));
  NOR4_X1   g581(.A1(new_n637), .A2(new_n767), .A3(new_n737), .A4(new_n763), .ZN(new_n768));
  OAI211_X1 g582(.A(new_n757), .B(new_n761), .C1(new_n766), .C2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G122), .ZN(G24));
  NOR3_X1   g584(.A1(new_n637), .A2(new_n699), .A3(new_n763), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n771), .A2(new_n672), .A3(new_n732), .A4(new_n756), .ZN(new_n772));
  XOR2_X1   g586(.A(KEYINPUT107), .B(G125), .Z(new_n773));
  XNOR2_X1  g587(.A(new_n772), .B(new_n773), .ZN(G27));
  AND2_X1   g588(.A1(new_n574), .A2(new_n581), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n737), .B1(new_n775), .B2(new_n592), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n302), .A2(G469), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n738), .B1(new_n308), .B2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT108), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n779), .B1(new_n495), .B2(new_n429), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n489), .A2(KEYINPUT108), .A3(new_n496), .A4(new_n490), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n732), .A2(new_n778), .A3(new_n780), .A4(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n776), .A2(new_n783), .A3(KEYINPUT110), .A4(KEYINPUT42), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT110), .ZN(new_n785));
  OAI211_X1 g599(.A(KEYINPUT42), .B(new_n632), .C1(new_n582), .C2(new_n589), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n785), .B1(new_n786), .B2(new_n782), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n784), .A2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(KEYINPUT109), .B(KEYINPUT42), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n790), .B1(new_n633), .B2(new_n782), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G131), .ZN(G33));
  AND4_X1   g607(.A1(new_n710), .A2(new_n778), .A3(new_n780), .A4(new_n781), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n794), .A2(new_n590), .A3(new_n594), .A4(new_n632), .ZN(new_n795));
  XOR2_X1   g609(.A(KEYINPUT111), .B(G134), .Z(new_n796));
  XNOR2_X1  g610(.A(new_n795), .B(new_n796), .ZN(G36));
  AOI21_X1  g611(.A(KEYINPUT45), .B1(new_n283), .B2(new_n290), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT112), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n283), .A2(new_n290), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT45), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n799), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n283), .A2(new_n290), .A3(KEYINPUT112), .A4(KEYINPUT45), .ZN(new_n803));
  AOI211_X1 g617(.A(new_n292), .B(new_n798), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n292), .A2(new_n294), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(KEYINPUT46), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT46), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n808), .B1(new_n804), .B2(new_n805), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n807), .A2(new_n308), .A3(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n810), .A2(new_n425), .A3(new_n717), .ZN(new_n811));
  INV_X1    g625(.A(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT44), .ZN(new_n813));
  INV_X1    g627(.A(new_n421), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n814), .A2(new_n667), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(KEYINPUT43), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(new_n698), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n637), .A2(new_n639), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n813), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n640), .A2(KEYINPUT44), .A3(new_n698), .A4(new_n816), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n780), .A2(new_n781), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n819), .A2(new_n820), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n812), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(G137), .ZN(G39));
  NAND3_X1  g639(.A1(new_n822), .A2(new_n737), .A3(new_n732), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n826), .B1(new_n590), .B2(new_n594), .ZN(new_n827));
  XNOR2_X1  g641(.A(KEYINPUT113), .B(KEYINPUT47), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n810), .A2(new_n425), .A3(new_n829), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n810), .A2(new_n425), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT113), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n832), .A2(KEYINPUT47), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n827), .B(new_n830), .C1(new_n831), .C2(new_n833), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(G140), .ZN(G42));
  XOR2_X1   g649(.A(new_n751), .B(KEYINPUT49), .Z(new_n836));
  NAND4_X1  g650(.A1(new_n815), .A2(new_n632), .A3(new_n427), .A4(new_n496), .ZN(new_n837));
  OR4_X1    g651(.A1(new_n724), .A2(new_n836), .A3(new_n725), .A4(new_n837), .ZN(new_n838));
  OR2_X1    g652(.A1(G952), .A2(G953), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n816), .A2(new_n408), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n840), .A2(new_n756), .A3(new_n822), .ZN(new_n841));
  INV_X1    g655(.A(new_n776), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(KEYINPUT48), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n840), .B1(new_n766), .B2(new_n768), .ZN(new_n845));
  INV_X1    g659(.A(new_n752), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n724), .A2(new_n737), .A3(new_n407), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n848), .A2(new_n425), .A3(new_n751), .A4(new_n822), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n405), .B1(new_n849), .B2(new_n731), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n844), .A2(new_n847), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT50), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n725), .A2(new_n496), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(new_n756), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n855), .A2(KEYINPUT117), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n853), .A2(KEYINPUT117), .A3(new_n756), .ZN(new_n857));
  OR4_X1    g671(.A1(new_n852), .A2(new_n856), .A3(new_n845), .A4(new_n857), .ZN(new_n858));
  XOR2_X1   g672(.A(new_n854), .B(KEYINPUT117), .Z(new_n859));
  OAI21_X1  g673(.A(new_n852), .B1(new_n859), .B2(new_n845), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n667), .A2(new_n421), .ZN(new_n862));
  INV_X1    g676(.A(new_n771), .ZN(new_n863));
  OAI22_X1  g677(.A1(new_n849), .A2(new_n862), .B1(new_n841), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n751), .A2(new_n426), .ZN(new_n865));
  INV_X1    g679(.A(new_n830), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n833), .B1(new_n810), .B2(new_n425), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n865), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n845), .A2(new_n821), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n864), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT51), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n861), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n871), .B1(new_n861), .B2(new_n870), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n851), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n754), .A2(new_n749), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT114), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n652), .A2(new_n399), .ZN(new_n877));
  INV_X1    g691(.A(new_n400), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n398), .A2(KEYINPUT114), .A3(new_n400), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n731), .B1(new_n814), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n882), .A2(new_n678), .A3(new_n491), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n640), .A2(new_n883), .A3(new_n641), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n494), .A2(new_n499), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n590), .A2(new_n594), .A3(new_n632), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n884), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n746), .A2(new_n701), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n875), .A2(new_n887), .A3(new_n888), .A4(new_n769), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n881), .A2(new_n680), .A3(new_n418), .A4(new_n709), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n890), .B1(new_n693), .B2(new_n697), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n309), .A2(new_n891), .A3(new_n427), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n892), .A2(new_n821), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n893), .A2(new_n590), .A3(new_n594), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n783), .A2(new_n771), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n795), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(new_n790), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n897), .B1(new_n886), .B2(new_n783), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n896), .B1(new_n898), .B2(new_n788), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n889), .A2(new_n899), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n629), .A2(new_n692), .A3(new_n708), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n778), .A2(KEYINPUT115), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(KEYINPUT115), .B1(new_n778), .B2(new_n901), .ZN(new_n903));
  OAI211_X1 g717(.A(new_n724), .B(new_n761), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n735), .A2(new_n713), .A3(new_n772), .A4(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT52), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI211_X1 g721(.A(new_n590), .B(new_n594), .C1(new_n734), .C2(new_n712), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n908), .A2(KEYINPUT52), .A3(new_n772), .A4(new_n904), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(KEYINPUT53), .B1(new_n900), .B2(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n769), .A2(new_n749), .A3(new_n754), .ZN(new_n912));
  INV_X1    g726(.A(new_n883), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n913), .A2(new_n632), .A3(new_n715), .A4(new_n818), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n914), .B1(new_n500), .B2(new_n633), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n746), .A2(new_n701), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n912), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n795), .A2(new_n894), .A3(new_n895), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n918), .B1(new_n789), .B2(new_n791), .ZN(new_n919));
  AND4_X1   g733(.A1(KEYINPUT53), .A2(new_n917), .A3(new_n910), .A4(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(KEYINPUT54), .B1(new_n911), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n917), .A2(new_n910), .A3(new_n919), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT53), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n900), .A2(KEYINPUT53), .A3(new_n910), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT54), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n921), .A2(KEYINPUT116), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n924), .A2(new_n925), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT116), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n929), .A2(new_n930), .A3(KEYINPUT54), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n874), .B1(new_n928), .B2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT118), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n839), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  AOI211_X1 g748(.A(KEYINPUT118), .B(new_n874), .C1(new_n928), .C2(new_n931), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n838), .B1(new_n934), .B2(new_n935), .ZN(G75));
  NOR2_X1   g750(.A1(new_n267), .A2(G952), .ZN(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n911), .A2(new_n920), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n939), .A2(new_n294), .ZN(new_n940));
  AOI21_X1  g754(.A(KEYINPUT56), .B1(new_n940), .B2(G210), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n457), .A2(new_n459), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(new_n465), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT55), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n938), .B1(new_n941), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n946), .B1(new_n941), .B2(new_n945), .ZN(G51));
  INV_X1    g761(.A(KEYINPUT119), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n921), .A2(new_n948), .A3(new_n927), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n929), .A2(KEYINPUT119), .A3(KEYINPUT54), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n805), .B(KEYINPUT57), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n952), .B1(new_n306), .B2(new_n307), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n940), .A2(new_n804), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n937), .B1(new_n953), .B2(new_n954), .ZN(G54));
  NAND3_X1  g769(.A1(new_n940), .A2(KEYINPUT58), .A3(G475), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n956), .A2(new_n364), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n956), .A2(new_n364), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n957), .A2(new_n958), .A3(new_n937), .ZN(G60));
  NAND2_X1  g773(.A1(G478), .A2(G902), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(KEYINPUT59), .Z(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n949), .A2(new_n665), .A3(new_n950), .A4(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(new_n938), .ZN(new_n964));
  INV_X1    g778(.A(new_n665), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n928), .A2(new_n931), .A3(new_n962), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n964), .B1(new_n965), .B2(new_n966), .ZN(G63));
  NAND2_X1  g781(.A1(G217), .A2(G902), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(KEYINPUT60), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n969), .B1(new_n924), .B2(new_n925), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n970), .A2(new_n626), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n971), .A2(new_n937), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT120), .ZN(new_n973));
  AND3_X1   g787(.A1(new_n970), .A2(new_n973), .A3(new_n690), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n973), .B1(new_n970), .B2(new_n690), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n972), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT61), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n972), .B(KEYINPUT61), .C1(new_n974), .C2(new_n975), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(G66));
  OAI21_X1  g794(.A(G953), .B1(new_n409), .B2(new_n463), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(KEYINPUT121), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n982), .B1(new_n917), .B2(G953), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(KEYINPUT122), .ZN(new_n984));
  INV_X1    g798(.A(G898), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n942), .B1(new_n985), .B2(G953), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n984), .B(new_n986), .ZN(G69));
  NAND2_X1  g801(.A1(new_n707), .A2(G953), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(KEYINPUT125), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n831), .A2(new_n717), .A3(new_n761), .A4(new_n776), .ZN(new_n990));
  AND2_X1   g804(.A1(new_n908), .A2(new_n772), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n990), .A2(new_n824), .A3(new_n795), .A4(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n834), .A2(new_n792), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n989), .B1(new_n994), .B2(G953), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n991), .A2(new_n729), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n996), .A2(KEYINPUT62), .ZN(new_n997));
  AND4_X1   g811(.A1(new_n715), .A2(new_n822), .A3(new_n717), .A4(new_n882), .ZN(new_n998));
  AOI22_X1  g812(.A1(new_n812), .A2(new_n823), .B1(new_n886), .B2(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT62), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n991), .A2(new_n1000), .A3(new_n729), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n997), .A2(new_n834), .A3(new_n999), .A4(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT123), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n537), .B1(new_n535), .B2(new_n534), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n322), .A2(new_n323), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1004), .B(new_n1005), .ZN(new_n1006));
  AOI22_X1  g820(.A1(new_n1002), .A2(new_n267), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g821(.A(KEYINPUT123), .B1(new_n1002), .B2(new_n267), .ZN(new_n1008));
  OAI22_X1  g822(.A1(new_n995), .A2(new_n1007), .B1(new_n1008), .B2(new_n1006), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1009), .A2(KEYINPUT124), .ZN(new_n1010));
  INV_X1    g824(.A(KEYINPUT124), .ZN(new_n1011));
  OAI221_X1 g825(.A(new_n1011), .B1(new_n1008), .B2(new_n1006), .C1(new_n995), .C2(new_n1007), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n267), .B1(G227), .B2(G900), .ZN(new_n1013));
  AND3_X1   g827(.A1(new_n1010), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1013), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n1014), .A2(new_n1015), .ZN(G72));
  NAND2_X1  g830(.A1(G472), .A2(G902), .ZN(new_n1017));
  XOR2_X1   g831(.A(new_n1017), .B(KEYINPUT63), .Z(new_n1018));
  INV_X1    g832(.A(new_n1018), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1019), .B1(new_n994), .B2(new_n917), .ZN(new_n1020));
  XOR2_X1   g834(.A(new_n577), .B(KEYINPUT126), .Z(new_n1021));
  NAND2_X1  g835(.A1(new_n1021), .A2(new_n555), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n938), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g837(.A(new_n1023), .B(KEYINPUT127), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n572), .B1(new_n577), .B2(new_n555), .ZN(new_n1025));
  NOR3_X1   g839(.A1(new_n939), .A2(new_n1019), .A3(new_n1025), .ZN(new_n1026));
  OR2_X1    g840(.A1(new_n1002), .A2(new_n889), .ZN(new_n1027));
  AOI211_X1 g841(.A(new_n555), .B(new_n1021), .C1(new_n1027), .C2(new_n1018), .ZN(new_n1028));
  NOR3_X1   g842(.A1(new_n1024), .A2(new_n1026), .A3(new_n1028), .ZN(G57));
endmodule


