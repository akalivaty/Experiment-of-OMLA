

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583;

  XNOR2_X1 U325 ( .A(n421), .B(n420), .ZN(n560) );
  NOR2_X1 U326 ( .A1(n560), .A2(n429), .ZN(n430) );
  XNOR2_X1 U327 ( .A(n385), .B(n384), .ZN(n571) );
  NOR2_X1 U328 ( .A1(n464), .A2(n564), .ZN(n453) );
  XOR2_X1 U329 ( .A(G162GAT), .B(G218GAT), .Z(n293) );
  XOR2_X1 U330 ( .A(KEYINPUT13), .B(KEYINPUT72), .Z(n294) );
  XNOR2_X1 U331 ( .A(n406), .B(n293), .ZN(n410) );
  XNOR2_X1 U332 ( .A(n410), .B(n409), .ZN(n415) );
  XNOR2_X1 U333 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U334 ( .A(KEYINPUT36), .B(n560), .Z(n580) );
  XNOR2_X1 U335 ( .A(n433), .B(KEYINPUT48), .ZN(n545) );
  NOR2_X1 U336 ( .A1(n524), .A2(n454), .ZN(n561) );
  XNOR2_X1 U337 ( .A(n475), .B(KEYINPUT41), .ZN(n549) );
  XNOR2_X1 U338 ( .A(n317), .B(n316), .ZN(n524) );
  XNOR2_X1 U339 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U340 ( .A(n458), .B(n457), .ZN(G1349GAT) );
  XOR2_X1 U341 ( .A(KEYINPUT90), .B(KEYINPUT65), .Z(n296) );
  XNOR2_X1 U342 ( .A(G120GAT), .B(G71GAT), .ZN(n295) );
  XNOR2_X1 U343 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U344 ( .A(G183GAT), .B(KEYINPUT89), .Z(n298) );
  XNOR2_X1 U345 ( .A(G15GAT), .B(G176GAT), .ZN(n297) );
  XNOR2_X1 U346 ( .A(n298), .B(n297), .ZN(n299) );
  XNOR2_X1 U347 ( .A(n300), .B(n299), .ZN(n317) );
  XOR2_X1 U348 ( .A(G127GAT), .B(KEYINPUT91), .Z(n302) );
  XNOR2_X1 U349 ( .A(G43GAT), .B(G99GAT), .ZN(n301) );
  XNOR2_X1 U350 ( .A(n302), .B(n301), .ZN(n304) );
  XOR2_X1 U351 ( .A(G134GAT), .B(G190GAT), .Z(n303) );
  XNOR2_X1 U352 ( .A(n304), .B(n303), .ZN(n313) );
  XOR2_X1 U353 ( .A(KEYINPUT94), .B(KEYINPUT20), .Z(n311) );
  XNOR2_X1 U354 ( .A(KEYINPUT17), .B(KEYINPUT19), .ZN(n305) );
  XNOR2_X1 U355 ( .A(n305), .B(KEYINPUT18), .ZN(n306) );
  XOR2_X1 U356 ( .A(n306), .B(KEYINPUT93), .Z(n308) );
  XNOR2_X1 U357 ( .A(G169GAT), .B(KEYINPUT92), .ZN(n307) );
  XNOR2_X1 U358 ( .A(n308), .B(n307), .ZN(n339) );
  XNOR2_X1 U359 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n309) );
  XNOR2_X1 U360 ( .A(n309), .B(KEYINPUT88), .ZN(n439) );
  XNOR2_X1 U361 ( .A(n339), .B(n439), .ZN(n310) );
  XNOR2_X1 U362 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U363 ( .A(n313), .B(n312), .ZN(n315) );
  NAND2_X1 U364 ( .A1(G227GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U365 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U366 ( .A(KEYINPUT96), .B(KEYINPUT24), .Z(n319) );
  NAND2_X1 U367 ( .A1(G228GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U368 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U369 ( .A(n320), .B(KEYINPUT97), .Z(n326) );
  XOR2_X1 U370 ( .A(G211GAT), .B(KEYINPUT21), .Z(n322) );
  XNOR2_X1 U371 ( .A(G197GAT), .B(G218GAT), .ZN(n321) );
  XNOR2_X1 U372 ( .A(n322), .B(n321), .ZN(n347) );
  XOR2_X1 U373 ( .A(G78GAT), .B(G204GAT), .Z(n324) );
  XNOR2_X1 U374 ( .A(G106GAT), .B(KEYINPUT74), .ZN(n323) );
  XNOR2_X1 U375 ( .A(n324), .B(n323), .ZN(n377) );
  XNOR2_X1 U376 ( .A(n347), .B(n377), .ZN(n325) );
  XNOR2_X1 U377 ( .A(n326), .B(n325), .ZN(n330) );
  XOR2_X1 U378 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n328) );
  XNOR2_X1 U379 ( .A(G50GAT), .B(KEYINPUT98), .ZN(n327) );
  XNOR2_X1 U380 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U381 ( .A(n330), .B(n329), .Z(n338) );
  XOR2_X1 U382 ( .A(KEYINPUT3), .B(G162GAT), .Z(n332) );
  XNOR2_X1 U383 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n331) );
  XNOR2_X1 U384 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U385 ( .A(G141GAT), .B(n333), .Z(n451) );
  XOR2_X1 U386 ( .A(KEYINPUT99), .B(KEYINPUT95), .Z(n335) );
  XNOR2_X1 U387 ( .A(G22GAT), .B(G148GAT), .ZN(n334) );
  XNOR2_X1 U388 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U389 ( .A(n451), .B(n336), .ZN(n337) );
  XNOR2_X1 U390 ( .A(n338), .B(n337), .ZN(n464) );
  XOR2_X1 U391 ( .A(G36GAT), .B(G190GAT), .Z(n411) );
  XOR2_X1 U392 ( .A(G8GAT), .B(G183GAT), .Z(n395) );
  XOR2_X1 U393 ( .A(n395), .B(KEYINPUT103), .Z(n341) );
  XNOR2_X1 U394 ( .A(n339), .B(G204GAT), .ZN(n340) );
  XNOR2_X1 U395 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U396 ( .A(n411), .B(n342), .Z(n344) );
  NAND2_X1 U397 ( .A1(G226GAT), .A2(G233GAT), .ZN(n343) );
  XNOR2_X1 U398 ( .A(n344), .B(n343), .ZN(n349) );
  XOR2_X1 U399 ( .A(G64GAT), .B(KEYINPUT77), .Z(n346) );
  XNOR2_X1 U400 ( .A(G176GAT), .B(G92GAT), .ZN(n345) );
  XNOR2_X1 U401 ( .A(n346), .B(n345), .ZN(n381) );
  XOR2_X1 U402 ( .A(n347), .B(n381), .Z(n348) );
  XNOR2_X1 U403 ( .A(n349), .B(n348), .ZN(n521) );
  XOR2_X1 U404 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n351) );
  XNOR2_X1 U405 ( .A(KEYINPUT71), .B(KEYINPUT66), .ZN(n350) );
  XNOR2_X1 U406 ( .A(n351), .B(n350), .ZN(n365) );
  XOR2_X1 U407 ( .A(G113GAT), .B(G141GAT), .Z(n353) );
  XNOR2_X1 U408 ( .A(G169GAT), .B(G197GAT), .ZN(n352) );
  XNOR2_X1 U409 ( .A(n353), .B(n352), .ZN(n357) );
  XOR2_X1 U410 ( .A(KEYINPUT67), .B(KEYINPUT70), .Z(n355) );
  XNOR2_X1 U411 ( .A(G8GAT), .B(G1GAT), .ZN(n354) );
  XNOR2_X1 U412 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U413 ( .A(n357), .B(n356), .Z(n363) );
  XNOR2_X1 U414 ( .A(G22GAT), .B(G15GAT), .ZN(n358) );
  XNOR2_X1 U415 ( .A(n358), .B(KEYINPUT69), .ZN(n392) );
  XOR2_X1 U416 ( .A(G36GAT), .B(n392), .Z(n360) );
  NAND2_X1 U417 ( .A1(G229GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U418 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U419 ( .A(G29GAT), .B(n361), .ZN(n362) );
  XNOR2_X1 U420 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U421 ( .A(n365), .B(n364), .ZN(n369) );
  XOR2_X1 U422 ( .A(KEYINPUT68), .B(KEYINPUT8), .Z(n367) );
  XNOR2_X1 U423 ( .A(G50GAT), .B(G43GAT), .ZN(n366) );
  XNOR2_X1 U424 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U425 ( .A(KEYINPUT7), .B(n368), .ZN(n416) );
  XOR2_X1 U426 ( .A(n369), .B(n416), .Z(n505) );
  INV_X1 U427 ( .A(n505), .ZN(n566) );
  XNOR2_X1 U428 ( .A(G71GAT), .B(KEYINPUT73), .ZN(n370) );
  XNOR2_X1 U429 ( .A(n294), .B(n370), .ZN(n391) );
  XOR2_X1 U430 ( .A(n391), .B(KEYINPUT32), .Z(n372) );
  XOR2_X1 U431 ( .A(G99GAT), .B(G85GAT), .Z(n406) );
  XNOR2_X1 U432 ( .A(n406), .B(KEYINPUT78), .ZN(n371) );
  XNOR2_X1 U433 ( .A(n372), .B(n371), .ZN(n376) );
  XOR2_X1 U434 ( .A(KEYINPUT75), .B(KEYINPUT33), .Z(n374) );
  XNOR2_X1 U435 ( .A(KEYINPUT31), .B(KEYINPUT79), .ZN(n373) );
  XNOR2_X1 U436 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U437 ( .A(n376), .B(n375), .Z(n385) );
  XOR2_X1 U438 ( .A(n377), .B(KEYINPUT76), .Z(n379) );
  NAND2_X1 U439 ( .A1(G230GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U440 ( .A(n379), .B(n378), .ZN(n383) );
  XNOR2_X1 U441 ( .A(G120GAT), .B(G148GAT), .ZN(n380) );
  XNOR2_X1 U442 ( .A(n380), .B(G57GAT), .ZN(n438) );
  XNOR2_X1 U443 ( .A(n438), .B(n381), .ZN(n382) );
  XOR2_X1 U444 ( .A(KEYINPUT86), .B(KEYINPUT84), .Z(n387) );
  XNOR2_X1 U445 ( .A(G57GAT), .B(KEYINPUT85), .ZN(n386) );
  XNOR2_X1 U446 ( .A(n387), .B(n386), .ZN(n403) );
  XOR2_X1 U447 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n389) );
  NAND2_X1 U448 ( .A1(G231GAT), .A2(G233GAT), .ZN(n388) );
  XNOR2_X1 U449 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U450 ( .A(n390), .B(KEYINPUT14), .Z(n394) );
  XNOR2_X1 U451 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U452 ( .A(n394), .B(n393), .ZN(n399) );
  XOR2_X1 U453 ( .A(n395), .B(G64GAT), .Z(n397) );
  XOR2_X1 U454 ( .A(G1GAT), .B(G127GAT), .Z(n446) );
  XNOR2_X1 U455 ( .A(G78GAT), .B(n446), .ZN(n396) );
  XNOR2_X1 U456 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U457 ( .A(n399), .B(n398), .Z(n401) );
  XNOR2_X1 U458 ( .A(G155GAT), .B(G211GAT), .ZN(n400) );
  XNOR2_X1 U459 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U460 ( .A(n403), .B(n402), .Z(n536) );
  XOR2_X1 U461 ( .A(KEYINPUT82), .B(KEYINPUT9), .Z(n405) );
  XNOR2_X1 U462 ( .A(G106GAT), .B(KEYINPUT10), .ZN(n404) );
  XNOR2_X1 U463 ( .A(n405), .B(n404), .ZN(n421) );
  XOR2_X1 U464 ( .A(KEYINPUT11), .B(KEYINPUT83), .Z(n408) );
  XNOR2_X1 U465 ( .A(G92GAT), .B(KEYINPUT64), .ZN(n407) );
  XNOR2_X1 U466 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U467 ( .A(n411), .B(KEYINPUT81), .Z(n413) );
  NAND2_X1 U468 ( .A1(G232GAT), .A2(G233GAT), .ZN(n412) );
  XNOR2_X1 U469 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U470 ( .A(n415), .B(n414), .Z(n419) );
  INV_X1 U471 ( .A(n416), .ZN(n417) );
  XOR2_X1 U472 ( .A(G29GAT), .B(G134GAT), .Z(n447) );
  XNOR2_X1 U473 ( .A(n417), .B(n447), .ZN(n418) );
  XNOR2_X1 U474 ( .A(n419), .B(n418), .ZN(n420) );
  NOR2_X1 U475 ( .A1(n536), .A2(n580), .ZN(n422) );
  XOR2_X1 U476 ( .A(KEYINPUT45), .B(n422), .Z(n423) );
  NOR2_X1 U477 ( .A1(n571), .A2(n423), .ZN(n424) );
  XOR2_X1 U478 ( .A(KEYINPUT118), .B(n424), .Z(n425) );
  NOR2_X1 U479 ( .A1(n566), .A2(n425), .ZN(n432) );
  XOR2_X1 U480 ( .A(KEYINPUT46), .B(KEYINPUT117), .Z(n427) );
  INV_X1 U481 ( .A(n571), .ZN(n475) );
  NAND2_X1 U482 ( .A1(n549), .A2(n566), .ZN(n426) );
  XNOR2_X1 U483 ( .A(n427), .B(n426), .ZN(n428) );
  NAND2_X1 U484 ( .A1(n536), .A2(n428), .ZN(n429) );
  XOR2_X1 U485 ( .A(KEYINPUT47), .B(n430), .Z(n431) );
  NOR2_X1 U486 ( .A1(n432), .A2(n431), .ZN(n433) );
  NOR2_X1 U487 ( .A1(n521), .A2(n545), .ZN(n434) );
  XNOR2_X1 U488 ( .A(n434), .B(KEYINPUT54), .ZN(n452) );
  XOR2_X1 U489 ( .A(KEYINPUT1), .B(KEYINPUT5), .Z(n436) );
  NAND2_X1 U490 ( .A1(G225GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U491 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U492 ( .A(n437), .B(KEYINPUT100), .Z(n441) );
  XNOR2_X1 U493 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U494 ( .A(n441), .B(n440), .ZN(n445) );
  XOR2_X1 U495 ( .A(KEYINPUT101), .B(KEYINPUT4), .Z(n443) );
  XNOR2_X1 U496 ( .A(G85GAT), .B(KEYINPUT6), .ZN(n442) );
  XNOR2_X1 U497 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U498 ( .A(n445), .B(n444), .Z(n449) );
  XNOR2_X1 U499 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U500 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U501 ( .A(n451), .B(n450), .ZN(n468) );
  XNOR2_X1 U502 ( .A(KEYINPUT102), .B(n468), .ZN(n544) );
  NAND2_X1 U503 ( .A1(n452), .A2(n544), .ZN(n564) );
  XNOR2_X1 U504 ( .A(n453), .B(KEYINPUT55), .ZN(n454) );
  NAND2_X1 U505 ( .A1(n561), .A2(n549), .ZN(n458) );
  XOR2_X1 U506 ( .A(KEYINPUT56), .B(KEYINPUT122), .Z(n456) );
  XNOR2_X1 U507 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n455) );
  XNOR2_X1 U508 ( .A(KEYINPUT27), .B(KEYINPUT104), .ZN(n459) );
  XNOR2_X1 U509 ( .A(n459), .B(n521), .ZN(n466) );
  INV_X1 U510 ( .A(n544), .ZN(n478) );
  XNOR2_X1 U511 ( .A(n464), .B(KEYINPUT28), .ZN(n487) );
  INV_X1 U512 ( .A(n487), .ZN(n527) );
  NAND2_X1 U513 ( .A1(n478), .A2(n527), .ZN(n460) );
  NOR2_X1 U514 ( .A1(n466), .A2(n460), .ZN(n531) );
  XOR2_X1 U515 ( .A(n531), .B(KEYINPUT105), .Z(n461) );
  NAND2_X1 U516 ( .A1(n461), .A2(n524), .ZN(n471) );
  NOR2_X1 U517 ( .A1(n524), .A2(n521), .ZN(n462) );
  NOR2_X1 U518 ( .A1(n464), .A2(n462), .ZN(n463) );
  XNOR2_X1 U519 ( .A(n463), .B(KEYINPUT25), .ZN(n467) );
  NAND2_X1 U520 ( .A1(n464), .A2(n524), .ZN(n465) );
  XNOR2_X1 U521 ( .A(n465), .B(KEYINPUT26), .ZN(n565) );
  OR2_X1 U522 ( .A1(n565), .A2(n466), .ZN(n547) );
  NAND2_X1 U523 ( .A1(n467), .A2(n547), .ZN(n469) );
  NAND2_X1 U524 ( .A1(n469), .A2(n468), .ZN(n470) );
  NAND2_X1 U525 ( .A1(n471), .A2(n470), .ZN(n490) );
  NOR2_X1 U526 ( .A1(n560), .A2(n536), .ZN(n472) );
  XNOR2_X1 U527 ( .A(n472), .B(KEYINPUT16), .ZN(n473) );
  XOR2_X1 U528 ( .A(KEYINPUT87), .B(n473), .Z(n474) );
  AND2_X1 U529 ( .A1(n490), .A2(n474), .ZN(n507) );
  NAND2_X1 U530 ( .A1(n566), .A2(n475), .ZN(n476) );
  XOR2_X1 U531 ( .A(KEYINPUT80), .B(n476), .Z(n494) );
  NAND2_X1 U532 ( .A1(n507), .A2(n494), .ZN(n477) );
  XOR2_X1 U533 ( .A(KEYINPUT106), .B(n477), .Z(n488) );
  NAND2_X1 U534 ( .A1(n488), .A2(n478), .ZN(n481) );
  XOR2_X1 U535 ( .A(G1GAT), .B(KEYINPUT34), .Z(n479) );
  XNOR2_X1 U536 ( .A(KEYINPUT107), .B(n479), .ZN(n480) );
  XNOR2_X1 U537 ( .A(n481), .B(n480), .ZN(G1324GAT) );
  XNOR2_X1 U538 ( .A(G8GAT), .B(KEYINPUT108), .ZN(n484) );
  INV_X1 U539 ( .A(n521), .ZN(n482) );
  NAND2_X1 U540 ( .A1(n482), .A2(n488), .ZN(n483) );
  XNOR2_X1 U541 ( .A(n484), .B(n483), .ZN(G1325GAT) );
  XOR2_X1 U542 ( .A(G15GAT), .B(KEYINPUT35), .Z(n486) );
  INV_X1 U543 ( .A(n524), .ZN(n530) );
  NAND2_X1 U544 ( .A1(n488), .A2(n530), .ZN(n485) );
  XNOR2_X1 U545 ( .A(n486), .B(n485), .ZN(G1326GAT) );
  NAND2_X1 U546 ( .A1(n488), .A2(n487), .ZN(n489) );
  XNOR2_X1 U547 ( .A(n489), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U548 ( .A1(n536), .A2(n490), .ZN(n491) );
  NOR2_X1 U549 ( .A1(n580), .A2(n491), .ZN(n493) );
  XNOR2_X1 U550 ( .A(KEYINPUT109), .B(KEYINPUT37), .ZN(n492) );
  XNOR2_X1 U551 ( .A(n493), .B(n492), .ZN(n519) );
  NAND2_X1 U552 ( .A1(n494), .A2(n519), .ZN(n495) );
  XNOR2_X1 U553 ( .A(n495), .B(KEYINPUT110), .ZN(n496) );
  XNOR2_X1 U554 ( .A(KEYINPUT38), .B(n496), .ZN(n503) );
  NOR2_X1 U555 ( .A1(n544), .A2(n503), .ZN(n498) );
  XNOR2_X1 U556 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n497) );
  XNOR2_X1 U557 ( .A(n498), .B(n497), .ZN(G1328GAT) );
  NOR2_X1 U558 ( .A1(n521), .A2(n503), .ZN(n499) );
  XOR2_X1 U559 ( .A(G36GAT), .B(n499), .Z(G1329GAT) );
  NOR2_X1 U560 ( .A1(n524), .A2(n503), .ZN(n501) );
  XNOR2_X1 U561 ( .A(KEYINPUT40), .B(KEYINPUT111), .ZN(n500) );
  XNOR2_X1 U562 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U563 ( .A(G43GAT), .B(n502), .ZN(G1330GAT) );
  NOR2_X1 U564 ( .A1(n527), .A2(n503), .ZN(n504) );
  XOR2_X1 U565 ( .A(G50GAT), .B(n504), .Z(G1331GAT) );
  NAND2_X1 U566 ( .A1(n549), .A2(n505), .ZN(n506) );
  XOR2_X1 U567 ( .A(KEYINPUT112), .B(n506), .Z(n518) );
  NAND2_X1 U568 ( .A1(n507), .A2(n518), .ZN(n515) );
  NOR2_X1 U569 ( .A1(n544), .A2(n515), .ZN(n509) );
  XNOR2_X1 U570 ( .A(KEYINPUT113), .B(KEYINPUT42), .ZN(n508) );
  XNOR2_X1 U571 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U572 ( .A(G57GAT), .B(n510), .ZN(G1332GAT) );
  NOR2_X1 U573 ( .A1(n521), .A2(n515), .ZN(n511) );
  XOR2_X1 U574 ( .A(KEYINPUT114), .B(n511), .Z(n512) );
  XNOR2_X1 U575 ( .A(G64GAT), .B(n512), .ZN(G1333GAT) );
  NOR2_X1 U576 ( .A1(n524), .A2(n515), .ZN(n514) );
  XNOR2_X1 U577 ( .A(G71GAT), .B(KEYINPUT115), .ZN(n513) );
  XNOR2_X1 U578 ( .A(n514), .B(n513), .ZN(G1334GAT) );
  NOR2_X1 U579 ( .A1(n527), .A2(n515), .ZN(n517) );
  XNOR2_X1 U580 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n517), .B(n516), .ZN(G1335GAT) );
  NAND2_X1 U582 ( .A1(n519), .A2(n518), .ZN(n526) );
  NOR2_X1 U583 ( .A1(n544), .A2(n526), .ZN(n520) );
  XOR2_X1 U584 ( .A(G85GAT), .B(n520), .Z(G1336GAT) );
  NOR2_X1 U585 ( .A1(n521), .A2(n526), .ZN(n522) );
  XOR2_X1 U586 ( .A(KEYINPUT116), .B(n522), .Z(n523) );
  XNOR2_X1 U587 ( .A(G92GAT), .B(n523), .ZN(G1337GAT) );
  NOR2_X1 U588 ( .A1(n524), .A2(n526), .ZN(n525) );
  XOR2_X1 U589 ( .A(G99GAT), .B(n525), .Z(G1338GAT) );
  NOR2_X1 U590 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U591 ( .A(KEYINPUT44), .B(n528), .Z(n529) );
  XNOR2_X1 U592 ( .A(G106GAT), .B(n529), .ZN(G1339GAT) );
  NAND2_X1 U593 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U594 ( .A1(n545), .A2(n532), .ZN(n540) );
  NAND2_X1 U595 ( .A1(n566), .A2(n540), .ZN(n533) );
  XNOR2_X1 U596 ( .A(n533), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U597 ( .A(G120GAT), .B(KEYINPUT49), .Z(n535) );
  NAND2_X1 U598 ( .A1(n540), .A2(n549), .ZN(n534) );
  XNOR2_X1 U599 ( .A(n535), .B(n534), .ZN(G1341GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT119), .B(KEYINPUT50), .Z(n538) );
  INV_X1 U601 ( .A(n536), .ZN(n575) );
  NAND2_X1 U602 ( .A1(n540), .A2(n575), .ZN(n537) );
  XNOR2_X1 U603 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U604 ( .A(G127GAT), .B(n539), .ZN(G1342GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT51), .B(KEYINPUT120), .Z(n542) );
  NAND2_X1 U606 ( .A1(n540), .A2(n560), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U608 ( .A(G134GAT), .B(n543), .ZN(G1343GAT) );
  OR2_X1 U609 ( .A1(n545), .A2(n544), .ZN(n546) );
  NOR2_X1 U610 ( .A1(n547), .A2(n546), .ZN(n555) );
  NAND2_X1 U611 ( .A1(n566), .A2(n555), .ZN(n548) );
  XNOR2_X1 U612 ( .A(n548), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT121), .B(KEYINPUT52), .Z(n551) );
  NAND2_X1 U614 ( .A1(n555), .A2(n549), .ZN(n550) );
  XNOR2_X1 U615 ( .A(n551), .B(n550), .ZN(n553) );
  XOR2_X1 U616 ( .A(G148GAT), .B(KEYINPUT53), .Z(n552) );
  XNOR2_X1 U617 ( .A(n553), .B(n552), .ZN(G1345GAT) );
  NAND2_X1 U618 ( .A1(n575), .A2(n555), .ZN(n554) );
  XNOR2_X1 U619 ( .A(n554), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U620 ( .A1(n560), .A2(n555), .ZN(n556) );
  XNOR2_X1 U621 ( .A(n556), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U622 ( .A1(n566), .A2(n561), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n557), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U624 ( .A(G183GAT), .B(KEYINPUT123), .Z(n559) );
  NAND2_X1 U625 ( .A1(n561), .A2(n575), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(G1350GAT) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(KEYINPUT58), .ZN(n563) );
  XNOR2_X1 U629 ( .A(G190GAT), .B(n563), .ZN(G1351GAT) );
  NOR2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n578) );
  NAND2_X1 U631 ( .A1(n566), .A2(n578), .ZN(n570) );
  XOR2_X1 U632 ( .A(KEYINPUT59), .B(KEYINPUT124), .Z(n568) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(G1352GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n573) );
  NAND2_X1 U637 ( .A1(n578), .A2(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n574) );
  XOR2_X1 U639 ( .A(G204GAT), .B(n574), .Z(G1353GAT) );
  NAND2_X1 U640 ( .A1(n575), .A2(n578), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n576), .B(KEYINPUT126), .ZN(n577) );
  XNOR2_X1 U642 ( .A(G211GAT), .B(n577), .ZN(G1354GAT) );
  INV_X1 U643 ( .A(n578), .ZN(n579) );
  NOR2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n582) );
  XNOR2_X1 U645 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(n583), .ZN(G1355GAT) );
endmodule

