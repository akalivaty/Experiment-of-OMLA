//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 0 0 0 0 0 1 0 0 1 0 0 1 1 1 0 0 0 1 0 0 1 1 1 0 0 1 1 0 1 1 1 0 1 1 0 1 0 1 1 1 0 0 0 0 1 1 0 0 0 1 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:56 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n757,
    new_n758, new_n759, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n791, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(G110), .B(G140), .ZN(new_n190));
  INV_X1    g004(.A(G227), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G953), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n190), .B(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  XOR2_X1   g008(.A(KEYINPUT78), .B(KEYINPUT12), .Z(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G143), .ZN(new_n197));
  OAI21_X1  g011(.A(KEYINPUT64), .B1(new_n197), .B2(G146), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT64), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(new_n200), .A3(G143), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n197), .A2(G146), .ZN(new_n202));
  INV_X1    g016(.A(G128), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n203), .A2(KEYINPUT1), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n198), .A2(new_n201), .A3(new_n202), .A4(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n203), .A2(KEYINPUT67), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT67), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G128), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n200), .A2(G143), .ZN(new_n210));
  AOI22_X1  g024(.A1(new_n207), .A2(new_n209), .B1(new_n210), .B2(KEYINPUT1), .ZN(new_n211));
  AND2_X1   g025(.A1(new_n210), .A2(new_n202), .ZN(new_n212));
  OAI21_X1  g026(.A(KEYINPUT68), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n210), .A2(new_n202), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT68), .ZN(new_n215));
  XNOR2_X1  g029(.A(KEYINPUT67), .B(G128), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT1), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n217), .B1(G143), .B2(new_n200), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n214), .B(new_n215), .C1(new_n216), .C2(new_n218), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n206), .B1(new_n213), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n221));
  INV_X1    g035(.A(G104), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n221), .B1(new_n222), .B2(G107), .ZN(new_n223));
  INV_X1    g037(.A(G107), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n224), .A2(KEYINPUT3), .A3(G104), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G101), .ZN(new_n227));
  OAI21_X1  g041(.A(KEYINPUT75), .B1(new_n224), .B2(G104), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT75), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n229), .A2(new_n222), .A3(G107), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n226), .A2(new_n227), .A3(new_n228), .A4(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n222), .A2(G107), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n224), .A2(G104), .ZN(new_n233));
  OAI21_X1  g047(.A(G101), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n231), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n220), .A2(new_n235), .ZN(new_n236));
  AND3_X1   g050(.A1(new_n198), .A2(new_n201), .A3(new_n202), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n218), .A2(new_n203), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n205), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n239), .A2(new_n231), .A3(new_n234), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n236), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(KEYINPUT11), .A2(G134), .ZN(new_n242));
  OAI21_X1  g056(.A(KEYINPUT66), .B1(new_n242), .B2(G137), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT66), .ZN(new_n244));
  INV_X1    g058(.A(G137), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n244), .A2(new_n245), .A3(KEYINPUT11), .A4(G134), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT65), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT11), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n245), .A2(G134), .ZN(new_n251));
  NAND2_X1  g065(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n250), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n245), .A2(G134), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n247), .A2(new_n253), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G131), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n254), .A2(G131), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n247), .A2(new_n253), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n196), .B1(new_n241), .B2(new_n260), .ZN(new_n261));
  AOI22_X1  g075(.A1(new_n248), .A2(new_n249), .B1(new_n245), .B2(G134), .ZN(new_n262));
  AOI22_X1  g076(.A1(new_n252), .A2(new_n262), .B1(new_n243), .B2(new_n246), .ZN(new_n263));
  AOI22_X1  g077(.A1(G131), .A2(new_n256), .B1(new_n263), .B2(new_n258), .ZN(new_n264));
  NOR2_X1   g078(.A1(KEYINPUT78), .A2(KEYINPUT12), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  AOI211_X1 g080(.A(new_n264), .B(new_n266), .C1(new_n236), .C2(new_n240), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n261), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT77), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n264), .B(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n219), .ZN(new_n271));
  OAI21_X1  g085(.A(KEYINPUT1), .B1(new_n197), .B2(G146), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n208), .A2(G128), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n203), .A2(KEYINPUT67), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n215), .B1(new_n275), .B2(new_n214), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n205), .B1(new_n271), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT10), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n235), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(KEYINPUT0), .A2(G128), .ZN(new_n280));
  OR2_X1    g094(.A1(KEYINPUT0), .A2(G128), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n214), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n280), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n198), .A2(new_n201), .A3(new_n202), .A4(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n228), .A2(new_n230), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n227), .B1(new_n286), .B2(new_n226), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT4), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n285), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n226), .A2(new_n228), .A3(new_n230), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(G101), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n291), .A2(KEYINPUT4), .A3(new_n231), .ZN(new_n292));
  AOI22_X1  g106(.A1(new_n277), .A2(new_n279), .B1(new_n289), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT76), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n294), .B1(new_n240), .B2(new_n278), .ZN(new_n295));
  AND2_X1   g109(.A1(new_n231), .A2(new_n234), .ZN(new_n296));
  AOI211_X1 g110(.A(KEYINPUT76), .B(KEYINPUT10), .C1(new_n296), .C2(new_n239), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n270), .B(new_n293), .C1(new_n295), .C2(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n194), .B1(new_n268), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n298), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n293), .B1(new_n297), .B2(new_n295), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT79), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n264), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n293), .B(KEYINPUT79), .C1(new_n297), .C2(new_n295), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n300), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n299), .B1(new_n305), .B2(new_n194), .ZN(new_n306));
  OAI21_X1  g120(.A(G469), .B1(new_n306), .B2(G902), .ZN(new_n307));
  INV_X1    g121(.A(G469), .ZN(new_n308));
  INV_X1    g122(.A(G902), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n301), .A2(new_n302), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n310), .A2(new_n260), .A3(new_n304), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n194), .B1(new_n311), .B2(new_n298), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n241), .A2(new_n260), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(new_n195), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n241), .A2(new_n260), .A3(new_n265), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n298), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n316), .A2(new_n193), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n308), .B(new_n309), .C1(new_n312), .C2(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n189), .B1(new_n307), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G953), .ZN(new_n320));
  AND2_X1   g134(.A1(new_n320), .A2(G952), .ZN(new_n321));
  NAND2_X1  g135(.A1(G234), .A2(G237), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n323), .B(KEYINPUT92), .ZN(new_n324));
  AND3_X1   g138(.A1(new_n322), .A2(G902), .A3(G953), .ZN(new_n325));
  XNOR2_X1  g139(.A(KEYINPUT21), .B(G898), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AND2_X1   g141(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(G214), .B1(G237), .B2(G902), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n329), .B(KEYINPUT80), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(G110), .B(G122), .ZN(new_n332));
  XOR2_X1   g146(.A(new_n332), .B(KEYINPUT8), .Z(new_n333));
  XNOR2_X1  g147(.A(KEYINPUT81), .B(KEYINPUT5), .ZN(new_n334));
  INV_X1    g148(.A(G116), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n335), .A2(G119), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G113), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(KEYINPUT84), .ZN(new_n339));
  XNOR2_X1  g153(.A(G116), .B(G119), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT5), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT84), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n337), .A2(new_n342), .A3(G113), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n339), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  XOR2_X1   g158(.A(KEYINPUT2), .B(G113), .Z(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n340), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n344), .A2(new_n346), .A3(new_n296), .ZN(new_n347));
  INV_X1    g161(.A(new_n340), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n337), .B(G113), .C1(new_n348), .C2(new_n334), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n346), .ZN(new_n350));
  AOI22_X1  g164(.A1(new_n347), .A2(KEYINPUT85), .B1(new_n235), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT85), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n344), .A2(new_n352), .A3(new_n346), .A4(new_n296), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n333), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  OR2_X1    g168(.A1(new_n345), .A2(new_n340), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n346), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n290), .A2(new_n288), .A3(G101), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n231), .A2(KEYINPUT4), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n356), .B(new_n357), .C1(new_n358), .C2(new_n287), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n296), .A2(new_n346), .A3(new_n349), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(new_n360), .A3(new_n332), .ZN(new_n361));
  INV_X1    g175(.A(G125), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n220), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n285), .A2(G125), .ZN(new_n364));
  INV_X1    g178(.A(G224), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n365), .A2(G953), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(KEYINPUT7), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n363), .A2(new_n364), .A3(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n368), .B1(new_n363), .B2(new_n364), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n361), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n309), .B1(new_n354), .B2(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n364), .B1(new_n277), .B2(G125), .ZN(new_n374));
  XNOR2_X1  g188(.A(new_n374), .B(new_n367), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n359), .A2(new_n360), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n332), .B(KEYINPUT82), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT83), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT6), .ZN(new_n381));
  AND2_X1   g195(.A1(new_n359), .A2(new_n360), .ZN(new_n382));
  AOI22_X1  g196(.A1(new_n380), .A2(new_n381), .B1(new_n382), .B2(new_n332), .ZN(new_n383));
  INV_X1    g197(.A(new_n379), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n384), .B1(new_n359), .B2(new_n360), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(KEYINPUT6), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n375), .B1(new_n383), .B2(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(G210), .B1(G237), .B2(G902), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  NOR3_X1   g203(.A1(new_n373), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n347), .A2(KEYINPUT85), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n350), .A2(new_n235), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(new_n353), .A3(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n333), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n374), .A2(KEYINPUT7), .A3(new_n367), .ZN(new_n396));
  AOI22_X1  g210(.A1(new_n396), .A2(new_n369), .B1(new_n382), .B2(new_n332), .ZN(new_n397));
  AOI21_X1  g211(.A(G902), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n374), .B(new_n366), .ZN(new_n399));
  INV_X1    g213(.A(new_n386), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n361), .B1(new_n385), .B2(KEYINPUT6), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n399), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n388), .B1(new_n398), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n331), .B1(new_n390), .B2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT86), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n328), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  OAI211_X1 g220(.A(KEYINPUT86), .B(new_n331), .C1(new_n390), .C2(new_n403), .ZN(new_n407));
  XNOR2_X1  g221(.A(KEYINPUT71), .B(G217), .ZN(new_n408));
  NOR3_X1   g222(.A1(new_n408), .A2(new_n187), .A3(G953), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT90), .ZN(new_n410));
  INV_X1    g224(.A(G122), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n410), .B1(new_n411), .B2(G116), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n335), .A2(KEYINPUT90), .A3(G122), .ZN(new_n413));
  AOI22_X1  g227(.A1(new_n412), .A2(new_n413), .B1(G116), .B2(new_n411), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n411), .A2(G116), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n224), .B1(new_n415), .B2(KEYINPUT14), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n414), .B(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(G134), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n216), .A2(G143), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(KEYINPUT91), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT91), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n216), .A2(new_n421), .A3(G143), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n197), .A2(G128), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n418), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n424), .ZN(new_n426));
  AOI211_X1 g240(.A(G134), .B(new_n426), .C1(new_n420), .C2(new_n422), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n417), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n423), .A2(new_n418), .A3(new_n424), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n414), .B(new_n224), .ZN(new_n430));
  XOR2_X1   g244(.A(new_n424), .B(KEYINPUT13), .Z(new_n431));
  AOI21_X1  g245(.A(new_n431), .B1(new_n420), .B2(new_n422), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n429), .B(new_n430), .C1(new_n432), .C2(new_n418), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n409), .B1(new_n428), .B2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n428), .A2(new_n433), .A3(new_n409), .ZN(new_n436));
  AOI21_X1  g250(.A(G902), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(G478), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n438), .A2(KEYINPUT15), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n437), .B(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT20), .ZN(new_n442));
  XNOR2_X1  g256(.A(G113), .B(G122), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n443), .B(new_n222), .ZN(new_n444));
  INV_X1    g258(.A(G237), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n445), .A2(new_n320), .A3(G214), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n446), .B(new_n197), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n447), .A2(KEYINPUT18), .A3(G131), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n446), .A2(new_n197), .ZN(new_n449));
  NOR2_X1   g263(.A1(G237), .A2(G953), .ZN(new_n450));
  AOI21_X1  g264(.A(G143), .B1(new_n450), .B2(G214), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT18), .ZN(new_n453));
  INV_X1    g267(.A(G131), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  XNOR2_X1  g269(.A(G125), .B(G140), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n456), .B(new_n200), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n448), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT87), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n448), .A2(new_n455), .A3(KEYINPUT87), .A4(new_n457), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT88), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n447), .A2(new_n463), .A3(KEYINPUT17), .A4(G131), .ZN(new_n464));
  OAI211_X1 g278(.A(KEYINPUT17), .B(G131), .C1(new_n449), .C2(new_n451), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(KEYINPUT88), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(G140), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(G125), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n362), .A2(G140), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n469), .A2(new_n470), .A3(KEYINPUT16), .ZN(new_n471));
  OR3_X1    g285(.A1(new_n362), .A2(KEYINPUT16), .A3(G140), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n471), .A2(new_n472), .A3(G146), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(KEYINPUT73), .ZN(new_n474));
  AOI21_X1  g288(.A(G146), .B1(new_n471), .B2(new_n472), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n471), .A2(G146), .A3(new_n472), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT73), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n467), .A2(KEYINPUT89), .A3(new_n474), .A4(new_n478), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n452), .B(G131), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT17), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n474), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n473), .A2(KEYINPUT73), .ZN(new_n485));
  NOR3_X1   g299(.A1(new_n484), .A2(new_n475), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(KEYINPUT89), .B1(new_n486), .B2(new_n467), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n444), .B(new_n462), .C1(new_n483), .C2(new_n487), .ZN(new_n488));
  XOR2_X1   g302(.A(new_n456), .B(KEYINPUT19), .Z(new_n489));
  OAI21_X1  g303(.A(new_n473), .B1(new_n489), .B2(G146), .ZN(new_n490));
  OR2_X1    g304(.A1(new_n490), .A2(new_n480), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n462), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n444), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n488), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g309(.A1(G475), .A2(G902), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n442), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n496), .ZN(new_n498));
  AOI211_X1 g312(.A(KEYINPUT20), .B(new_n498), .C1(new_n488), .C2(new_n494), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n462), .B1(new_n483), .B2(new_n487), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(new_n493), .ZN(new_n501));
  AOI21_X1  g315(.A(G902), .B1(new_n501), .B2(new_n488), .ZN(new_n502));
  INV_X1    g316(.A(G475), .ZN(new_n503));
  OAI22_X1  g317(.A1(new_n497), .A2(new_n499), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n441), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n319), .A2(new_n406), .A3(new_n407), .A4(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT70), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n255), .A2(new_n251), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(G131), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n259), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n213), .A2(new_n219), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n510), .B1(new_n511), .B2(new_n205), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n285), .B1(new_n257), .B2(new_n259), .ZN(new_n513));
  NOR3_X1   g327(.A1(new_n512), .A2(new_n513), .A3(new_n356), .ZN(new_n514));
  INV_X1    g328(.A(new_n356), .ZN(new_n515));
  INV_X1    g329(.A(new_n510), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n277), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n285), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n454), .B1(new_n263), .B2(new_n255), .ZN(new_n519));
  INV_X1    g333(.A(new_n259), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n515), .B1(new_n517), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(KEYINPUT28), .B1(new_n514), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n450), .A2(G210), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n524), .B(KEYINPUT27), .ZN(new_n525));
  XNOR2_X1  g339(.A(KEYINPUT26), .B(G101), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n525), .B(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n517), .A2(new_n521), .A3(new_n515), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT28), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n523), .A2(KEYINPUT29), .A3(new_n527), .A4(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT29), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n527), .B1(new_n514), .B2(KEYINPUT28), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n356), .B1(new_n512), .B2(new_n513), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n529), .B1(new_n534), .B2(new_n528), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n532), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT30), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n537), .B1(new_n512), .B2(new_n513), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n517), .A2(KEYINPUT30), .A3(new_n521), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n538), .A2(new_n539), .A3(new_n356), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n527), .B1(new_n540), .B2(new_n528), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n531), .B(new_n309), .C1(new_n536), .C2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(G472), .ZN(new_n543));
  OAI21_X1  g357(.A(KEYINPUT30), .B1(new_n220), .B2(new_n510), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n356), .B1(new_n544), .B2(new_n513), .ZN(new_n545));
  AOI21_X1  g359(.A(KEYINPUT30), .B1(new_n517), .B2(new_n521), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n528), .A2(new_n527), .ZN(new_n548));
  OAI21_X1  g362(.A(KEYINPUT31), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n527), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n512), .A2(new_n513), .ZN(new_n551));
  AOI21_X1  g365(.A(KEYINPUT28), .B1(new_n551), .B2(new_n515), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n550), .B1(new_n535), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n550), .B1(new_n551), .B2(new_n515), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT31), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n540), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(KEYINPUT69), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT69), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n540), .A2(new_n555), .A3(new_n559), .A4(new_n556), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n554), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g375(.A1(G472), .A2(G902), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT32), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n543), .B1(new_n561), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n558), .A2(new_n560), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n523), .A2(new_n530), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n540), .A2(new_n555), .ZN(new_n570));
  AOI22_X1  g384(.A1(new_n569), .A2(new_n550), .B1(new_n570), .B2(KEYINPUT31), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(KEYINPUT32), .B1(new_n572), .B2(new_n562), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n507), .B1(new_n567), .B2(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n564), .B1(new_n561), .B2(new_n563), .ZN(new_n575));
  AOI22_X1  g389(.A1(new_n572), .A2(new_n565), .B1(G472), .B2(new_n542), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n575), .A2(new_n576), .A3(KEYINPUT70), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n408), .B1(G234), .B2(new_n309), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n478), .A2(new_n474), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n216), .A2(G119), .ZN(new_n581));
  INV_X1    g395(.A(G119), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(G128), .ZN(new_n583));
  XOR2_X1   g397(.A(KEYINPUT24), .B(G110), .Z(new_n584));
  NAND3_X1  g398(.A1(new_n581), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n216), .A2(KEYINPUT23), .A3(G119), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT23), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n587), .B1(new_n582), .B2(G128), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n586), .A2(new_n583), .A3(new_n588), .ZN(new_n589));
  AND3_X1   g403(.A1(new_n589), .A2(KEYINPUT72), .A3(G110), .ZN(new_n590));
  AOI21_X1  g404(.A(KEYINPUT72), .B1(new_n589), .B2(G110), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n580), .B(new_n585), .C1(new_n590), .C2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n456), .A2(new_n200), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n589), .A2(G110), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n584), .B1(new_n581), .B2(new_n583), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n473), .B(new_n593), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(KEYINPUT22), .B(G137), .ZN(new_n598));
  AND3_X1   g412(.A1(new_n320), .A2(G221), .A3(G234), .ZN(new_n599));
  XOR2_X1   g413(.A(new_n598), .B(new_n599), .Z(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n592), .A2(new_n596), .A3(new_n600), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n602), .A2(new_n309), .A3(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT25), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n602), .A2(KEYINPUT25), .A3(new_n309), .A4(new_n603), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n579), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n603), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n600), .B1(new_n592), .B2(new_n596), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n578), .A2(G902), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n608), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n574), .A2(new_n577), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(KEYINPUT74), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT74), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n574), .A2(new_n577), .A3(new_n616), .A4(new_n613), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n506), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(new_n227), .ZN(G3));
  INV_X1    g433(.A(new_n329), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n389), .B1(new_n373), .B2(new_n387), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n398), .A2(new_n388), .A3(new_n402), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n620), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  OR2_X1    g438(.A1(new_n624), .A2(new_n328), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n438), .A2(new_n309), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n626), .B1(new_n437), .B2(new_n438), .ZN(new_n627));
  INV_X1    g441(.A(new_n436), .ZN(new_n628));
  OAI21_X1  g442(.A(KEYINPUT33), .B1(new_n628), .B2(new_n434), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT33), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n435), .A2(new_n630), .A3(new_n436), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n629), .A2(new_n631), .A3(G478), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n627), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n495), .A2(new_n496), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(KEYINPUT20), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n495), .A2(new_n442), .A3(new_n496), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AND2_X1   g451(.A1(new_n501), .A2(new_n488), .ZN(new_n638));
  OAI21_X1  g452(.A(G475), .B1(new_n638), .B2(G902), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n633), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n625), .A2(new_n641), .ZN(new_n642));
  OAI21_X1  g456(.A(G472), .B1(new_n561), .B2(G902), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n572), .A2(new_n562), .ZN(new_n644));
  AND3_X1   g458(.A1(new_n643), .A2(new_n613), .A3(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n642), .A2(new_n319), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT34), .B(G104), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G6));
  NAND3_X1  g462(.A1(new_n635), .A2(KEYINPUT93), .A3(new_n636), .ZN(new_n649));
  OR2_X1    g463(.A1(new_n636), .A2(KEYINPUT93), .ZN(new_n650));
  AND3_X1   g464(.A1(new_n649), .A2(new_n639), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n441), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n652), .A2(new_n625), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n653), .A2(new_n319), .A3(new_n645), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT35), .B(G107), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G9));
  AND2_X1   g470(.A1(new_n643), .A2(new_n644), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n606), .A2(new_n607), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n578), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n597), .A2(KEYINPUT94), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT94), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n592), .A2(new_n661), .A3(new_n596), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n601), .A2(KEYINPUT36), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n660), .A2(new_n664), .A3(new_n662), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n612), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n659), .A2(KEYINPUT95), .A3(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT95), .ZN(new_n671));
  INV_X1    g485(.A(new_n612), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n672), .B1(new_n666), .B2(new_n667), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n671), .B1(new_n608), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n657), .A2(new_n675), .ZN(new_n676));
  OR2_X1    g490(.A1(new_n676), .A2(KEYINPUT96), .ZN(new_n677));
  INV_X1    g491(.A(new_n506), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n676), .A2(KEYINPUT96), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT37), .B(G110), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G12));
  NAND4_X1  g496(.A1(new_n574), .A2(new_n577), .A3(new_n319), .A4(new_n675), .ZN(new_n683));
  INV_X1    g497(.A(G900), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n325), .A2(new_n684), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n324), .A2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n651), .A2(new_n441), .A3(new_n623), .A4(new_n687), .ZN(new_n688));
  OR2_X1    g502(.A1(new_n683), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(KEYINPUT97), .B(G128), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G30));
  XOR2_X1   g505(.A(new_n686), .B(KEYINPUT39), .Z(new_n692));
  NAND2_X1  g506(.A1(new_n319), .A2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT40), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT100), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n693), .B(KEYINPUT40), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(KEYINPUT100), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n390), .A2(new_n403), .ZN(new_n700));
  XNOR2_X1  g514(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(new_n675), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n702), .A2(new_n329), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n441), .A2(new_n504), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n527), .B1(new_n534), .B2(new_n528), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n570), .B1(KEYINPUT99), .B2(new_n706), .ZN(new_n707));
  AND2_X1   g521(.A1(new_n706), .A2(KEYINPUT99), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n309), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  AOI22_X1  g523(.A1(new_n572), .A2(new_n565), .B1(new_n709), .B2(G472), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n575), .A2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NOR3_X1   g526(.A1(new_n704), .A2(new_n705), .A3(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n697), .A2(new_n699), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(KEYINPUT101), .B(G143), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G45));
  AND2_X1   g530(.A1(new_n627), .A2(new_n632), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n623), .A2(new_n504), .A3(new_n717), .A4(new_n687), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT102), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n640), .A2(KEYINPUT102), .A3(new_n623), .A4(new_n687), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n683), .A2(new_n722), .ZN(new_n723));
  XOR2_X1   g537(.A(KEYINPUT103), .B(G146), .Z(new_n724));
  XNOR2_X1  g538(.A(new_n723), .B(new_n724), .ZN(G48));
  NAND2_X1  g539(.A1(new_n311), .A2(new_n298), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n317), .B1(new_n726), .B2(new_n193), .ZN(new_n727));
  OAI21_X1  g541(.A(G469), .B1(new_n727), .B2(G902), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n728), .A2(new_n188), .A3(new_n318), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(KEYINPUT104), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT104), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n728), .A2(new_n731), .A3(new_n188), .A4(new_n318), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n574), .A2(new_n577), .A3(new_n613), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n733), .A2(new_n734), .A3(new_n642), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(KEYINPUT105), .ZN(new_n736));
  XOR2_X1   g550(.A(KEYINPUT41), .B(G113), .Z(new_n737));
  XNOR2_X1  g551(.A(new_n736), .B(new_n737), .ZN(G15));
  NAND3_X1  g552(.A1(new_n733), .A2(new_n734), .A3(new_n653), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G116), .ZN(G18));
  NAND3_X1  g554(.A1(new_n574), .A2(new_n577), .A3(new_n675), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n728), .A2(new_n188), .A3(new_n318), .A4(new_n623), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n441), .A2(new_n504), .A3(new_n328), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n742), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G119), .ZN(G21));
  NAND2_X1  g561(.A1(new_n644), .A2(KEYINPUT106), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT106), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n572), .A2(new_n749), .A3(new_n562), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n751), .A2(new_n613), .A3(new_n643), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n625), .A2(new_n705), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n753), .A2(new_n754), .A3(new_n730), .A4(new_n732), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G122), .ZN(G24));
  AND3_X1   g570(.A1(new_n504), .A2(new_n717), .A3(new_n687), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n751), .A2(new_n675), .A3(new_n757), .A4(new_n643), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n758), .A2(new_n743), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(new_n362), .ZN(G27));
  NAND2_X1  g574(.A1(new_n316), .A2(new_n193), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT108), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n311), .A2(new_n194), .A3(new_n298), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n316), .A2(KEYINPUT108), .A3(new_n193), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n763), .A2(G469), .A3(new_n764), .A4(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT109), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  AOI211_X1 g582(.A(new_n762), .B(new_n194), .C1(new_n268), .C2(new_n298), .ZN(new_n769));
  AOI21_X1  g583(.A(KEYINPUT108), .B1(new_n316), .B2(new_n193), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n771), .A2(KEYINPUT109), .A3(G469), .A4(new_n764), .ZN(new_n772));
  NAND2_X1  g586(.A1(G469), .A2(G902), .ZN(new_n773));
  XOR2_X1   g587(.A(new_n773), .B(KEYINPUT107), .Z(new_n774));
  NAND4_X1  g588(.A1(new_n768), .A2(new_n772), .A3(new_n318), .A4(new_n774), .ZN(new_n775));
  NOR3_X1   g589(.A1(new_n390), .A2(new_n403), .A3(new_n620), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n776), .A2(new_n188), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n775), .A2(new_n777), .A3(KEYINPUT110), .ZN(new_n778));
  AOI21_X1  g592(.A(KEYINPUT110), .B1(new_n775), .B2(new_n777), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n734), .B(new_n757), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(KEYINPUT111), .B(KEYINPUT42), .ZN(new_n781));
  INV_X1    g595(.A(new_n779), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n775), .A2(new_n777), .A3(KEYINPUT110), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n575), .A2(new_n576), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n613), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  AND3_X1   g601(.A1(new_n787), .A2(KEYINPUT42), .A3(new_n757), .ZN(new_n788));
  AOI22_X1  g602(.A1(new_n780), .A2(new_n781), .B1(new_n784), .B2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(new_n454), .ZN(G33));
  NOR2_X1   g604(.A1(new_n652), .A2(new_n686), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n734), .B(new_n791), .C1(new_n778), .C2(new_n779), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G134), .ZN(G36));
  NAND3_X1  g607(.A1(new_n771), .A2(KEYINPUT45), .A3(new_n764), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n764), .A2(new_n761), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT45), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n308), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n798), .A2(KEYINPUT46), .A3(new_n774), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n799), .A2(KEYINPUT112), .A3(new_n318), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT46), .ZN(new_n801));
  INV_X1    g615(.A(new_n798), .ZN(new_n802));
  INV_X1    g616(.A(new_n774), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n801), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n800), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(KEYINPUT112), .B1(new_n799), .B2(new_n318), .ZN(new_n806));
  OR2_X1    g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n807), .A2(new_n188), .A3(new_n692), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT113), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n807), .A2(KEYINPUT113), .A3(new_n188), .A4(new_n692), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n717), .A2(new_n637), .A3(new_n639), .ZN(new_n812));
  OR2_X1    g626(.A1(new_n812), .A2(KEYINPUT43), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(KEYINPUT43), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n815), .A2(new_n657), .A3(new_n703), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n776), .B1(new_n816), .B2(KEYINPUT44), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n817), .B1(KEYINPUT44), .B2(new_n816), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n810), .A2(new_n811), .A3(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(G137), .ZN(G39));
  INV_X1    g634(.A(new_n776), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n821), .A2(new_n613), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(new_n757), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n823), .B1(new_n574), .B2(new_n577), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n807), .A2(KEYINPUT47), .A3(new_n188), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(KEYINPUT47), .B1(new_n807), .B2(new_n188), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n824), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(G140), .ZN(G42));
  NAND3_X1  g643(.A1(new_n613), .A2(new_n331), .A3(new_n188), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n830), .A2(new_n812), .ZN(new_n831));
  XOR2_X1   g645(.A(new_n831), .B(KEYINPUT114), .Z(new_n832));
  NAND2_X1  g646(.A1(new_n728), .A2(new_n318), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(KEYINPUT49), .ZN(new_n834));
  OR2_X1    g648(.A1(new_n833), .A2(KEYINPUT49), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n702), .A2(new_n711), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n832), .A2(new_n834), .A3(new_n835), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n645), .A2(new_n319), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n406), .A2(new_n407), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n504), .A2(new_n440), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n680), .A2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n615), .A2(new_n617), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(new_n678), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n838), .A2(new_n839), .A3(new_n641), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(KEYINPUT115), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT115), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n618), .A2(new_n850), .A3(new_n847), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n844), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  AND4_X1   g666(.A1(new_n735), .A2(new_n739), .A3(new_n746), .A4(new_n755), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n780), .A2(new_n781), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n784), .A2(new_n788), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n821), .A2(new_n441), .A3(new_n686), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n742), .A2(new_n319), .A3(new_n651), .A4(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n758), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n859), .B1(new_n778), .B2(new_n779), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n792), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n853), .A2(new_n856), .A3(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n852), .A2(new_n862), .ZN(new_n863));
  OAI22_X1  g677(.A1(new_n683), .A2(new_n688), .B1(new_n758), .B2(new_n743), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n659), .A2(new_n669), .A3(new_n188), .A4(new_n687), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n865), .B1(new_n575), .B2(new_n710), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n705), .A2(new_n624), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n866), .A2(new_n775), .A3(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n864), .A2(new_n723), .A3(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(KEYINPUT116), .B1(new_n870), .B2(KEYINPUT52), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(KEYINPUT52), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n870), .A2(KEYINPUT116), .A3(KEYINPUT52), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(KEYINPUT53), .B1(new_n863), .B2(new_n875), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n735), .A2(new_n739), .A3(new_n746), .A4(new_n755), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n792), .A2(new_n858), .A3(new_n860), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n789), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n846), .A2(new_n848), .A3(KEYINPUT115), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n850), .B1(new_n618), .B2(new_n847), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n843), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(new_n723), .ZN(new_n883));
  INV_X1    g697(.A(new_n759), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n883), .A2(new_n689), .A3(new_n884), .A4(new_n868), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT52), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(new_n872), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n879), .A2(new_n882), .A3(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT53), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(KEYINPUT54), .B1(new_n876), .B2(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n863), .A2(new_n875), .A3(KEYINPUT53), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT54), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n889), .A2(new_n890), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n892), .A2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT51), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n815), .A2(new_n324), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n729), .A2(new_n821), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n751), .A2(new_n643), .A3(new_n675), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT119), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n815), .A2(new_n752), .A3(new_n324), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n702), .A2(new_n329), .A3(new_n729), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n907), .B(KEYINPUT50), .Z(new_n908));
  INV_X1    g722(.A(new_n324), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n900), .A2(new_n613), .A3(new_n909), .A4(new_n712), .ZN(new_n910));
  OR3_X1    g724(.A1(new_n910), .A2(new_n504), .A3(new_n717), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n904), .A2(new_n908), .A3(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n827), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n728), .A2(new_n189), .A3(new_n318), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n913), .A2(new_n825), .A3(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT120), .ZN(new_n916));
  OR2_X1    g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n905), .A2(new_n776), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(KEYINPUT117), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n920), .B1(new_n915), .B2(new_n916), .ZN(new_n921));
  AOI211_X1 g735(.A(new_n898), .B(new_n912), .C1(new_n917), .C2(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n321), .B1(new_n910), .B2(new_n641), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n901), .A2(new_n786), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT48), .ZN(new_n925));
  AOI211_X1 g739(.A(new_n923), .B(new_n925), .C1(new_n744), .C2(new_n905), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n914), .B(KEYINPUT118), .Z(new_n927));
  NAND3_X1  g741(.A1(new_n913), .A2(new_n825), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n912), .B1(new_n919), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n926), .B1(new_n929), .B2(KEYINPUT51), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n897), .A2(new_n922), .A3(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(G952), .A2(G953), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n837), .B1(new_n931), .B2(new_n932), .ZN(G75));
  INV_X1    g747(.A(KEYINPUT56), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n893), .A2(new_n895), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(G902), .ZN(new_n936));
  INV_X1    g750(.A(G210), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n934), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n383), .A2(new_n375), .A3(new_n386), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(new_n402), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT55), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n941), .ZN(new_n943));
  OAI211_X1 g757(.A(new_n934), .B(new_n943), .C1(new_n936), .C2(new_n937), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n320), .A2(G952), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  AND3_X1   g760(.A1(new_n942), .A2(new_n944), .A3(new_n946), .ZN(G51));
  INV_X1    g761(.A(new_n896), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n894), .B1(new_n893), .B2(new_n895), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n774), .B(KEYINPUT57), .ZN(new_n951));
  OAI22_X1  g765(.A1(new_n950), .A2(new_n951), .B1(new_n312), .B2(new_n317), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n935), .A2(G902), .A3(new_n802), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n945), .B1(new_n952), .B2(new_n953), .ZN(G54));
  INV_X1    g768(.A(KEYINPUT121), .ZN(new_n955));
  NAND2_X1  g769(.A1(KEYINPUT58), .A2(G475), .ZN(new_n956));
  AOI211_X1 g770(.A(new_n309), .B(new_n956), .C1(new_n893), .C2(new_n895), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n946), .B1(new_n957), .B2(new_n495), .ZN(new_n958));
  INV_X1    g772(.A(new_n956), .ZN(new_n959));
  AND4_X1   g773(.A1(G902), .A2(new_n935), .A3(new_n495), .A4(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n955), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n495), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n962), .B1(new_n936), .B2(new_n956), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n957), .A2(new_n495), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n963), .A2(new_n964), .A3(KEYINPUT121), .A4(new_n946), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n961), .A2(new_n965), .ZN(G60));
  AND2_X1   g780(.A1(new_n629), .A2(new_n631), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n626), .B(KEYINPUT59), .Z(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n946), .B1(new_n950), .B2(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n968), .B1(new_n897), .B2(new_n969), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n971), .A2(new_n972), .ZN(G63));
  NAND2_X1  g787(.A1(G217), .A2(G902), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT60), .ZN(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n935), .A2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n611), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n945), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n975), .B1(new_n893), .B2(new_n895), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(new_n668), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT122), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n979), .B(new_n981), .C1(new_n982), .C2(KEYINPUT61), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT61), .ZN(new_n984));
  OAI211_X1 g798(.A(new_n982), .B(new_n946), .C1(new_n980), .C2(new_n611), .ZN(new_n985));
  INV_X1    g799(.A(new_n981), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n946), .B1(new_n980), .B2(new_n611), .ZN(new_n987));
  OAI211_X1 g801(.A(new_n984), .B(new_n985), .C1(new_n986), .C2(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n983), .A2(new_n988), .ZN(G66));
  OAI21_X1  g803(.A(G953), .B1(new_n326), .B2(new_n365), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n882), .A2(new_n853), .ZN(new_n991));
  AND3_X1   g805(.A1(new_n991), .A2(KEYINPUT123), .A3(new_n320), .ZN(new_n992));
  AOI21_X1  g806(.A(KEYINPUT123), .B1(new_n991), .B2(new_n320), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n990), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(KEYINPUT124), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT124), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n996), .B(new_n990), .C1(new_n992), .C2(new_n993), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n320), .A2(G898), .ZN(new_n999));
  NOR3_X1   g813(.A1(new_n400), .A2(new_n401), .A3(new_n999), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n998), .B(new_n1000), .ZN(G69));
  INV_X1    g815(.A(KEYINPUT62), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n864), .A2(new_n723), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n714), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT126), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1004), .B(new_n1005), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n1002), .B1(new_n714), .B2(new_n1003), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n776), .B1(new_n841), .B2(new_n640), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n693), .A2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1007), .B1(new_n845), .B2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n1006), .A2(new_n819), .A3(new_n828), .A4(new_n1010), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1011), .A2(new_n320), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n538), .A2(new_n539), .ZN(new_n1013));
  XOR2_X1   g827(.A(new_n1013), .B(KEYINPUT125), .Z(new_n1014));
  XOR2_X1   g828(.A(new_n1014), .B(new_n489), .Z(new_n1015));
  INV_X1    g829(.A(new_n1015), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1012), .A2(new_n1016), .ZN(new_n1017));
  NAND4_X1  g831(.A1(new_n810), .A2(new_n787), .A3(new_n811), .A4(new_n867), .ZN(new_n1018));
  AND3_X1   g832(.A1(new_n856), .A2(new_n792), .A3(new_n1003), .ZN(new_n1019));
  NAND4_X1  g833(.A1(new_n1018), .A2(new_n819), .A3(new_n828), .A4(new_n1019), .ZN(new_n1020));
  NOR2_X1   g834(.A1(new_n1020), .A2(G953), .ZN(new_n1021));
  NAND2_X1  g835(.A1(G900), .A2(G953), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1015), .A2(new_n1022), .ZN(new_n1023));
  OR2_X1    g837(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g838(.A(G953), .B1(new_n191), .B2(new_n684), .ZN(new_n1025));
  OR2_X1    g839(.A1(new_n1025), .A2(KEYINPUT127), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1025), .A2(KEYINPUT127), .ZN(new_n1027));
  NAND4_X1  g841(.A1(new_n1017), .A2(new_n1024), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1015), .B1(new_n1011), .B2(new_n320), .ZN(new_n1029));
  NOR2_X1   g843(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1030));
  OAI211_X1 g844(.A(KEYINPUT127), .B(new_n1025), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1031));
  AND2_X1   g845(.A1(new_n1028), .A2(new_n1031), .ZN(G72));
  NAND2_X1  g846(.A1(G472), .A2(G902), .ZN(new_n1033));
  XOR2_X1   g847(.A(new_n1033), .B(KEYINPUT63), .Z(new_n1034));
  OAI21_X1  g848(.A(new_n1034), .B1(new_n1011), .B2(new_n991), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n540), .A2(new_n528), .ZN(new_n1036));
  NAND3_X1  g850(.A1(new_n1035), .A2(new_n527), .A3(new_n1036), .ZN(new_n1037));
  NAND3_X1  g851(.A1(new_n540), .A2(new_n528), .A3(new_n550), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1036), .A2(new_n527), .ZN(new_n1039));
  AND2_X1   g853(.A1(new_n1039), .A2(new_n1034), .ZN(new_n1040));
  OAI211_X1 g854(.A(new_n1038), .B(new_n1040), .C1(new_n876), .C2(new_n891), .ZN(new_n1041));
  OAI21_X1  g855(.A(new_n1034), .B1(new_n1020), .B2(new_n991), .ZN(new_n1042));
  INV_X1    g856(.A(new_n1038), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  AND4_X1   g858(.A1(new_n946), .A2(new_n1037), .A3(new_n1041), .A4(new_n1044), .ZN(G57));
endmodule


