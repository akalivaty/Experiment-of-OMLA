//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 0 0 1 0 0 1 0 0 1 1 0 0 0 1 0 0 1 0 1 1 0 0 1 1 1 0 0 0 0 1 1 0 1 0 1 0 0 0 0 0 0 0 0 0 1 0 1 1 1 0 0 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n743, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n833, new_n834,
    new_n836, new_n837, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n949, new_n950, new_n951, new_n952;
  INV_X1    g000(.A(KEYINPUT82), .ZN(new_n202));
  XOR2_X1   g001(.A(G155gat), .B(G162gat), .Z(new_n203));
  INV_X1    g002(.A(KEYINPUT2), .ZN(new_n204));
  AND2_X1   g003(.A1(KEYINPUT76), .A2(G162gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(KEYINPUT76), .A2(G162gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n204), .B1(new_n207), .B2(G155gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT77), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n203), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G141gat), .B(G148gat), .ZN(new_n211));
  XNOR2_X1  g010(.A(KEYINPUT76), .B(G162gat), .ZN(new_n212));
  INV_X1    g011(.A(G155gat), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT2), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n211), .B1(new_n214), .B2(KEYINPUT77), .ZN(new_n215));
  INV_X1    g014(.A(G148gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G141gat), .ZN(new_n217));
  INV_X1    g016(.A(G141gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(G148gat), .ZN(new_n219));
  AOI21_X1  g018(.A(KEYINPUT2), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(G155gat), .B(G162gat), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT75), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT75), .ZN(new_n223));
  OAI211_X1 g022(.A(new_n203), .B(new_n223), .C1(KEYINPUT2), .C2(new_n211), .ZN(new_n224));
  AOI22_X1  g023(.A1(new_n210), .A2(new_n215), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT3), .ZN(new_n226));
  AOI21_X1  g025(.A(KEYINPUT29), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(G218gat), .ZN(new_n228));
  OR2_X1    g027(.A1(G197gat), .A2(G204gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(G197gat), .A2(G204gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT71), .ZN(new_n231));
  INV_X1    g030(.A(G211gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(KEYINPUT71), .A2(G211gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n233), .A2(G218gat), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT22), .ZN(new_n236));
  AOI221_X4 g035(.A(G211gat), .B1(new_n229), .B2(new_n230), .C1(new_n235), .C2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(new_n236), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n229), .A2(new_n230), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n232), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n228), .B1(new_n237), .B2(new_n240), .ZN(new_n241));
  AND2_X1   g040(.A1(KEYINPUT71), .A2(G211gat), .ZN(new_n242));
  NOR2_X1   g041(.A1(KEYINPUT71), .A2(G211gat), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(KEYINPUT22), .B1(new_n244), .B2(G218gat), .ZN(new_n245));
  INV_X1    g044(.A(new_n239), .ZN(new_n246));
  OAI21_X1  g045(.A(G211gat), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n238), .A2(new_n232), .A3(new_n239), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n247), .A2(G218gat), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n241), .A2(new_n249), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n202), .B1(new_n227), .B2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n250), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n224), .A2(new_n222), .ZN(new_n253));
  INV_X1    g052(.A(new_n211), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n254), .B1(new_n208), .B2(new_n209), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n221), .B1(new_n214), .B2(KEYINPUT77), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n226), .B(new_n253), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT29), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n252), .A2(new_n259), .A3(KEYINPUT82), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n251), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(G228gat), .ZN(new_n262));
  INV_X1    g061(.A(G233gat), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NOR3_X1   g063(.A1(new_n237), .A2(new_n240), .A3(new_n228), .ZN(new_n265));
  AOI21_X1  g064(.A(G218gat), .B1(new_n247), .B2(new_n248), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n258), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(new_n226), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n253), .B1(new_n255), .B2(new_n256), .ZN(new_n269));
  AOI21_X1  g068(.A(KEYINPUT81), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(KEYINPUT29), .B1(new_n241), .B2(new_n249), .ZN(new_n271));
  OAI211_X1 g070(.A(KEYINPUT81), .B(new_n269), .C1(new_n271), .C2(KEYINPUT3), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  OAI211_X1 g072(.A(new_n261), .B(new_n264), .C1(new_n270), .C2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT83), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT81), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n271), .A2(KEYINPUT3), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n277), .B1(new_n278), .B2(new_n225), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(new_n272), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n280), .A2(KEYINPUT83), .A3(new_n261), .A4(new_n264), .ZN(new_n281));
  INV_X1    g080(.A(new_n264), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n225), .B1(new_n267), .B2(new_n226), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n227), .A2(new_n250), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT80), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI211_X1 g086(.A(KEYINPUT80), .B(new_n282), .C1(new_n283), .C2(new_n284), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n276), .A2(new_n281), .A3(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(G78gat), .B(G106gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(KEYINPUT31), .B(G50gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n291), .B(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n293), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n276), .A2(new_n289), .A3(new_n281), .A4(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(KEYINPUT84), .B(G22gat), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n294), .A2(new_n298), .A3(new_n296), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT25), .ZN(new_n302));
  NOR2_X1   g101(.A1(G169gat), .A2(G176gat), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT23), .ZN(new_n304));
  XNOR2_X1  g103(.A(new_n303), .B(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(G169gat), .A2(G176gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  OR2_X1    g106(.A1(G183gat), .A2(G190gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(G183gat), .A2(G190gat), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n308), .A2(KEYINPUT24), .A3(new_n309), .ZN(new_n310));
  OR2_X1    g109(.A1(new_n309), .A2(KEYINPUT24), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n302), .B1(new_n307), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n312), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n306), .A2(KEYINPUT65), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n315), .A2(new_n302), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n306), .A2(KEYINPUT65), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n314), .A2(new_n305), .A3(new_n316), .A4(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n313), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(G190gat), .ZN(new_n320));
  AND2_X1   g119(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n321));
  NOR2_X1   g120(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT28), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(KEYINPUT27), .B(G183gat), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n326), .A2(KEYINPUT28), .A3(new_n320), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G169gat), .ZN(new_n329));
  INV_X1    g128(.A(G176gat), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n329), .A2(new_n330), .A3(KEYINPUT66), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(KEYINPUT26), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT26), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n303), .A2(KEYINPUT66), .A3(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n332), .A2(new_n306), .A3(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n328), .A2(new_n309), .A3(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT67), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  AND2_X1   g137(.A1(new_n335), .A2(new_n309), .ZN(new_n339));
  AOI21_X1  g138(.A(KEYINPUT67), .B1(new_n339), .B2(new_n328), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n319), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(G113gat), .B(G120gat), .ZN(new_n342));
  OAI21_X1  g141(.A(G127gat), .B1(new_n342), .B2(KEYINPUT1), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT1), .ZN(new_n344));
  INV_X1    g143(.A(G127gat), .ZN(new_n345));
  INV_X1    g144(.A(G113gat), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n346), .A2(G120gat), .ZN(new_n347));
  INV_X1    g146(.A(G120gat), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n348), .A2(G113gat), .ZN(new_n349));
  OAI211_X1 g148(.A(new_n344), .B(new_n345), .C1(new_n347), .C2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n343), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(G134gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n343), .A2(new_n350), .A3(G134gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n341), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n336), .A2(new_n337), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n339), .A2(KEYINPUT67), .A3(new_n328), .ZN(new_n358));
  AOI22_X1  g157(.A1(new_n357), .A2(new_n358), .B1(new_n313), .B2(new_n318), .ZN(new_n359));
  AND3_X1   g158(.A1(new_n343), .A2(new_n350), .A3(G134gat), .ZN(new_n360));
  AOI21_X1  g159(.A(G134gat), .B1(new_n343), .B2(new_n350), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(G227gat), .A2(G233gat), .ZN(new_n364));
  XOR2_X1   g163(.A(new_n364), .B(KEYINPUT64), .Z(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n356), .A2(new_n363), .A3(new_n366), .ZN(new_n367));
  XOR2_X1   g166(.A(new_n367), .B(KEYINPUT34), .Z(new_n368));
  NAND2_X1  g167(.A1(new_n356), .A2(new_n363), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(new_n365), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT32), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT33), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(G15gat), .B(G43gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(KEYINPUT68), .B(KEYINPUT69), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n374), .B(new_n375), .ZN(new_n376));
  XOR2_X1   g175(.A(G71gat), .B(G99gat), .Z(new_n377));
  XOR2_X1   g176(.A(new_n376), .B(new_n377), .Z(new_n378));
  NAND3_X1  g177(.A1(new_n371), .A2(new_n373), .A3(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n378), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n370), .B(KEYINPUT32), .C1(new_n372), .C2(new_n380), .ZN(new_n381));
  AND3_X1   g180(.A1(new_n368), .A2(new_n379), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n368), .B1(new_n379), .B2(new_n381), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n300), .A2(new_n301), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(KEYINPUT92), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT74), .ZN(new_n387));
  NAND2_X1  g186(.A1(G226gat), .A2(G233gat), .ZN(new_n388));
  XOR2_X1   g187(.A(new_n388), .B(KEYINPUT72), .Z(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n359), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n319), .A2(new_n336), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n389), .B1(new_n392), .B2(new_n258), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n250), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  AOI22_X1  g193(.A1(new_n313), .A2(new_n318), .B1(new_n339), .B2(new_n328), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(new_n389), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n359), .A2(KEYINPUT29), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n397), .B1(new_n398), .B2(new_n390), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n394), .B1(new_n399), .B2(new_n250), .ZN(new_n400));
  XOR2_X1   g199(.A(G8gat), .B(G36gat), .Z(new_n401));
  XNOR2_X1  g200(.A(new_n401), .B(G64gat), .ZN(new_n402));
  INV_X1    g201(.A(G92gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n402), .B(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n387), .B1(new_n400), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT30), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n400), .A2(new_n387), .A3(new_n405), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n407), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(KEYINPUT4), .B1(new_n269), .B2(new_n355), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT4), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n225), .A2(new_n412), .A3(new_n362), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n225), .A2(new_n362), .ZN(new_n415));
  NAND2_X1  g214(.A1(G225gat), .A2(G233gat), .ZN(new_n416));
  XOR2_X1   g215(.A(new_n416), .B(KEYINPUT78), .Z(new_n417));
  NAND2_X1  g216(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n269), .A2(KEYINPUT3), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n419), .A2(new_n355), .A3(new_n257), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n414), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT5), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n269), .A2(new_n355), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n415), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n422), .B1(new_n424), .B2(new_n417), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n421), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n417), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n414), .A2(new_n420), .A3(new_n422), .A4(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  XOR2_X1   g228(.A(G1gat), .B(G29gat), .Z(new_n430));
  XNOR2_X1  g229(.A(G57gat), .B(G85gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n430), .B(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n432), .B(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n429), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT6), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n426), .A2(new_n428), .A3(new_n434), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n434), .B1(new_n426), .B2(new_n428), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(KEYINPUT6), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT73), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n400), .A2(KEYINPUT30), .A3(new_n405), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n341), .A2(new_n258), .A3(new_n390), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n250), .B1(new_n445), .B2(new_n396), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n447), .A2(new_n394), .A3(new_n404), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n444), .A2(new_n448), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n410), .B(new_n442), .C1(new_n443), .C2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n449), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n451), .A2(KEYINPUT73), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT92), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n300), .A2(new_n454), .A3(new_n301), .A4(new_n384), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n386), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT35), .ZN(new_n457));
  AOI21_X1  g256(.A(KEYINPUT89), .B1(new_n440), .B2(KEYINPUT6), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n458), .B1(new_n442), .B2(KEYINPUT89), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n410), .A2(new_n451), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT91), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  AOI211_X1 g260(.A(KEYINPUT74), .B(new_n404), .C1(new_n447), .C2(new_n394), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n462), .A2(new_n406), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n449), .B1(new_n463), .B2(new_n408), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT91), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT89), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n466), .B1(new_n439), .B2(new_n441), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n464), .B(new_n465), .C1(new_n467), .C2(new_n458), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n461), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT35), .ZN(new_n470));
  AND2_X1   g269(.A1(new_n300), .A2(new_n301), .ZN(new_n471));
  NOR3_X1   g270(.A1(new_n382), .A2(new_n383), .A3(KEYINPUT70), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n382), .A2(KEYINPUT70), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n469), .A2(new_n470), .A3(new_n471), .A4(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT90), .ZN(new_n477));
  AND3_X1   g276(.A1(new_n426), .A2(new_n434), .A3(new_n428), .ZN(new_n478));
  NOR3_X1   g277(.A1(new_n478), .A2(new_n440), .A3(KEYINPUT6), .ZN(new_n479));
  INV_X1    g278(.A(new_n441), .ZN(new_n480));
  OAI21_X1  g279(.A(KEYINPUT89), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n458), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT37), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n341), .A2(new_n389), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n390), .B1(new_n395), .B2(KEYINPUT29), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n252), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n483), .B1(new_n446), .B2(new_n486), .ZN(new_n487));
  XOR2_X1   g286(.A(KEYINPUT87), .B(KEYINPUT38), .Z(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n445), .A2(new_n250), .A3(new_n396), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n484), .A2(new_n252), .A3(new_n485), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n490), .A2(KEYINPUT37), .A3(new_n491), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n487), .A2(new_n404), .A3(new_n489), .A4(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT88), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n481), .A2(new_n463), .A3(new_n482), .A4(new_n495), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n493), .A2(new_n494), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n477), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AND2_X1   g297(.A1(new_n493), .A2(new_n494), .ZN(new_n499));
  NOR3_X1   g298(.A1(new_n467), .A2(new_n458), .A3(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n497), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n500), .A2(KEYINPUT90), .A3(new_n463), .A4(new_n501), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n400), .A2(new_n483), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n404), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n488), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n498), .A2(new_n502), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n414), .A2(new_n420), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(new_n417), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n508), .A2(KEYINPUT39), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n509), .A2(new_n435), .ZN(new_n510));
  OAI211_X1 g309(.A(new_n508), .B(KEYINPUT39), .C1(new_n417), .C2(new_n424), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT40), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  XOR2_X1   g313(.A(new_n514), .B(KEYINPUT86), .Z(new_n515));
  OR2_X1    g314(.A1(new_n512), .A2(KEYINPUT85), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n512), .A2(KEYINPUT85), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(new_n513), .A3(new_n517), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n515), .A2(new_n518), .A3(new_n436), .A4(new_n460), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n506), .A2(new_n471), .A3(new_n519), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n471), .A2(new_n453), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT36), .ZN(new_n522));
  INV_X1    g321(.A(new_n474), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n522), .B1(new_n472), .B2(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(KEYINPUT36), .B1(new_n382), .B2(new_n383), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n521), .A2(new_n526), .ZN(new_n527));
  AOI22_X1  g326(.A1(new_n457), .A2(new_n476), .B1(new_n520), .B2(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(G15gat), .B(G22gat), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT16), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n529), .B1(new_n530), .B2(G1gat), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n531), .B1(G1gat), .B2(new_n529), .ZN(new_n532));
  OR2_X1    g331(.A1(new_n532), .A2(G8gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(G8gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  XOR2_X1   g334(.A(G71gat), .B(G78gat), .Z(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT9), .ZN(new_n538));
  INV_X1    g337(.A(G71gat), .ZN(new_n539));
  INV_X1    g338(.A(G78gat), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  XOR2_X1   g340(.A(G57gat), .B(G64gat), .Z(new_n542));
  NAND3_X1  g341(.A1(new_n537), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n541), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(new_n536), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n535), .B1(KEYINPUT21), .B2(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(G183gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(G231gat), .A2(G233gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(G127gat), .B(G155gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(new_n232), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n551), .B(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n547), .A2(KEYINPUT21), .ZN(new_n555));
  XNOR2_X1  g354(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n555), .B(new_n556), .ZN(new_n557));
  OR2_X1    g356(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n554), .A2(new_n557), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(G43gat), .B(G50gat), .ZN(new_n561));
  OR2_X1    g360(.A1(new_n561), .A2(KEYINPUT15), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(KEYINPUT15), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT14), .ZN(new_n564));
  INV_X1    g363(.A(G29gat), .ZN(new_n565));
  INV_X1    g364(.A(G36gat), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(G29gat), .A2(G36gat), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n562), .A2(new_n563), .A3(new_n569), .A4(new_n570), .ZN(new_n571));
  AND3_X1   g370(.A1(new_n567), .A2(KEYINPUT93), .A3(new_n568), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n570), .B1(new_n567), .B2(KEYINPUT93), .ZN(new_n573));
  OAI211_X1 g372(.A(KEYINPUT15), .B(new_n561), .C1(new_n572), .C2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(KEYINPUT17), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT96), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n577), .A2(G85gat), .A3(G92gat), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT7), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(G99gat), .A2(G106gat), .ZN(new_n581));
  INV_X1    g380(.A(G85gat), .ZN(new_n582));
  AOI22_X1  g381(.A1(KEYINPUT8), .A2(new_n581), .B1(new_n582), .B2(new_n403), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n577), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n580), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(G99gat), .ZN(new_n586));
  INV_X1    g385(.A(G106gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n585), .A2(new_n581), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n581), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n580), .A2(new_n583), .A3(new_n590), .A4(new_n584), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n592), .ZN(new_n593));
  AND2_X1   g392(.A1(new_n589), .A2(new_n591), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(new_n575), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT41), .ZN(new_n596));
  NAND2_X1  g395(.A1(G232gat), .A2(G233gat), .ZN(new_n597));
  XOR2_X1   g396(.A(new_n597), .B(KEYINPUT95), .Z(new_n598));
  OAI211_X1 g397(.A(new_n593), .B(new_n595), .C1(new_n596), .C2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G134gat), .B(G162gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n598), .A2(new_n596), .ZN(new_n602));
  XOR2_X1   g401(.A(G190gat), .B(G218gat), .Z(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n601), .B(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n560), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n535), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n576), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n535), .A2(new_n575), .ZN(new_n609));
  NAND2_X1  g408(.A1(G229gat), .A2(G233gat), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT18), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n611), .A2(KEYINPUT94), .A3(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n535), .B(new_n575), .ZN(new_n614));
  XOR2_X1   g413(.A(new_n610), .B(KEYINPUT13), .Z(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n612), .A2(KEYINPUT94), .ZN(new_n617));
  NAND4_X1  g416(.A1(new_n608), .A2(new_n609), .A3(new_n610), .A4(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n613), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(KEYINPUT11), .B(G169gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(G197gat), .ZN(new_n621));
  XOR2_X1   g420(.A(G113gat), .B(G141gat), .Z(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(KEYINPUT12), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n619), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n613), .A2(new_n624), .A3(new_n616), .A4(new_n618), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(G230gat), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n630), .A2(new_n263), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n594), .A2(new_n547), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT10), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n592), .A2(new_n546), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n594), .A2(new_n547), .A3(KEYINPUT10), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n631), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n632), .A2(new_n634), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(new_n631), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(G176gat), .B(G204gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(KEYINPUT97), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(G120gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(new_n216), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n641), .B(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n629), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NOR3_X1   g447(.A1(new_n528), .A2(new_n606), .A3(new_n648), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n442), .B(KEYINPUT98), .Z(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(G1gat), .ZN(G1324gat));
  INV_X1    g452(.A(new_n649), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n654), .A2(new_n464), .ZN(new_n655));
  NAND2_X1  g454(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n656));
  INV_X1    g455(.A(G8gat), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n530), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n655), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(KEYINPUT42), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n660), .B1(new_n657), .B2(new_n655), .ZN(G1325gat));
  AOI21_X1  g460(.A(G15gat), .B1(new_n649), .B2(new_n475), .ZN(new_n662));
  INV_X1    g461(.A(new_n526), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n654), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n662), .B1(new_n664), .B2(G15gat), .ZN(G1326gat));
  INV_X1    g464(.A(new_n471), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n649), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(KEYINPUT43), .B(G22gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(G1327gat));
  NOR2_X1   g468(.A1(new_n560), .A2(new_n648), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NOR3_X1   g470(.A1(new_n528), .A2(new_n605), .A3(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n672), .A2(new_n565), .A3(new_n651), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(KEYINPUT45), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT99), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n675), .A2(KEYINPUT44), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n677), .B1(new_n528), .B2(new_n605), .ZN(new_n678));
  INV_X1    g477(.A(new_n605), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT99), .B(KEYINPUT44), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  AND2_X1   g480(.A1(new_n520), .A2(new_n527), .ZN(new_n682));
  AND3_X1   g481(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n683));
  AOI22_X1  g482(.A1(new_n475), .A2(new_n683), .B1(new_n456), .B2(KEYINPUT35), .ZN(new_n684));
  OAI211_X1 g483(.A(new_n679), .B(new_n681), .C1(new_n682), .C2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n678), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(KEYINPUT100), .B1(new_n686), .B2(new_n670), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT100), .ZN(new_n689));
  AOI211_X1 g488(.A(new_n689), .B(new_n671), .C1(new_n678), .C2(new_n685), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n650), .B1(new_n688), .B2(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n674), .B1(new_n692), .B2(new_n565), .ZN(G1328gat));
  NAND3_X1  g492(.A1(new_n672), .A2(new_n566), .A3(new_n460), .ZN(new_n694));
  XOR2_X1   g493(.A(new_n694), .B(KEYINPUT46), .Z(new_n695));
  AOI21_X1  g494(.A(new_n464), .B1(new_n688), .B2(new_n691), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n695), .B1(new_n696), .B2(new_n566), .ZN(G1329gat));
  NAND2_X1  g496(.A1(new_n686), .A2(new_n670), .ZN(new_n698));
  OAI21_X1  g497(.A(G43gat), .B1(new_n698), .B2(new_n663), .ZN(new_n699));
  INV_X1    g498(.A(G43gat), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n672), .A2(new_n700), .A3(new_n475), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n699), .A2(KEYINPUT47), .A3(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n701), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n526), .B1(new_n687), .B2(new_n690), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n703), .B1(new_n704), .B2(G43gat), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n702), .B1(new_n705), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g505(.A(G50gat), .ZN(new_n707));
  AND3_X1   g506(.A1(new_n672), .A2(new_n707), .A3(new_n666), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT101), .ZN(new_n709));
  OR2_X1    g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(G50gat), .B1(new_n698), .B2(new_n471), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n708), .A2(new_n709), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n710), .A2(new_n711), .A3(new_n712), .A4(KEYINPUT48), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n666), .B1(new_n687), .B2(new_n690), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n708), .B1(new_n714), .B2(G50gat), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n713), .B1(new_n715), .B2(KEYINPUT48), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(KEYINPUT102), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT102), .ZN(new_n718));
  OAI211_X1 g517(.A(new_n718), .B(new_n713), .C1(new_n715), .C2(KEYINPUT48), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n717), .A2(new_n719), .ZN(G1331gat));
  INV_X1    g519(.A(new_n646), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n528), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n606), .A2(new_n628), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(new_n651), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(G57gat), .ZN(G1332gat));
  INV_X1    g526(.A(KEYINPUT103), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n724), .B(new_n728), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n729), .A2(new_n464), .ZN(new_n730));
  NOR2_X1   g529(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n731));
  AND2_X1   g530(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n733), .B1(new_n730), .B2(new_n731), .ZN(G1333gat));
  OAI21_X1  g533(.A(G71gat), .B1(new_n729), .B2(new_n663), .ZN(new_n735));
  AOI21_X1  g534(.A(KEYINPUT104), .B1(new_n725), .B2(new_n475), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT104), .ZN(new_n737));
  INV_X1    g536(.A(new_n475), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n724), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n539), .B1(new_n736), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n735), .A2(new_n740), .ZN(new_n741));
  XOR2_X1   g540(.A(new_n741), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g541(.A1(new_n729), .A2(new_n471), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(new_n540), .ZN(G1335gat));
  NOR2_X1   g543(.A1(new_n560), .A2(new_n628), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n679), .B(new_n745), .C1(new_n682), .C2(new_n684), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT51), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n747), .A2(new_n721), .ZN(new_n748));
  AOI21_X1  g547(.A(G85gat), .B1(new_n748), .B2(new_n651), .ZN(new_n749));
  AND2_X1   g548(.A1(new_n686), .A2(new_n745), .ZN(new_n750));
  AND3_X1   g549(.A1(new_n750), .A2(new_n651), .A3(new_n646), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n749), .B1(G85gat), .B2(new_n751), .ZN(G1336gat));
  NAND3_X1  g551(.A1(new_n748), .A2(new_n403), .A3(new_n460), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT52), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n686), .A2(new_n460), .A3(new_n646), .A4(new_n745), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(G92gat), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n753), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n756), .A2(KEYINPUT105), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n756), .A2(KEYINPUT105), .ZN(new_n759));
  NOR2_X1   g558(.A1(KEYINPUT106), .A2(KEYINPUT51), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n746), .B(new_n760), .ZN(new_n761));
  AND4_X1   g560(.A1(new_n403), .A2(new_n761), .A3(new_n460), .A4(new_n646), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n758), .A2(new_n759), .A3(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n757), .B1(new_n763), .B2(new_n754), .ZN(G1337gat));
  NAND3_X1  g563(.A1(new_n748), .A2(new_n586), .A3(new_n475), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n750), .A2(new_n526), .A3(new_n646), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n765), .B1(new_n586), .B2(new_n766), .ZN(G1338gat));
  NAND4_X1  g566(.A1(new_n686), .A2(new_n666), .A3(new_n646), .A4(new_n745), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(G106gat), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT53), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n666), .A2(new_n587), .A3(new_n646), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n769), .B(new_n770), .C1(new_n747), .C2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(new_n771), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n761), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n769), .A2(new_n774), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n775), .A2(KEYINPUT107), .A3(KEYINPUT53), .ZN(new_n776));
  AOI21_X1  g575(.A(KEYINPUT107), .B1(new_n775), .B2(KEYINPUT53), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n772), .B1(new_n776), .B2(new_n777), .ZN(G1339gat));
  NOR2_X1   g577(.A1(new_n650), .A2(new_n460), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT113), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT108), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n635), .A2(new_n782), .A3(new_n636), .A4(new_n631), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n783), .A2(KEYINPUT54), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n635), .A2(new_n636), .A3(new_n631), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n785), .B1(new_n637), .B2(KEYINPUT108), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n645), .B1(new_n638), .B2(KEYINPUT54), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n781), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(KEYINPUT109), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n641), .A2(new_n645), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n788), .B1(new_n784), .B2(new_n786), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n791), .B1(new_n792), .B2(KEYINPUT55), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT109), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n794), .B(new_n781), .C1(new_n787), .C2(new_n788), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n790), .A2(new_n793), .A3(new_n795), .A4(new_n628), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT111), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n610), .B1(new_n608), .B2(new_n609), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n614), .A2(new_n615), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n623), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n627), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n646), .ZN(new_n802));
  AND3_X1   g601(.A1(new_n796), .A2(new_n797), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n797), .B1(new_n796), .B2(new_n802), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n803), .A2(new_n804), .A3(new_n679), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n790), .A2(new_n793), .A3(new_n801), .A4(new_n795), .ZN(new_n806));
  OR3_X1    g605(.A1(new_n806), .A2(KEYINPUT110), .A3(new_n605), .ZN(new_n807));
  OAI21_X1  g606(.A(KEYINPUT110), .B1(new_n806), .B2(new_n605), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(KEYINPUT112), .B1(new_n805), .B2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(new_n560), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n796), .A2(new_n802), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(KEYINPUT111), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n796), .A2(new_n797), .A3(new_n802), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n813), .A2(new_n605), .A3(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT112), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n815), .A2(new_n816), .A3(new_n808), .A4(new_n807), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n810), .A2(new_n811), .A3(new_n817), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n606), .A2(new_n646), .A3(new_n628), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n780), .B1(new_n821), .B2(new_n471), .ZN(new_n822));
  AOI211_X1 g621(.A(KEYINPUT113), .B(new_n666), .C1(new_n818), .C2(new_n820), .ZN(new_n823));
  OAI211_X1 g622(.A(new_n475), .B(new_n779), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  XNOR2_X1  g623(.A(new_n824), .B(KEYINPUT114), .ZN(new_n825));
  OAI21_X1  g624(.A(G113gat), .B1(new_n825), .B2(new_n629), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n650), .B1(new_n818), .B2(new_n820), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n386), .A2(new_n455), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n828), .A2(new_n460), .A3(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n830), .A2(new_n346), .A3(new_n628), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n826), .A2(new_n831), .ZN(G1340gat));
  OAI21_X1  g631(.A(G120gat), .B1(new_n825), .B2(new_n721), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n830), .A2(new_n348), .A3(new_n646), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(G1341gat));
  NOR3_X1   g634(.A1(new_n825), .A2(new_n345), .A3(new_n811), .ZN(new_n836));
  AOI21_X1  g635(.A(G127gat), .B1(new_n830), .B2(new_n560), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n836), .A2(new_n837), .ZN(G1342gat));
  OAI21_X1  g637(.A(G134gat), .B1(new_n825), .B2(new_n605), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n460), .A2(new_n605), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  NOR4_X1   g640(.A1(new_n828), .A2(G134gat), .A3(new_n829), .A4(new_n841), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n842), .B(KEYINPUT56), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n839), .A2(new_n843), .ZN(G1343gat));
  AOI21_X1  g643(.A(new_n471), .B1(new_n818), .B2(new_n820), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT57), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n663), .A2(new_n779), .ZN(new_n848));
  OR2_X1    g647(.A1(new_n789), .A2(KEYINPUT115), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n789), .A2(KEYINPUT115), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n849), .A2(new_n628), .A3(new_n793), .A4(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n679), .B1(new_n851), .B2(new_n802), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n809), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n853), .A2(new_n560), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n666), .B1(new_n854), .B2(new_n819), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n848), .B1(new_n855), .B2(KEYINPUT57), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n847), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(G141gat), .B1(new_n857), .B2(new_n629), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n471), .B1(new_n828), .B2(KEYINPUT116), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT116), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n526), .B1(new_n827), .B2(new_n860), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n859), .A2(new_n218), .A3(new_n464), .A4(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n858), .B1(new_n862), .B2(new_n629), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(KEYINPUT117), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT117), .ZN(new_n865));
  OAI211_X1 g664(.A(new_n865), .B(new_n858), .C1(new_n862), .C2(new_n629), .ZN(new_n866));
  AND3_X1   g665(.A1(new_n864), .A2(KEYINPUT58), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(KEYINPUT58), .B1(new_n864), .B2(new_n866), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n867), .A2(new_n868), .ZN(G1344gat));
  AND3_X1   g668(.A1(new_n859), .A2(new_n464), .A3(new_n861), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n870), .A2(new_n216), .A3(new_n646), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT59), .ZN(new_n872));
  OR2_X1    g671(.A1(new_n845), .A2(new_n846), .ZN(new_n873));
  INV_X1    g672(.A(new_n852), .ZN(new_n874));
  AND3_X1   g673(.A1(new_n790), .A2(new_n793), .A3(new_n795), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n875), .A2(new_n679), .A3(new_n801), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n560), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n846), .B(new_n666), .C1(new_n819), .C2(new_n877), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n873), .A2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(new_n848), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n879), .A2(new_n646), .A3(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT118), .ZN(new_n882));
  OR2_X1    g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n216), .B1(new_n881), .B2(new_n882), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n872), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(new_n857), .ZN(new_n886));
  AOI211_X1 g685(.A(KEYINPUT59), .B(new_n216), .C1(new_n886), .C2(new_n646), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n871), .B1(new_n885), .B2(new_n887), .ZN(G1345gat));
  NAND3_X1  g687(.A1(new_n870), .A2(new_n213), .A3(new_n560), .ZN(new_n889));
  OAI21_X1  g688(.A(G155gat), .B1(new_n857), .B2(new_n811), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  XOR2_X1   g690(.A(new_n891), .B(KEYINPUT119), .Z(G1346gat));
  NAND4_X1  g691(.A1(new_n859), .A2(new_n212), .A3(new_n840), .A4(new_n861), .ZN(new_n893));
  OR3_X1    g692(.A1(new_n857), .A2(KEYINPUT120), .A3(new_n605), .ZN(new_n894));
  OAI21_X1  g693(.A(KEYINPUT120), .B1(new_n857), .B2(new_n605), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n893), .B1(new_n896), .B2(new_n212), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT121), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n897), .B(new_n898), .ZN(G1347gat));
  NOR3_X1   g698(.A1(new_n829), .A2(new_n651), .A3(new_n464), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n821), .A2(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n902), .A2(new_n329), .A3(new_n628), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n651), .A2(new_n464), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(new_n475), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(KEYINPUT122), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n906), .B1(new_n822), .B2(new_n823), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT123), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OAI211_X1 g708(.A(KEYINPUT123), .B(new_n906), .C1(new_n822), .C2(new_n823), .ZN(new_n910));
  AND3_X1   g709(.A1(new_n909), .A2(new_n628), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n903), .B1(new_n911), .B2(new_n329), .ZN(G1348gat));
  NAND4_X1  g711(.A1(new_n909), .A2(G176gat), .A3(new_n646), .A4(new_n910), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n330), .B1(new_n901), .B2(new_n721), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n913), .A2(new_n914), .ZN(G1349gat));
  AND3_X1   g714(.A1(new_n902), .A2(new_n326), .A3(new_n560), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n909), .A2(new_n560), .A3(new_n910), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n916), .B1(new_n917), .B2(G183gat), .ZN(new_n918));
  NAND2_X1  g717(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n918), .B(new_n919), .ZN(G1350gat));
  NAND3_X1  g719(.A1(new_n909), .A2(new_n679), .A3(new_n910), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(G190gat), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(KEYINPUT125), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT125), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n921), .A2(new_n924), .A3(G190gat), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n923), .A2(KEYINPUT61), .A3(new_n925), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n902), .A2(new_n320), .A3(new_n679), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT61), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n922), .A2(KEYINPUT125), .A3(new_n928), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n926), .A2(new_n927), .A3(new_n929), .ZN(G1351gat));
  NAND2_X1  g729(.A1(new_n663), .A2(new_n904), .ZN(new_n931));
  INV_X1    g730(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n879), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g732(.A(G197gat), .B1(new_n933), .B2(new_n629), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n845), .A2(new_n932), .ZN(new_n935));
  OR3_X1    g734(.A1(new_n935), .A2(G197gat), .A3(new_n629), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n936), .ZN(G1352gat));
  NAND3_X1  g736(.A1(new_n879), .A2(new_n646), .A3(new_n932), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(G204gat), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n935), .A2(G204gat), .A3(new_n721), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT62), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n941), .ZN(G1353gat));
  OAI21_X1  g741(.A(G211gat), .B1(new_n933), .B2(new_n811), .ZN(new_n943));
  OR2_X1    g742(.A1(new_n943), .A2(KEYINPUT63), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(KEYINPUT63), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n935), .A2(new_n244), .A3(new_n811), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n946), .B(KEYINPUT126), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n944), .A2(new_n945), .A3(new_n947), .ZN(G1354gat));
  OAI21_X1  g747(.A(new_n228), .B1(new_n935), .B2(new_n605), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n605), .A2(new_n228), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT127), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n949), .B1(new_n933), .B2(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(new_n952), .ZN(G1355gat));
endmodule


