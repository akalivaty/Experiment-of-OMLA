//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 0 1 1 0 0 0 0 1 1 1 0 1 1 0 0 0 1 1 0 1 0 1 0 0 1 1 0 0 1 1 1 0 1 0 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n751, new_n753, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n812, new_n814,
    new_n815, new_n816, new_n817, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n864, new_n865, new_n866, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n875, new_n876, new_n878,
    new_n879, new_n880, new_n881, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924;
  INV_X1    g000(.A(KEYINPUT9), .ZN(new_n202));
  INV_X1    g001(.A(G71gat), .ZN(new_n203));
  INV_X1    g002(.A(G78gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n205), .A2(KEYINPUT93), .ZN(new_n206));
  XOR2_X1   g005(.A(G71gat), .B(G78gat), .Z(new_n207));
  NOR2_X1   g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G57gat), .B(G64gat), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n209), .B1(KEYINPUT93), .B2(new_n205), .ZN(new_n210));
  OR2_X1    g009(.A1(new_n209), .A2(new_n202), .ZN(new_n211));
  AOI22_X1  g010(.A1(new_n208), .A2(new_n210), .B1(new_n211), .B2(new_n207), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n212), .A2(KEYINPUT21), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n213), .B(G211gat), .ZN(new_n214));
  XNOR2_X1  g013(.A(G127gat), .B(G155gat), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n214), .B(new_n215), .ZN(new_n216));
  XOR2_X1   g015(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n217));
  XNOR2_X1  g016(.A(new_n216), .B(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(G15gat), .B(G22gat), .ZN(new_n220));
  INV_X1    g019(.A(G1gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT16), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n223), .B1(G1gat), .B2(new_n220), .ZN(new_n224));
  XOR2_X1   g023(.A(new_n224), .B(G8gat), .Z(new_n225));
  INV_X1    g024(.A(KEYINPUT21), .ZN(new_n226));
  INV_X1    g025(.A(new_n212), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n225), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n228), .B(G183gat), .ZN(new_n229));
  INV_X1    g028(.A(G231gat), .ZN(new_n230));
  INV_X1    g029(.A(G233gat), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n229), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(G183gat), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n228), .B(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n234), .A2(G231gat), .A3(G233gat), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT94), .B(KEYINPUT95), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n232), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n237), .B1(new_n232), .B2(new_n235), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n219), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n240), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n242), .A2(new_n218), .A3(new_n238), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(G50gat), .ZN(new_n246));
  OR2_X1    g045(.A1(new_n246), .A2(G43gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(G43gat), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n247), .A2(KEYINPUT15), .A3(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(KEYINPUT89), .B(G43gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(new_n246), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT15), .B1(new_n251), .B2(new_n247), .ZN(new_n252));
  NOR2_X1   g051(.A1(G29gat), .A2(G36gat), .ZN(new_n253));
  OR2_X1    g052(.A1(new_n253), .A2(KEYINPUT14), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(KEYINPUT14), .ZN(new_n255));
  INV_X1    g054(.A(G36gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(KEYINPUT88), .B(G29gat), .ZN(new_n257));
  OAI211_X1 g056(.A(new_n254), .B(new_n255), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n249), .B1(new_n252), .B2(new_n258), .ZN(new_n259));
  OR2_X1    g058(.A1(new_n258), .A2(new_n249), .ZN(new_n260));
  AND2_X1   g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT17), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n261), .A2(KEYINPUT90), .A3(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT90), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n259), .A2(new_n260), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n264), .B1(new_n265), .B2(KEYINPUT17), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n265), .A2(KEYINPUT17), .ZN(new_n268));
  NAND2_X1  g067(.A1(G99gat), .A2(G106gat), .ZN(new_n269));
  INV_X1    g068(.A(G85gat), .ZN(new_n270));
  INV_X1    g069(.A(G92gat), .ZN(new_n271));
  AOI22_X1  g070(.A1(KEYINPUT8), .A2(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT7), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n273), .B1(new_n270), .B2(new_n271), .ZN(new_n274));
  NAND3_X1  g073(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n272), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  XOR2_X1   g075(.A(G99gat), .B(G106gat), .Z(new_n277));
  NAND3_X1  g076(.A1(new_n276), .A2(KEYINPUT96), .A3(new_n277), .ZN(new_n278));
  OR2_X1    g077(.A1(new_n276), .A2(new_n277), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT96), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n276), .A2(new_n277), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n267), .A2(new_n268), .A3(new_n278), .A4(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n278), .ZN(new_n284));
  AND2_X1   g083(.A1(G232gat), .A2(G233gat), .ZN(new_n285));
  AOI22_X1  g084(.A1(new_n261), .A2(new_n284), .B1(KEYINPUT41), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G190gat), .B(G218gat), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n287), .B(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n285), .A2(KEYINPUT41), .ZN(new_n291));
  XNOR2_X1  g090(.A(G134gat), .B(G162gat), .ZN(new_n292));
  XOR2_X1   g091(.A(new_n291), .B(new_n292), .Z(new_n293));
  NAND2_X1  g092(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n287), .B(new_n288), .ZN(new_n295));
  INV_X1    g094(.A(new_n293), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  AND2_X1   g098(.A1(G230gat), .A2(G233gat), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT97), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n301), .B1(new_n284), .B2(new_n212), .ZN(new_n302));
  NAND4_X1  g101(.A1(new_n227), .A2(new_n282), .A3(KEYINPUT97), .A4(new_n278), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AND2_X1   g103(.A1(new_n279), .A2(new_n281), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(new_n212), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT98), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT98), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n305), .A2(new_n308), .A3(new_n212), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT10), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n304), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n284), .A2(KEYINPUT10), .A3(new_n212), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n300), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n300), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n315), .B1(new_n304), .B2(new_n310), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G120gat), .B(G148gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(G176gat), .B(G204gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n318), .B(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n317), .B(new_n321), .ZN(new_n322));
  NOR3_X1   g121(.A1(new_n245), .A2(new_n299), .A3(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT87), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT73), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT23), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n327), .A2(G169gat), .ZN(new_n328));
  INV_X1    g127(.A(G176gat), .ZN(new_n329));
  AND2_X1   g128(.A1(new_n329), .A2(KEYINPUT64), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n329), .A2(KEYINPUT64), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n328), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(G169gat), .A2(G176gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(G183gat), .A2(G190gat), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT24), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n337));
  INV_X1    g136(.A(G190gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n233), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n336), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(G169gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(new_n329), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(new_n327), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n332), .A2(new_n333), .A3(new_n340), .A4(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT25), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AOI22_X1  g145(.A1(new_n342), .A2(new_n327), .B1(KEYINPUT65), .B2(new_n333), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n328), .A2(new_n329), .ZN(new_n348));
  AND2_X1   g147(.A1(G169gat), .A2(G176gat), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT65), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n345), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n347), .A2(new_n340), .A3(new_n348), .A4(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(KEYINPUT66), .ZN(new_n353));
  OAI21_X1  g152(.A(KEYINPUT25), .B1(new_n333), .B2(KEYINPUT65), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n354), .B1(new_n329), .B2(new_n328), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT66), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n355), .A2(new_n356), .A3(new_n340), .A4(new_n347), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n346), .A2(new_n353), .A3(new_n357), .ZN(new_n358));
  AND2_X1   g157(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n359));
  NOR2_X1   g158(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT67), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n338), .B1(new_n362), .B2(KEYINPUT28), .ZN(new_n363));
  NOR3_X1   g162(.A1(new_n361), .A2(KEYINPUT68), .A3(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT68), .ZN(new_n365));
  XNOR2_X1  g164(.A(KEYINPUT27), .B(G183gat), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT28), .ZN(new_n367));
  AOI21_X1  g166(.A(G190gat), .B1(new_n367), .B2(KEYINPUT67), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n365), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  OAI22_X1  g168(.A1(new_n364), .A2(new_n369), .B1(KEYINPUT67), .B2(new_n367), .ZN(new_n370));
  NOR2_X1   g169(.A1(G169gat), .A2(G176gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n371), .B(KEYINPUT26), .ZN(new_n372));
  AOI22_X1  g171(.A1(new_n372), .A2(new_n333), .B1(G183gat), .B2(G190gat), .ZN(new_n373));
  OAI21_X1  g172(.A(KEYINPUT68), .B1(new_n361), .B2(new_n363), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n366), .A2(new_n365), .A3(new_n368), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n374), .A2(new_n362), .A3(new_n375), .A4(KEYINPUT28), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n370), .A2(new_n373), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n358), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(G113gat), .B(G120gat), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n379), .A2(KEYINPUT1), .ZN(new_n380));
  XNOR2_X1  g179(.A(G127gat), .B(G134gat), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  OR2_X1    g181(.A1(new_n381), .A2(KEYINPUT69), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n381), .A2(KEYINPUT69), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n379), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(KEYINPUT70), .B(KEYINPUT1), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n382), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n378), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(G227gat), .A2(G233gat), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n358), .A2(new_n387), .A3(new_n377), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n389), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(KEYINPUT34), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT34), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n389), .A2(new_n394), .A3(new_n390), .A4(new_n391), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n390), .ZN(new_n397));
  AND3_X1   g196(.A1(new_n358), .A2(new_n387), .A3(new_n377), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n387), .B1(new_n358), .B2(new_n377), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n397), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  XOR2_X1   g199(.A(G15gat), .B(G43gat), .Z(new_n401));
  XOR2_X1   g200(.A(G71gat), .B(G99gat), .Z(new_n402));
  XOR2_X1   g201(.A(new_n401), .B(new_n402), .Z(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  OR2_X1    g203(.A1(new_n404), .A2(KEYINPUT71), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(KEYINPUT71), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n405), .A2(KEYINPUT33), .A3(new_n406), .ZN(new_n407));
  AND3_X1   g206(.A1(new_n400), .A2(KEYINPUT32), .A3(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT32), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT33), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n404), .B1(new_n400), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n396), .B1(new_n408), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n390), .B1(new_n389), .B2(new_n391), .ZN(new_n413));
  INV_X1    g212(.A(new_n410), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n403), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n400), .A2(KEYINPUT32), .A3(new_n407), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n415), .A2(new_n416), .A3(new_n393), .A4(new_n395), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n412), .A2(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(KEYINPUT72), .B(KEYINPUT36), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n326), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  AOI211_X1 g221(.A(KEYINPUT73), .B(new_n419), .C1(new_n412), .C2(new_n417), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  AND3_X1   g223(.A1(new_n412), .A2(KEYINPUT36), .A3(new_n417), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n422), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(G226gat), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n428), .A2(new_n231), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT29), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n378), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n358), .A2(new_n377), .A3(new_n430), .ZN(new_n434));
  XNOR2_X1  g233(.A(G197gat), .B(G204gat), .ZN(new_n435));
  INV_X1    g234(.A(G211gat), .ZN(new_n436));
  INV_X1    g235(.A(G218gat), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n435), .B1(KEYINPUT22), .B2(new_n438), .ZN(new_n439));
  XOR2_X1   g238(.A(G211gat), .B(G218gat), .Z(new_n440));
  XNOR2_X1  g239(.A(new_n439), .B(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n433), .A2(new_n434), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT75), .ZN(new_n443));
  XOR2_X1   g242(.A(G64gat), .B(G92gat), .Z(new_n444));
  XNOR2_X1  g243(.A(G8gat), .B(G36gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n444), .B(new_n445), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n441), .B(KEYINPUT74), .ZN(new_n447));
  INV_X1    g246(.A(new_n434), .ZN(new_n448));
  AOI22_X1  g247(.A1(new_n358), .A2(new_n377), .B1(new_n431), .B2(new_n430), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT75), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n433), .A2(new_n451), .A3(new_n434), .A4(new_n441), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n443), .A2(new_n446), .A3(new_n450), .A4(new_n452), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n453), .A2(KEYINPUT30), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT30), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n443), .A2(new_n450), .A3(new_n452), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n446), .B(KEYINPUT76), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n455), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n454), .B1(new_n453), .B2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(G155gat), .ZN(new_n460));
  INV_X1    g259(.A(G162gat), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(G155gat), .A2(G162gat), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  XNOR2_X1  g263(.A(new_n464), .B(KEYINPUT77), .ZN(new_n465));
  INV_X1    g264(.A(G148gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(G141gat), .ZN(new_n467));
  INV_X1    g266(.A(G141gat), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(G148gat), .ZN(new_n469));
  AOI22_X1  g268(.A1(new_n467), .A2(new_n469), .B1(KEYINPUT2), .B2(new_n463), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT82), .ZN(new_n473));
  OR2_X1    g272(.A1(KEYINPUT80), .A2(G162gat), .ZN(new_n474));
  NAND2_X1  g273(.A1(KEYINPUT80), .A2(G162gat), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n474), .A2(G155gat), .A3(new_n475), .ZN(new_n476));
  AND3_X1   g275(.A1(new_n476), .A2(KEYINPUT81), .A3(KEYINPUT2), .ZN(new_n477));
  AOI21_X1  g276(.A(KEYINPUT81), .B1(new_n476), .B2(KEYINPUT2), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT78), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n480), .A2(G141gat), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n468), .A2(KEYINPUT78), .ZN(new_n482));
  OAI21_X1  g281(.A(G148gat), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  AND2_X1   g282(.A1(G155gat), .A2(G162gat), .ZN(new_n484));
  NOR2_X1   g283(.A1(G155gat), .A2(G162gat), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT79), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT79), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n462), .A2(new_n487), .A3(new_n463), .ZN(new_n488));
  AOI22_X1  g287(.A1(new_n483), .A2(new_n467), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n473), .B1(new_n479), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT81), .ZN(new_n491));
  AND2_X1   g290(.A1(KEYINPUT80), .A2(G162gat), .ZN(new_n492));
  NOR2_X1   g291(.A1(KEYINPUT80), .A2(G162gat), .ZN(new_n493));
  NOR3_X1   g292(.A1(new_n492), .A2(new_n493), .A3(new_n460), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT2), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n491), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n476), .A2(KEYINPUT81), .A3(KEYINPUT2), .ZN(new_n497));
  AND4_X1   g296(.A1(new_n473), .A2(new_n489), .A3(new_n496), .A4(new_n497), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n472), .B(new_n387), .C1(new_n490), .C2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT4), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT83), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n483), .A2(new_n467), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n488), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n496), .A2(new_n502), .A3(new_n503), .A4(new_n497), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(KEYINPUT82), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n489), .A2(new_n473), .A3(new_n496), .A4(new_n497), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n471), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT4), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n507), .A2(new_n508), .A3(new_n387), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n500), .A2(new_n501), .A3(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n472), .B1(new_n490), .B2(new_n498), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT3), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n505), .A2(new_n506), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT3), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n513), .A2(new_n514), .A3(new_n472), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n512), .A2(new_n388), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(G225gat), .A2(G233gat), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n508), .B1(new_n507), .B2(new_n387), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(KEYINPUT83), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n510), .A2(new_n516), .A3(new_n517), .A4(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT5), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n511), .A2(new_n388), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(new_n499), .ZN(new_n523));
  INV_X1    g322(.A(new_n517), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n521), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n514), .B1(new_n513), .B2(new_n472), .ZN(new_n526));
  AOI211_X1 g325(.A(KEYINPUT3), .B(new_n471), .C1(new_n505), .C2(new_n506), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AOI22_X1  g327(.A1(new_n528), .A2(new_n388), .B1(new_n500), .B2(new_n509), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n524), .A2(KEYINPUT5), .ZN(new_n530));
  AOI22_X1  g329(.A1(new_n520), .A2(new_n525), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(G1gat), .B(G29gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(new_n270), .ZN(new_n533));
  XNOR2_X1  g332(.A(KEYINPUT0), .B(G57gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(KEYINPUT6), .B1(new_n531), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n525), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n529), .A2(new_n530), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n535), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n536), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n539), .A2(KEYINPUT6), .A3(new_n540), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n459), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G78gat), .B(G106gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(KEYINPUT31), .B(G50gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n441), .B1(new_n515), .B2(new_n431), .ZN(new_n548));
  AOI21_X1  g347(.A(KEYINPUT3), .B1(new_n441), .B2(new_n431), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n507), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(G228gat), .ZN(new_n551));
  OAI22_X1  g350(.A1(new_n548), .A2(new_n550), .B1(new_n551), .B2(new_n231), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n447), .B1(new_n527), .B2(KEYINPUT29), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n551), .A2(new_n231), .ZN(new_n554));
  INV_X1    g353(.A(new_n550), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(G22gat), .ZN(new_n557));
  AND3_X1   g356(.A1(new_n552), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n557), .B1(new_n552), .B2(new_n556), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n547), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n552), .A2(new_n556), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(G22gat), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n552), .A2(new_n556), .A3(new_n557), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n547), .A2(KEYINPUT84), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n559), .A2(KEYINPUT84), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n560), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n427), .B1(new_n544), .B2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT40), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n500), .A2(new_n509), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n517), .B1(new_n571), .B2(new_n516), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n522), .A2(new_n517), .A3(new_n499), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT39), .ZN(new_n575));
  NOR3_X1   g374(.A1(new_n572), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n499), .A2(KEYINPUT4), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n577), .A2(new_n518), .ZN(new_n578));
  NOR3_X1   g377(.A1(new_n526), .A2(new_n527), .A3(new_n387), .ZN(new_n579));
  OAI211_X1 g378(.A(new_n575), .B(new_n524), .C1(new_n578), .C2(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n535), .B(KEYINPUT85), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n570), .B1(new_n576), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n539), .A2(new_n581), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n581), .B1(new_n572), .B2(new_n575), .ZN(new_n586));
  OAI211_X1 g385(.A(KEYINPUT39), .B(new_n573), .C1(new_n529), .C2(new_n517), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n586), .A2(new_n587), .A3(KEYINPUT40), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n584), .A2(new_n585), .A3(new_n459), .A4(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT86), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n536), .A2(new_n585), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT38), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n446), .B1(new_n456), .B2(KEYINPUT37), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT37), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n443), .A2(new_n594), .A3(new_n450), .A4(new_n452), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n592), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n595), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n441), .B1(new_n448), .B2(new_n449), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n433), .A2(new_n434), .A3(new_n447), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n598), .A2(new_n599), .A3(KEYINPUT37), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n600), .A2(new_n592), .A3(new_n457), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n453), .B1(new_n597), .B2(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n596), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n591), .A2(new_n603), .A3(new_n543), .ZN(new_n604));
  AND2_X1   g403(.A1(new_n604), .A2(new_n568), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n569), .B1(new_n590), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n543), .ZN(new_n607));
  NOR4_X1   g406(.A1(new_n567), .A2(KEYINPUT35), .A3(new_n459), .A4(new_n418), .ZN(new_n608));
  AND2_X1   g407(.A1(new_n412), .A2(new_n417), .ZN(new_n609));
  AND4_X1   g408(.A1(new_n560), .A2(new_n565), .A3(new_n609), .A4(new_n566), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n537), .A2(new_n535), .A3(new_n538), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT6), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n531), .A2(new_n535), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n543), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n459), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n610), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  AOI22_X1  g416(.A1(new_n607), .A2(new_n608), .B1(new_n617), .B2(KEYINPUT35), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n325), .B1(new_n606), .B2(new_n618), .ZN(new_n619));
  OR2_X1    g418(.A1(new_n225), .A2(new_n265), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT91), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n621), .B1(new_n225), .B2(new_n265), .ZN(new_n622));
  XOR2_X1   g421(.A(new_n620), .B(new_n622), .Z(new_n623));
  NAND2_X1  g422(.A1(G229gat), .A2(G233gat), .ZN(new_n624));
  XOR2_X1   g423(.A(new_n624), .B(KEYINPUT13), .Z(new_n625));
  NAND2_X1  g424(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n267), .A2(new_n225), .A3(new_n268), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n627), .A2(new_n624), .A3(new_n620), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT18), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n627), .A2(KEYINPUT18), .A3(new_n624), .A4(new_n620), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n626), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(G113gat), .B(G141gat), .ZN(new_n633));
  INV_X1    g432(.A(G197gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(KEYINPUT11), .B(G169gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g436(.A(new_n637), .B(KEYINPUT12), .Z(new_n638));
  NAND2_X1  g437(.A1(new_n632), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n638), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n626), .A2(new_n630), .A3(new_n631), .A4(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  AND3_X1   g441(.A1(new_n586), .A2(new_n587), .A3(KEYINPUT40), .ZN(new_n643));
  AOI21_X1  g442(.A(KEYINPUT40), .B1(new_n586), .B2(new_n587), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n645), .A2(KEYINPUT86), .A3(new_n459), .A4(new_n585), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT86), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n589), .A2(new_n647), .ZN(new_n648));
  NAND4_X1  g447(.A1(new_n646), .A2(new_n648), .A3(new_n568), .A4(new_n604), .ZN(new_n649));
  NOR3_X1   g448(.A1(new_n421), .A2(new_n423), .A3(new_n425), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n615), .A2(new_n616), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n650), .B1(new_n651), .B2(new_n567), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n617), .A2(KEYINPUT35), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT35), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n607), .A2(new_n610), .A3(new_n655), .A4(new_n616), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n653), .A2(new_n657), .A3(KEYINPUT87), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n619), .A2(new_n642), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(KEYINPUT92), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT92), .ZN(new_n661));
  NAND4_X1  g460(.A1(new_n619), .A2(new_n661), .A3(new_n642), .A4(new_n658), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n324), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n615), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g465(.A1(new_n663), .A2(new_n459), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT42), .ZN(new_n668));
  XNOR2_X1  g467(.A(KEYINPUT16), .B(G8gat), .ZN(new_n669));
  OR3_X1    g468(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n667), .A2(G8gat), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n668), .B1(new_n667), .B2(new_n669), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(G1325gat));
  OR2_X1    g472(.A1(new_n650), .A2(KEYINPUT100), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n650), .A2(KEYINPUT100), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n663), .A2(G15gat), .A3(new_n676), .ZN(new_n677));
  AOI211_X1 g476(.A(KEYINPUT99), .B(G15gat), .C1(new_n663), .C2(new_n609), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT99), .ZN(new_n679));
  AND3_X1   g478(.A1(new_n653), .A2(KEYINPUT87), .A3(new_n657), .ZN(new_n680));
  AOI21_X1  g479(.A(KEYINPUT87), .B1(new_n653), .B2(new_n657), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n661), .B1(new_n682), .B2(new_n642), .ZN(new_n683));
  INV_X1    g482(.A(new_n662), .ZN(new_n684));
  OAI211_X1 g483(.A(new_n609), .B(new_n323), .C1(new_n683), .C2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(G15gat), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n679), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n677), .B1(new_n678), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(KEYINPUT101), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT101), .ZN(new_n690));
  OAI211_X1 g489(.A(new_n690), .B(new_n677), .C1(new_n678), .C2(new_n687), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n689), .A2(new_n691), .ZN(G1326gat));
  NAND2_X1  g491(.A1(new_n663), .A2(new_n567), .ZN(new_n693));
  XNOR2_X1  g492(.A(KEYINPUT43), .B(G22gat), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n693), .B(new_n694), .ZN(G1327gat));
  AOI21_X1  g494(.A(new_n322), .B1(new_n660), .B2(new_n662), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n244), .A2(new_n298), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n696), .A2(new_n664), .A3(new_n257), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT45), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n682), .A2(KEYINPUT44), .A3(new_n299), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n244), .B(KEYINPUT102), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n298), .B1(new_n653), .B2(new_n657), .ZN(new_n703));
  OR2_X1    g502(.A1(new_n703), .A2(KEYINPUT44), .ZN(new_n704));
  INV_X1    g503(.A(new_n642), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n705), .A2(new_n322), .ZN(new_n706));
  NAND4_X1  g505(.A1(new_n700), .A2(new_n702), .A3(new_n704), .A4(new_n706), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n707), .A2(new_n615), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n699), .B1(new_n257), .B2(new_n708), .ZN(G1328gat));
  AND2_X1   g508(.A1(new_n696), .A2(new_n697), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n616), .A2(G36gat), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(KEYINPUT103), .B1(new_n712), .B2(KEYINPUT46), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT46), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n707), .A2(new_n616), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n714), .B1(new_n715), .B2(new_n256), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(new_n712), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT103), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n710), .A2(new_n718), .A3(new_n714), .A4(new_n711), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n713), .A2(new_n717), .A3(new_n719), .ZN(G1329gat));
  INV_X1    g519(.A(new_n676), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n250), .B1(new_n707), .B2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n250), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n696), .A2(new_n723), .A3(new_n609), .A4(new_n697), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT104), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n722), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT47), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  OAI211_X1 g527(.A(KEYINPUT47), .B(new_n250), .C1(new_n707), .C2(new_n427), .ZN(new_n729));
  OAI211_X1 g528(.A(new_n729), .B(new_n724), .C1(new_n725), .C2(KEYINPUT47), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n730), .ZN(G1330gat));
  OAI21_X1  g530(.A(G50gat), .B1(new_n707), .B2(new_n568), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n696), .A2(new_n246), .A3(new_n567), .A4(new_n697), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  XOR2_X1   g533(.A(new_n734), .B(KEYINPUT48), .Z(G1331gat));
  NAND2_X1  g534(.A1(new_n653), .A2(new_n657), .ZN(new_n736));
  INV_X1    g535(.A(new_n322), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n737), .A2(new_n642), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  AND3_X1   g538(.A1(new_n739), .A2(new_n244), .A3(new_n298), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n664), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g541(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n740), .A2(new_n459), .A3(new_n743), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT105), .ZN(new_n745));
  NOR2_X1   g544(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n745), .B(new_n746), .ZN(G1333gat));
  INV_X1    g546(.A(new_n740), .ZN(new_n748));
  OAI21_X1  g547(.A(G71gat), .B1(new_n748), .B2(new_n721), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n740), .A2(new_n203), .A3(new_n609), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  XOR2_X1   g550(.A(new_n751), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g551(.A1(new_n740), .A2(new_n567), .ZN(new_n753));
  XNOR2_X1  g552(.A(KEYINPUT106), .B(G78gat), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n753), .B(new_n754), .ZN(G1335gat));
  NAND3_X1  g554(.A1(new_n736), .A2(new_n705), .A3(new_n697), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT51), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n757), .A2(new_n737), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n758), .A2(new_n270), .A3(new_n664), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n700), .A2(new_n245), .A3(new_n704), .A4(new_n738), .ZN(new_n760));
  OAI21_X1  g559(.A(G85gat), .B1(new_n760), .B2(new_n615), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n759), .A2(new_n761), .ZN(G1336gat));
  OAI21_X1  g561(.A(G92gat), .B1(new_n760), .B2(new_n616), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n322), .A2(new_n271), .A3(new_n459), .ZN(new_n764));
  XOR2_X1   g563(.A(new_n764), .B(KEYINPUT108), .Z(new_n765));
  OAI22_X1  g564(.A1(new_n763), .A2(KEYINPUT107), .B1(new_n757), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(KEYINPUT52), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT52), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n763), .B1(KEYINPUT107), .B2(new_n768), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n757), .A2(KEYINPUT52), .A3(new_n764), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n767), .B1(new_n769), .B2(new_n770), .ZN(G1337gat));
  INV_X1    g570(.A(G99gat), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n758), .A2(new_n772), .A3(new_n609), .ZN(new_n773));
  OAI21_X1  g572(.A(G99gat), .B1(new_n760), .B2(new_n721), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(G1338gat));
  OAI21_X1  g574(.A(G106gat), .B1(new_n760), .B2(new_n568), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT109), .ZN(new_n777));
  OR3_X1    g576(.A1(new_n568), .A2(new_n737), .A3(G106gat), .ZN(new_n778));
  XOR2_X1   g577(.A(new_n778), .B(KEYINPUT110), .Z(new_n779));
  OAI22_X1  g578(.A1(new_n776), .A2(new_n777), .B1(new_n757), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(KEYINPUT53), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT53), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n776), .B1(new_n777), .B2(new_n782), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n757), .A2(KEYINPUT53), .A3(new_n778), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n781), .B1(new_n783), .B2(new_n784), .ZN(G1339gat));
  NAND4_X1  g584(.A1(new_n244), .A2(new_n705), .A3(new_n298), .A4(new_n737), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT55), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n312), .A2(new_n300), .A3(new_n313), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(KEYINPUT54), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n789), .A2(new_n314), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT54), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n314), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(new_n320), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n787), .B1(new_n790), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n317), .A2(new_n321), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n321), .B1(new_n314), .B2(new_n791), .ZN(new_n796));
  OAI211_X1 g595(.A(new_n796), .B(KEYINPUT55), .C1(new_n314), .C2(new_n789), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n794), .A2(new_n795), .A3(new_n797), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n623), .A2(new_n625), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n624), .B1(new_n627), .B2(new_n620), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n637), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n294), .A2(new_n297), .A3(new_n641), .A4(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n798), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n642), .A2(new_n795), .A3(new_n794), .A4(new_n797), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n322), .A2(new_n641), .A3(new_n801), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n803), .B1(new_n806), .B2(new_n298), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n786), .B1(new_n807), .B2(new_n701), .ZN(new_n808));
  AND4_X1   g607(.A1(new_n664), .A2(new_n808), .A3(new_n616), .A4(new_n610), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n642), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n810), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g610(.A1(new_n809), .A2(new_n322), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n812), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g612(.A1(new_n809), .A2(new_n244), .ZN(new_n814));
  XOR2_X1   g613(.A(new_n814), .B(KEYINPUT111), .Z(new_n815));
  INV_X1    g614(.A(G127gat), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n702), .A2(new_n816), .ZN(new_n817));
  AOI22_X1  g616(.A1(new_n815), .A2(new_n816), .B1(new_n809), .B2(new_n817), .ZN(G1342gat));
  NAND2_X1  g617(.A1(new_n809), .A2(new_n299), .ZN(new_n819));
  OR2_X1    g618(.A1(new_n819), .A2(G134gat), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n820), .A2(KEYINPUT56), .ZN(new_n821));
  OR2_X1    g620(.A1(new_n821), .A2(KEYINPUT112), .ZN(new_n822));
  OR2_X1    g621(.A1(new_n820), .A2(KEYINPUT56), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n819), .A2(G134gat), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n821), .A2(KEYINPUT112), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n822), .A2(new_n823), .A3(new_n824), .A4(new_n825), .ZN(G1343gat));
  NAND2_X1  g625(.A1(new_n664), .A2(new_n616), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n827), .A2(new_n650), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n808), .A2(new_n567), .ZN(new_n830));
  XNOR2_X1  g629(.A(KEYINPUT113), .B(KEYINPUT57), .ZN(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n299), .B1(new_n804), .B2(new_n805), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n245), .B1(new_n834), .B2(new_n803), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n786), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n836), .A2(KEYINPUT57), .A3(new_n567), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n829), .B1(new_n833), .B2(new_n837), .ZN(new_n838));
  AOI211_X1 g637(.A(new_n481), .B(new_n482), .C1(new_n838), .C2(new_n642), .ZN(new_n839));
  INV_X1    g638(.A(new_n827), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n676), .A2(new_n568), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n808), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n842), .A2(G141gat), .A3(new_n705), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n839), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g643(.A(KEYINPUT114), .B(KEYINPUT58), .ZN(new_n845));
  XNOR2_X1  g644(.A(new_n844), .B(new_n845), .ZN(G1344gat));
  INV_X1    g645(.A(new_n842), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n847), .A2(new_n466), .A3(new_n322), .ZN(new_n848));
  AOI211_X1 g647(.A(KEYINPUT59), .B(new_n466), .C1(new_n838), .C2(new_n322), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n849), .B(KEYINPUT115), .ZN(new_n850));
  XNOR2_X1  g649(.A(KEYINPUT116), .B(KEYINPUT59), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT57), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n835), .A2(KEYINPUT118), .A3(new_n786), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n567), .ZN(new_n854));
  AOI21_X1  g653(.A(KEYINPUT118), .B1(new_n835), .B2(new_n786), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n852), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n808), .A2(new_n567), .A3(new_n831), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n737), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n829), .A2(KEYINPUT117), .ZN(new_n859));
  OR2_X1    g658(.A1(new_n829), .A2(KEYINPUT117), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n851), .B1(new_n861), .B2(G148gat), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n848), .B1(new_n850), .B2(new_n862), .ZN(G1345gat));
  AOI21_X1  g662(.A(G155gat), .B1(new_n847), .B2(new_n244), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n701), .A2(G155gat), .ZN(new_n865));
  XOR2_X1   g664(.A(new_n865), .B(KEYINPUT119), .Z(new_n866));
  AOI21_X1  g665(.A(new_n864), .B1(new_n838), .B2(new_n866), .ZN(G1346gat));
  AOI22_X1  g666(.A1(new_n847), .A2(new_n299), .B1(new_n474), .B2(new_n475), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n298), .A2(new_n493), .A3(new_n492), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n868), .B1(new_n838), .B2(new_n869), .ZN(G1347gat));
  AND2_X1   g669(.A1(new_n808), .A2(new_n615), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n871), .A2(new_n459), .A3(new_n610), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n872), .A2(new_n705), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n873), .B(new_n341), .ZN(G1348gat));
  NOR2_X1   g673(.A1(new_n872), .A2(new_n737), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n875), .B1(new_n330), .B2(new_n331), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n876), .B1(new_n329), .B2(new_n875), .ZN(G1349gat));
  OAI21_X1  g676(.A(G183gat), .B1(new_n872), .B2(new_n702), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT120), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n244), .A2(new_n366), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n878), .B(new_n879), .C1(new_n872), .C2(new_n880), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(KEYINPUT60), .ZN(G1350gat));
  NAND4_X1  g681(.A1(new_n871), .A2(new_n459), .A3(new_n610), .A4(new_n299), .ZN(new_n883));
  AND3_X1   g682(.A1(new_n883), .A2(KEYINPUT121), .A3(G190gat), .ZN(new_n884));
  AOI21_X1  g683(.A(KEYINPUT121), .B1(new_n883), .B2(G190gat), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT122), .ZN(new_n886));
  OR3_X1    g685(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n886), .B1(new_n884), .B2(new_n885), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n887), .A2(new_n888), .A3(KEYINPUT61), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT61), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n886), .B(new_n890), .C1(new_n884), .C2(new_n885), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n889), .B(new_n891), .C1(G190gat), .C2(new_n883), .ZN(G1351gat));
  NOR3_X1   g691(.A1(new_n676), .A2(new_n664), .A3(new_n616), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n894), .B1(new_n856), .B2(new_n857), .ZN(new_n895));
  AND3_X1   g694(.A1(new_n895), .A2(KEYINPUT124), .A3(new_n642), .ZN(new_n896));
  AOI21_X1  g695(.A(KEYINPUT124), .B1(new_n895), .B2(new_n642), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n896), .A2(new_n897), .A3(new_n634), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n676), .A2(new_n616), .A3(new_n568), .ZN(new_n899));
  OR2_X1    g698(.A1(new_n899), .A2(KEYINPUT123), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(KEYINPUT123), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n900), .A2(new_n871), .A3(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n902), .A2(new_n634), .A3(new_n642), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(KEYINPUT125), .B1(new_n898), .B2(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(new_n897), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n895), .A2(KEYINPUT124), .A3(new_n642), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n906), .A2(G197gat), .A3(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT125), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n908), .A2(new_n909), .A3(new_n903), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n905), .A2(new_n910), .ZN(G1352gat));
  INV_X1    g710(.A(G204gat), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n902), .A2(new_n912), .A3(new_n322), .ZN(new_n913));
  XOR2_X1   g712(.A(new_n913), .B(KEYINPUT62), .Z(new_n914));
  AND2_X1   g713(.A1(new_n858), .A2(new_n893), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n914), .B1(new_n912), .B2(new_n915), .ZN(G1353gat));
  AOI21_X1  g715(.A(new_n436), .B1(new_n895), .B2(new_n244), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT63), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n902), .A2(new_n436), .A3(new_n244), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(G1354gat));
  AOI21_X1  g719(.A(G218gat), .B1(new_n902), .B2(new_n299), .ZN(new_n921));
  XOR2_X1   g720(.A(new_n895), .B(KEYINPUT126), .Z(new_n922));
  NOR2_X1   g721(.A1(new_n298), .A2(new_n437), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n923), .B(KEYINPUT127), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n921), .B1(new_n922), .B2(new_n924), .ZN(G1355gat));
endmodule


