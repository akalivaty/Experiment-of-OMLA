//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 1 0 1 1 1 0 1 0 1 0 1 0 1 0 0 1 0 0 1 0 1 1 0 0 0 0 0 0 0 1 1 1 1 1 0 0 0 0 1 0 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:18 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1294, new_n1295, new_n1296, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1371,
    new_n1372, new_n1373, new_n1374, new_n1375, new_n1376, new_n1377,
    new_n1378;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  INV_X1    g0008(.A(KEYINPUT0), .ZN(new_n209));
  INV_X1    g0009(.A(new_n201), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G50), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(new_n208), .A2(new_n209), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G87), .ZN(new_n218));
  INV_X1    g0018(.A(G250), .ZN(new_n219));
  INV_X1    g0019(.A(G97), .ZN(new_n220));
  INV_X1    g0020(.A(G257), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n206), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n216), .B1(new_n209), .B2(new_n208), .C1(new_n226), .C2(KEYINPUT1), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT2), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G226), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT64), .B(G232), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n233), .B(new_n236), .Z(G358));
  XOR2_X1   g0037(.A(G50), .B(G58), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT65), .ZN(new_n239));
  XOR2_X1   g0039(.A(G68), .B(G77), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XOR2_X1   g0042(.A(G107), .B(G116), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  INV_X1    g0045(.A(G33), .ZN(new_n246));
  INV_X1    g0046(.A(G41), .ZN(new_n247));
  OAI211_X1 g0047(.A(G1), .B(G13), .C1(new_n246), .C2(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n246), .A2(KEYINPUT3), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT3), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G33), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n249), .A2(new_n251), .A3(G1698), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(KEYINPUT66), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT3), .B(G33), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT66), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n254), .A2(new_n255), .A3(G1698), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G223), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n249), .A2(new_n251), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(G1698), .ZN(new_n260));
  AOI22_X1  g0060(.A1(new_n260), .A2(G222), .B1(G77), .B2(new_n259), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n248), .B1(new_n258), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G1), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n263), .B1(G41), .B2(G45), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G274), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n248), .A2(new_n264), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n267), .B1(new_n269), .B2(G226), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(G200), .B1(new_n262), .B2(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(G20), .A2(G33), .ZN(new_n273));
  AOI22_X1  g0073(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n214), .A2(G33), .ZN(new_n275));
  XNOR2_X1  g0075(.A(KEYINPUT8), .B(G58), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n213), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT67), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n278), .A2(KEYINPUT67), .A3(new_n213), .ZN(new_n282));
  AND2_X1   g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G13), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n284), .A2(G1), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G20), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n277), .A2(new_n283), .B1(new_n202), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n281), .A2(new_n282), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n263), .A2(G20), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n289), .A2(G50), .A3(new_n286), .A4(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n288), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT9), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G1698), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n254), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G222), .ZN(new_n297));
  INV_X1    g0097(.A(G77), .ZN(new_n298));
  OAI22_X1  g0098(.A1(new_n296), .A2(new_n297), .B1(new_n298), .B2(new_n254), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n299), .B1(G223), .B2(new_n257), .ZN(new_n300));
  OAI211_X1 g0100(.A(G190), .B(new_n270), .C1(new_n300), .C2(new_n248), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n288), .A2(KEYINPUT9), .A3(new_n291), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n272), .A2(new_n294), .A3(new_n301), .A4(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(KEYINPUT10), .ZN(new_n304));
  AND3_X1   g0104(.A1(new_n288), .A2(KEYINPUT9), .A3(new_n291), .ZN(new_n305));
  AOI21_X1  g0105(.A(KEYINPUT9), .B1(new_n288), .B2(new_n291), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT10), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n307), .A2(new_n308), .A3(new_n301), .A4(new_n272), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n304), .A2(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n262), .A2(new_n271), .ZN(new_n311));
  INV_X1    g0111(.A(G169), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G179), .ZN(new_n314));
  NOR3_X1   g0114(.A1(new_n262), .A2(new_n314), .A3(new_n271), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n292), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G200), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n318));
  INV_X1    g0118(.A(G238), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n319), .B1(new_n253), .B2(new_n256), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n254), .A2(G232), .A3(new_n295), .ZN(new_n321));
  INV_X1    g0121(.A(G107), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n321), .B1(new_n322), .B2(new_n254), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n318), .B1(new_n320), .B2(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n267), .B1(new_n269), .B2(G244), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n317), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT68), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n324), .A2(new_n325), .ZN(new_n328));
  INV_X1    g0128(.A(G190), .ZN(new_n329));
  OAI22_X1  g0129(.A1(new_n326), .A2(new_n327), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n324), .A2(KEYINPUT68), .A3(G190), .A4(new_n325), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n289), .A2(G77), .A3(new_n286), .A4(new_n290), .ZN(new_n332));
  XNOR2_X1  g0132(.A(new_n332), .B(KEYINPUT69), .ZN(new_n333));
  INV_X1    g0133(.A(new_n273), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n276), .A2(new_n334), .ZN(new_n335));
  XNOR2_X1  g0135(.A(KEYINPUT15), .B(G87), .ZN(new_n336));
  OAI22_X1  g0136(.A1(new_n336), .A2(new_n275), .B1(new_n214), .B2(new_n298), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n283), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n287), .A2(new_n298), .ZN(new_n339));
  AND2_X1   g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n330), .A2(new_n331), .A3(new_n333), .A4(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n328), .A2(G169), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n342), .B1(new_n314), .B2(new_n328), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n333), .A2(new_n339), .A3(new_n338), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AND4_X1   g0145(.A1(new_n310), .A2(new_n316), .A3(new_n341), .A4(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT75), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n347), .B1(new_n250), .B2(G33), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n246), .A2(KEYINPUT75), .A3(KEYINPUT3), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n348), .A2(new_n251), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n214), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(KEYINPUT7), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT7), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n350), .A2(new_n353), .A3(new_n214), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n352), .A2(G68), .A3(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G58), .ZN(new_n356));
  INV_X1    g0156(.A(G68), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(G20), .B1(new_n358), .B2(new_n201), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n273), .A2(G159), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n355), .A2(KEYINPUT16), .A3(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT16), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n353), .B1(new_n254), .B2(G20), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n259), .A2(KEYINPUT7), .A3(new_n214), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n357), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n364), .B1(new_n367), .B2(new_n361), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n363), .A2(new_n283), .A3(new_n368), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n283), .A2(new_n287), .ZN(new_n370));
  INV_X1    g0170(.A(new_n276), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n290), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n370), .A2(new_n373), .B1(new_n287), .B2(new_n276), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n369), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(G226), .A2(G1698), .ZN(new_n376));
  INV_X1    g0176(.A(G223), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n376), .B1(new_n377), .B2(G1698), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n378), .A2(new_n348), .A3(new_n251), .A4(new_n349), .ZN(new_n379));
  NAND2_X1  g0179(.A1(G33), .A2(G87), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n248), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(G232), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n266), .B1(new_n268), .B2(new_n382), .ZN(new_n383));
  NOR4_X1   g0183(.A1(new_n381), .A2(new_n383), .A3(KEYINPUT76), .A4(G179), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT76), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n381), .A2(new_n383), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n385), .B1(new_n386), .B2(G169), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n314), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n384), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n375), .A2(KEYINPUT18), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(KEYINPUT77), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT77), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n375), .A2(new_n392), .A3(KEYINPUT18), .A4(new_n389), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT18), .ZN(new_n394));
  INV_X1    g0194(.A(new_n374), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n357), .B1(new_n351), .B2(KEYINPUT7), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n361), .B1(new_n396), .B2(new_n354), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n289), .B1(new_n397), .B2(KEYINPUT16), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n395), .B1(new_n398), .B2(new_n368), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n387), .A2(new_n388), .ZN(new_n400));
  INV_X1    g0200(.A(new_n384), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n394), .B1(new_n399), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n391), .A2(new_n393), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n386), .A2(new_n329), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n405), .B1(G200), .B2(new_n386), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n369), .A2(new_n374), .A3(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT78), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n369), .A2(new_n406), .A3(KEYINPUT78), .A4(new_n374), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n409), .A2(KEYINPUT17), .A3(new_n410), .ZN(new_n411));
  OR2_X1    g0211(.A1(new_n407), .A2(KEYINPUT17), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n346), .A2(new_n404), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n370), .A2(G68), .A3(new_n290), .ZN(new_n415));
  XOR2_X1   g0215(.A(new_n415), .B(KEYINPUT73), .Z(new_n416));
  OAI22_X1  g0216(.A1(new_n275), .A2(new_n298), .B1(new_n214), .B2(G68), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT72), .ZN(new_n418));
  OAI22_X1  g0218(.A1(new_n417), .A2(new_n418), .B1(new_n202), .B2(new_n334), .ZN(new_n419));
  AND2_X1   g0219(.A1(new_n417), .A2(new_n418), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n283), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT11), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OR2_X1    g0223(.A1(new_n421), .A2(new_n422), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n285), .A2(G20), .A3(new_n357), .ZN(new_n425));
  XNOR2_X1  g0225(.A(new_n425), .B(KEYINPUT12), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n416), .A2(new_n423), .A3(new_n424), .A4(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT13), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n249), .A2(new_n251), .A3(G226), .A4(new_n295), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n249), .A2(new_n251), .A3(G232), .A4(G1698), .ZN(new_n431));
  NAND2_X1  g0231(.A1(G33), .A2(G97), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n318), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(KEYINPUT70), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT70), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n433), .A2(new_n436), .A3(new_n318), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n267), .B1(new_n269), .B2(G238), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n429), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  AND3_X1   g0240(.A1(new_n433), .A2(new_n436), .A3(new_n318), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n436), .B1(new_n433), .B2(new_n318), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n429), .B(new_n439), .C1(new_n441), .C2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(G169), .B1(new_n440), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(KEYINPUT14), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n444), .A2(KEYINPUT71), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n439), .B1(new_n441), .B2(new_n442), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT13), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT71), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n443), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n447), .A2(G179), .A3(new_n449), .A4(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n449), .A2(new_n443), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT14), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n453), .A2(new_n454), .A3(G169), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n446), .A2(new_n452), .A3(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT74), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n446), .A2(new_n452), .A3(KEYINPUT74), .A4(new_n455), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n428), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n447), .A2(G190), .A3(new_n449), .A4(new_n451), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n453), .A2(G200), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n428), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NOR3_X1   g0264(.A1(new_n414), .A2(new_n460), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n263), .A2(G33), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n289), .A2(new_n286), .A3(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n467), .A2(new_n322), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n285), .A2(G20), .A3(new_n322), .ZN(new_n469));
  XNOR2_X1  g0269(.A(new_n469), .B(KEYINPUT25), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g0271(.A(KEYINPUT85), .B1(new_n214), .B2(G107), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT23), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OAI211_X1 g0274(.A(KEYINPUT85), .B(KEYINPUT23), .C1(new_n214), .C2(G107), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n214), .A2(G33), .A3(G116), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n474), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n218), .A2(G20), .ZN(new_n478));
  AOI21_X1  g0278(.A(KEYINPUT22), .B1(new_n254), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  AND3_X1   g0280(.A1(new_n348), .A2(new_n251), .A3(new_n349), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n481), .A2(KEYINPUT22), .A3(new_n214), .A4(G87), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n480), .A2(new_n482), .A3(KEYINPUT24), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n283), .ZN(new_n484));
  AOI21_X1  g0284(.A(KEYINPUT24), .B1(new_n480), .B2(new_n482), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n471), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n263), .A2(G45), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT5), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n247), .ZN(new_n489));
  NAND2_X1  g0289(.A1(KEYINPUT5), .A2(G41), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n487), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n491), .A2(new_n318), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(G264), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n491), .A2(G274), .ZN(new_n494));
  NAND2_X1  g0294(.A1(G257), .A2(G1698), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n495), .B1(new_n219), .B2(G1698), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n496), .A2(new_n348), .A3(new_n251), .A4(new_n349), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT86), .ZN(new_n498));
  NAND2_X1  g0298(.A1(G33), .A2(G294), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n318), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n498), .B1(new_n497), .B2(new_n499), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n493), .B(new_n494), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n317), .ZN(new_n504));
  OR2_X1    g0304(.A1(new_n501), .A2(new_n502), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n505), .A2(new_n329), .A3(new_n493), .A4(new_n494), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n486), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n503), .A2(new_n314), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(KEYINPUT87), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT87), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n510), .B1(new_n503), .B2(G169), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n509), .B1(new_n508), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n507), .B1(new_n512), .B2(new_n486), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT82), .ZN(new_n514));
  INV_X1    g0314(.A(new_n467), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(G87), .ZN(new_n516));
  AOI21_X1  g0316(.A(KEYINPUT75), .B1(new_n246), .B2(KEYINPUT3), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n246), .A2(KEYINPUT3), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n519), .A2(new_n214), .A3(G68), .A4(new_n349), .ZN(new_n520));
  NOR2_X1   g0320(.A1(G87), .A2(G97), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n521), .A2(new_n322), .B1(new_n432), .B2(new_n214), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT19), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n214), .ZN(new_n524));
  OAI22_X1  g0324(.A1(new_n522), .A2(new_n523), .B1(new_n432), .B2(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n289), .B1(new_n520), .B2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT81), .ZN(new_n527));
  INV_X1    g0327(.A(new_n336), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n528), .A2(new_n286), .ZN(new_n529));
  NOR3_X1   g0329(.A1(new_n526), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n348), .A2(new_n349), .A3(new_n214), .A4(new_n251), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n531), .A2(new_n357), .ZN(new_n532));
  NOR3_X1   g0332(.A1(new_n432), .A2(KEYINPUT19), .A3(G20), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n218), .A2(new_n220), .A3(new_n322), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n432), .A2(new_n214), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n533), .B1(new_n536), .B2(KEYINPUT19), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n283), .B1(new_n532), .B2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n529), .ZN(new_n539));
  AOI21_X1  g0339(.A(KEYINPUT81), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n516), .B1(new_n530), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n319), .A2(G1698), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n348), .A2(new_n349), .A3(new_n542), .A4(new_n251), .ZN(new_n543));
  NAND2_X1  g0343(.A1(G33), .A2(G116), .ZN(new_n544));
  AND2_X1   g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT80), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n519), .A2(G244), .A3(G1698), .A4(new_n349), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n348), .A2(new_n349), .A3(G244), .A4(new_n251), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n544), .B(new_n543), .C1(new_n549), .C2(new_n295), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(KEYINPUT80), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n548), .A2(new_n551), .A3(new_n318), .ZN(new_n552));
  INV_X1    g0352(.A(G45), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n553), .A2(G1), .ZN(new_n554));
  AND2_X1   g0354(.A1(new_n554), .A2(G274), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n554), .A2(new_n219), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n248), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n317), .B1(new_n552), .B2(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n514), .B1(new_n541), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n527), .B1(new_n526), .B2(new_n529), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n538), .A2(KEYINPUT81), .A3(new_n539), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n560), .A2(new_n561), .B1(G87), .B2(new_n515), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n318), .B1(new_n550), .B2(KEYINPUT80), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n546), .B1(new_n545), .B2(new_n547), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n557), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(G200), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n562), .A2(new_n566), .A3(KEYINPUT82), .ZN(new_n567));
  OAI211_X1 g0367(.A(G190), .B(new_n557), .C1(new_n563), .C2(new_n564), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n559), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  OAI22_X1  g0369(.A1(new_n530), .A2(new_n540), .B1(new_n336), .B2(new_n467), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n314), .B(new_n557), .C1(new_n563), .C2(new_n564), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n565), .A2(new_n312), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  AND2_X1   g0373(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT6), .ZN(new_n575));
  NOR3_X1   g0375(.A1(new_n575), .A2(new_n220), .A3(G107), .ZN(new_n576));
  XNOR2_X1  g0376(.A(G97), .B(G107), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n576), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  OAI22_X1  g0378(.A1(new_n578), .A2(new_n214), .B1(new_n298), .B2(new_n334), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n322), .B1(new_n365), .B2(new_n366), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n283), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n515), .A2(G97), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n286), .A2(G97), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n581), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n249), .A2(new_n251), .A3(G250), .A4(G1698), .ZN(new_n586));
  AND2_X1   g0386(.A1(KEYINPUT4), .A2(G244), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n249), .A2(new_n251), .A3(new_n587), .A4(new_n295), .ZN(new_n588));
  NAND2_X1  g0388(.A1(G33), .A2(G283), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n586), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT4), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n591), .B1(new_n549), .B2(G1698), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n318), .ZN(new_n594));
  INV_X1    g0394(.A(new_n490), .ZN(new_n595));
  NOR2_X1   g0395(.A1(KEYINPUT5), .A2(G41), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n554), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n248), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n494), .B1(new_n598), .B2(new_n221), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n312), .B1(new_n594), .B2(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n248), .B1(new_n590), .B2(new_n592), .ZN(new_n602));
  NOR3_X1   g0402(.A1(new_n602), .A2(new_n314), .A3(new_n599), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n585), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(KEYINPUT79), .ZN(new_n605));
  INV_X1    g0405(.A(new_n585), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n594), .A2(new_n600), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n607), .A2(G190), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n602), .A2(new_n599), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n609), .A2(G200), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n606), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT79), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n585), .B(new_n612), .C1(new_n601), .C2(new_n603), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n605), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(G116), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n278), .A2(new_n213), .B1(G20), .B2(new_n615), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n589), .B(new_n214), .C1(G33), .C2(new_n220), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n616), .A2(KEYINPUT20), .A3(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT83), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n616), .A2(KEYINPUT83), .A3(new_n617), .A4(KEYINPUT20), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n616), .A2(new_n617), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT20), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n620), .A2(new_n621), .A3(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n289), .A2(G116), .A3(new_n286), .A4(new_n466), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n287), .A2(new_n615), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n492), .A2(G270), .B1(G274), .B2(new_n491), .ZN(new_n629));
  NAND2_X1  g0429(.A1(G264), .A2(G1698), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n630), .B1(new_n221), .B2(G1698), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n631), .A2(new_n348), .A3(new_n251), .A4(new_n349), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n259), .A2(G303), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n318), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n629), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n628), .A2(G169), .A3(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT21), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n629), .A2(G179), .A3(new_n635), .ZN(new_n639));
  INV_X1    g0439(.A(G270), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n494), .B1(new_n598), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n248), .B1(new_n632), .B2(new_n633), .ZN(new_n642));
  OAI211_X1 g0442(.A(KEYINPUT21), .B(G169), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  AOI22_X1  g0444(.A1(new_n637), .A2(new_n638), .B1(new_n644), .B2(new_n628), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT84), .ZN(new_n646));
  AOI21_X1  g0446(.A(G200), .B1(new_n629), .B2(new_n635), .ZN(new_n647));
  NOR3_X1   g0447(.A1(new_n641), .A2(new_n642), .A3(G190), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n646), .B1(new_n649), .B2(new_n628), .ZN(new_n650));
  INV_X1    g0450(.A(new_n628), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n651), .B(KEYINPUT84), .C1(new_n648), .C2(new_n647), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n645), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n614), .A2(new_n653), .ZN(new_n654));
  AND4_X1   g0454(.A1(new_n465), .A2(new_n513), .A3(new_n574), .A4(new_n654), .ZN(G372));
  INV_X1    g0455(.A(new_n316), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n454), .B1(new_n453), .B2(G169), .ZN(new_n657));
  AOI211_X1 g0457(.A(KEYINPUT14), .B(new_n312), .C1(new_n449), .C2(new_n443), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(KEYINPUT74), .B1(new_n659), .B2(new_n452), .ZN(new_n660));
  INV_X1    g0460(.A(new_n459), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n427), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n662), .B1(new_n464), .B2(new_n345), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(new_n413), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n403), .A2(new_n390), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n656), .B1(new_n666), .B2(new_n310), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n404), .A2(new_n413), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n662), .A2(new_n669), .A3(new_n463), .A4(new_n346), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n605), .A2(new_n613), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n569), .A2(new_n671), .A3(new_n573), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(KEYINPUT26), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n605), .A2(new_n613), .A3(new_n611), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n560), .A2(new_n561), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n675), .A2(new_n568), .A3(new_n516), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT88), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n677), .B1(new_n565), .B2(G200), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n558), .A2(new_n677), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n507), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NOR3_X1   g0481(.A1(new_n503), .A2(new_n510), .A3(new_n314), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n503), .A2(G169), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(KEYINPUT87), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n503), .A2(new_n314), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n682), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n486), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n645), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n674), .A2(new_n681), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n571), .ZN(new_n690));
  AOI21_X1  g0490(.A(G169), .B1(new_n552), .B2(new_n557), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AOI22_X1  g0492(.A1(new_n679), .A2(new_n680), .B1(new_n570), .B2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT26), .ZN(new_n694));
  INV_X1    g0494(.A(new_n604), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n673), .A2(new_n573), .A3(new_n689), .A4(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n667), .B1(new_n670), .B2(new_n698), .ZN(G369));
  AND2_X1   g0499(.A1(new_n653), .A2(KEYINPUT89), .ZN(new_n700));
  INV_X1    g0500(.A(new_n285), .ZN(new_n701));
  OR3_X1    g0501(.A1(new_n701), .A2(KEYINPUT27), .A3(G20), .ZN(new_n702));
  OAI21_X1  g0502(.A(KEYINPUT27), .B1(new_n701), .B2(G20), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n702), .A2(G213), .A3(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(G343), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n628), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n707), .B1(new_n653), .B2(KEYINPUT89), .ZN(new_n708));
  OAI22_X1  g0508(.A1(new_n700), .A2(new_n708), .B1(new_n645), .B2(new_n707), .ZN(new_n709));
  XOR2_X1   g0509(.A(new_n709), .B(KEYINPUT90), .Z(new_n710));
  AND2_X1   g0510(.A1(new_n710), .A2(G330), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n512), .A2(new_n486), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n506), .A2(new_n504), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n687), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n486), .A2(new_n706), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n712), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT91), .ZN(new_n717));
  XNOR2_X1  g0517(.A(new_n716), .B(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n706), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n712), .A2(new_n719), .ZN(new_n720));
  OR2_X1    g0520(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n711), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n512), .A2(new_n486), .A3(new_n719), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n645), .A2(new_n706), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n718), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n722), .A2(new_n723), .A3(new_n725), .ZN(G399));
  INV_X1    g0526(.A(new_n207), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(G41), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(G1), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n521), .A2(new_n322), .A3(new_n615), .ZN(new_n731));
  OAI22_X1  g0531(.A1(new_n730), .A2(new_n731), .B1(new_n211), .B2(new_n729), .ZN(new_n732));
  XOR2_X1   g0532(.A(KEYINPUT92), .B(KEYINPUT28), .Z(new_n733));
  XNOR2_X1  g0533(.A(new_n732), .B(new_n733), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n574), .A2(new_n654), .A3(new_n513), .A4(new_n719), .ZN(new_n735));
  NOR3_X1   g0535(.A1(new_n641), .A2(new_n642), .A3(new_n314), .ZN(new_n736));
  AND3_X1   g0536(.A1(new_n505), .A2(new_n493), .A3(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n565), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT93), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(KEYINPUT30), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n737), .A2(new_n738), .A3(new_n609), .A4(new_n740), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n609), .A2(new_n505), .A3(new_n493), .A4(new_n736), .ZN(new_n742));
  OAI22_X1  g0542(.A1(new_n742), .A2(new_n565), .B1(new_n739), .B2(KEYINPUT30), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  AND3_X1   g0544(.A1(new_n565), .A2(new_n314), .A3(new_n636), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT94), .ZN(new_n746));
  AND3_X1   g0546(.A1(new_n607), .A2(new_n746), .A3(new_n503), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n746), .B1(new_n607), .B2(new_n503), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n745), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n719), .B1(new_n744), .B2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT31), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n735), .A2(new_n752), .ZN(new_n753));
  AOI211_X1 g0553(.A(KEYINPUT31), .B(new_n719), .C1(new_n744), .C2(new_n749), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n753), .A2(G330), .A3(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n672), .A2(new_n694), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT95), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n693), .A2(new_n759), .A3(KEYINPUT26), .A4(new_n695), .ZN(new_n760));
  OAI211_X1 g0560(.A(new_n562), .B(new_n568), .C1(new_n558), .C2(new_n677), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n566), .A2(KEYINPUT88), .ZN(new_n762));
  OAI211_X1 g0562(.A(new_n573), .B(new_n695), .C1(new_n761), .C2(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(KEYINPUT95), .B1(new_n763), .B2(new_n694), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n758), .A2(new_n760), .A3(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n714), .B1(new_n761), .B2(new_n762), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n614), .ZN(new_n767));
  AOI22_X1  g0567(.A1(new_n767), .A2(new_n688), .B1(new_n570), .B2(new_n692), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n769), .A2(KEYINPUT29), .A3(new_n719), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(KEYINPUT96), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n706), .B1(new_n765), .B2(new_n768), .ZN(new_n772));
  INV_X1    g0572(.A(KEYINPUT96), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n772), .A2(new_n773), .A3(KEYINPUT29), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n771), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n697), .A2(new_n719), .ZN(new_n776));
  INV_X1    g0576(.A(KEYINPUT29), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n757), .B1(new_n775), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n734), .B1(new_n779), .B2(G1), .ZN(G364));
  NOR2_X1   g0580(.A1(new_n284), .A2(G20), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G45), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n729), .A2(G1), .A3(new_n782), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT97), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n711), .A2(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n785), .B1(G330), .B2(new_n710), .ZN(new_n786));
  INV_X1    g0586(.A(new_n784), .ZN(new_n787));
  OAI211_X1 g0587(.A(G1), .B(G13), .C1(new_n214), .C2(G169), .ZN(new_n788));
  OR2_X1    g0588(.A1(new_n788), .A2(KEYINPUT98), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(KEYINPUT98), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n329), .A2(G20), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  OR2_X1    g0594(.A1(new_n794), .A2(KEYINPUT100), .ZN(new_n795));
  NOR2_X1   g0595(.A1(G179), .A2(G200), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n794), .A2(KEYINPUT100), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(G159), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n800), .B(KEYINPUT32), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n214), .A2(new_n329), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n314), .A2(G200), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n317), .A2(G179), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n804), .A2(new_n356), .B1(new_n806), .B2(new_n218), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n214), .B1(new_n796), .B2(G190), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n314), .A2(new_n317), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n794), .A2(new_n809), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n254), .B1(new_n808), .B2(new_n220), .C1(new_n810), .C2(new_n357), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n809), .A2(new_n802), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n807), .B(new_n811), .C1(G50), .C2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n794), .A2(new_n803), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT99), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n815), .A2(new_n816), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n795), .A2(new_n797), .A3(new_n805), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n821), .A2(G77), .B1(G107), .B2(new_n823), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n801), .A2(new_n814), .A3(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n798), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n821), .A2(G311), .B1(new_n826), .B2(G329), .ZN(new_n827));
  INV_X1    g0627(.A(G322), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n259), .B1(new_n804), .B2(new_n828), .ZN(new_n829));
  XOR2_X1   g0629(.A(KEYINPUT33), .B(G317), .Z(new_n830));
  INV_X1    g0630(.A(G326), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n810), .A2(new_n830), .B1(new_n812), .B2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n808), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n829), .B(new_n832), .C1(G294), .C2(new_n833), .ZN(new_n834));
  XOR2_X1   g0634(.A(new_n806), .B(KEYINPUT101), .Z(new_n835));
  AOI22_X1  g0635(.A1(G303), .A2(new_n835), .B1(new_n823), .B2(G283), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n827), .A2(new_n834), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n792), .B1(new_n825), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(G13), .A2(G33), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n840), .A2(G20), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n791), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n481), .A2(new_n727), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n241), .A2(new_n553), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n212), .A2(G45), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n843), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n727), .A2(new_n259), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n847), .A2(G355), .B1(new_n615), .B2(new_n727), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  AOI211_X1 g0649(.A(new_n787), .B(new_n838), .C1(new_n842), .C2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n841), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n850), .B1(new_n710), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n786), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g0653(.A(new_n853), .B(KEYINPUT102), .ZN(G396));
  NAND2_X1  g0654(.A1(new_n344), .A2(new_n706), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n341), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n345), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n345), .A2(new_n706), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n776), .B(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n784), .B1(new_n862), .B2(new_n757), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n863), .B1(new_n757), .B2(new_n862), .ZN(new_n864));
  INV_X1    g0664(.A(new_n810), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n865), .A2(G150), .B1(new_n813), .B2(G137), .ZN(new_n866));
  XNOR2_X1  g0666(.A(KEYINPUT103), .B(G143), .ZN(new_n867));
  OAI221_X1 g0667(.A(new_n866), .B1(new_n804), .B2(new_n867), .C1(new_n820), .C2(new_n799), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n868), .B(KEYINPUT34), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n481), .B1(new_n356), .B2(new_n808), .ZN(new_n870));
  INV_X1    g0670(.A(new_n835), .ZN(new_n871));
  OAI22_X1  g0671(.A1(new_n871), .A2(new_n202), .B1(new_n357), .B2(new_n822), .ZN(new_n872));
  AOI211_X1 g0672(.A(new_n870), .B(new_n872), .C1(G132), .C2(new_n826), .ZN(new_n873));
  INV_X1    g0673(.A(G283), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n259), .B1(new_n810), .B2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(G303), .ZN(new_n876));
  INV_X1    g0676(.A(G294), .ZN(new_n877));
  OAI22_X1  g0677(.A1(new_n812), .A2(new_n876), .B1(new_n804), .B2(new_n877), .ZN(new_n878));
  AOI211_X1 g0678(.A(new_n875), .B(new_n878), .C1(G97), .C2(new_n833), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n821), .A2(G116), .B1(new_n826), .B2(G311), .ZN(new_n880));
  AOI22_X1  g0680(.A1(G107), .A2(new_n835), .B1(new_n823), .B2(G87), .ZN(new_n881));
  AND2_X1   g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AOI22_X1  g0682(.A1(new_n869), .A2(new_n873), .B1(new_n879), .B2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT104), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n792), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n885), .B1(new_n884), .B2(new_n883), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n792), .A2(new_n840), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n886), .B(new_n784), .C1(G77), .C2(new_n887), .ZN(new_n888));
  XOR2_X1   g0688(.A(new_n888), .B(KEYINPUT105), .Z(new_n889));
  NOR2_X1   g0689(.A1(new_n861), .A2(new_n840), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n864), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n891), .B(KEYINPUT106), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(G384));
  NAND2_X1  g0693(.A1(new_n215), .A2(G116), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT35), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n894), .B1(new_n578), .B2(new_n895), .ZN(new_n896));
  OAI22_X1  g0696(.A1(new_n896), .A2(KEYINPUT107), .B1(new_n895), .B2(new_n578), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n897), .B1(KEYINPUT107), .B2(new_n896), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n898), .B(KEYINPUT36), .ZN(new_n899));
  OR3_X1    g0699(.A1(new_n211), .A2(new_n298), .A3(new_n358), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n202), .A2(G68), .ZN(new_n901));
  AOI211_X1 g0701(.A(new_n263), .B(G13), .C1(new_n900), .C2(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n763), .A2(KEYINPUT26), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n904), .B1(KEYINPUT26), .B2(new_n672), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n706), .B1(new_n905), .B2(new_n768), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n465), .B1(new_n906), .B2(KEYINPUT29), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n774), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n773), .B1(new_n772), .B2(KEYINPUT29), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n667), .ZN(new_n912));
  INV_X1    g0712(.A(new_n704), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n665), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n697), .A2(new_n719), .A3(new_n861), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n858), .B(KEYINPUT108), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n427), .A2(new_n706), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n662), .A2(new_n463), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n458), .A2(new_n459), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n427), .B(new_n706), .C1(new_n919), .C2(new_n464), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n915), .A2(new_n916), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n363), .A2(new_n283), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n397), .A2(KEYINPUT16), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n913), .B1(new_n924), .B2(new_n395), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n668), .A2(new_n926), .ZN(new_n927));
  OAI22_X1  g0727(.A1(new_n924), .A2(new_n395), .B1(new_n389), .B2(new_n913), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n928), .A2(new_n409), .A3(new_n410), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(KEYINPUT37), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT37), .B1(new_n375), .B2(new_n389), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n375), .A2(new_n913), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n931), .A2(new_n409), .A3(new_n410), .A4(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n927), .A2(KEYINPUT38), .A3(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT38), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n925), .B1(new_n404), .B2(new_n413), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n409), .A2(new_n410), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n931), .A2(new_n932), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n938), .A2(new_n939), .B1(new_n929), .B2(KEYINPUT37), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n936), .B1(new_n937), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n935), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n914), .B1(new_n921), .B2(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n662), .A2(new_n706), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT109), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n407), .B1(new_n399), .B2(new_n402), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n399), .A2(new_n704), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n945), .B(KEYINPUT37), .C1(new_n946), .C2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n933), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n932), .B(new_n407), .C1(new_n399), .C2(new_n402), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n945), .B1(new_n950), .B2(KEYINPUT37), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n411), .A2(new_n412), .B1(new_n390), .B2(new_n403), .ZN(new_n952));
  OAI22_X1  g0752(.A1(new_n949), .A2(new_n951), .B1(new_n952), .B2(new_n932), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n936), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT39), .ZN(new_n955));
  AND3_X1   g0755(.A1(new_n954), .A2(new_n935), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n955), .B1(new_n935), .B2(new_n941), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n944), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n943), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n912), .B(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n918), .A2(new_n920), .ZN(new_n961));
  AOI211_X1 g0761(.A(new_n860), .B(new_n754), .C1(new_n735), .C2(new_n752), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n954), .A2(new_n935), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(KEYINPUT40), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n753), .A2(new_n755), .A3(new_n861), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n967), .B1(new_n918), .B2(new_n920), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT40), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n968), .A2(new_n969), .A3(new_n942), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n966), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n753), .A2(new_n755), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n972), .A2(new_n670), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n971), .B(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(G330), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n960), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n263), .B2(new_n781), .ZN(new_n977));
  NOR3_X1   g0777(.A1(new_n960), .A2(new_n974), .A3(new_n975), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n903), .B1(new_n977), .B2(new_n978), .ZN(G367));
  NOR2_X1   g0779(.A1(new_n562), .A2(new_n719), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n693), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(new_n573), .B2(new_n980), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n982), .B(KEYINPUT43), .Z(new_n983));
  INV_X1    g0783(.A(KEYINPUT110), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n674), .B1(new_n606), .B2(new_n719), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n725), .A2(new_n985), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT42), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n695), .A2(new_n706), .ZN(new_n988));
  AND2_X1   g0788(.A1(new_n985), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n989), .A2(new_n712), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n719), .B1(new_n990), .B2(new_n671), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n984), .B1(new_n987), .B2(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n986), .A2(KEYINPUT42), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT42), .ZN(new_n994));
  NOR3_X1   g0794(.A1(new_n725), .A2(new_n994), .A3(new_n985), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n991), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n996), .A2(KEYINPUT110), .ZN(new_n997));
  OAI211_X1 g0797(.A(KEYINPUT111), .B(new_n983), .C1(new_n992), .C2(new_n997), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n987), .A2(new_n984), .A3(new_n991), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n996), .A2(KEYINPUT110), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n998), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n999), .A2(new_n1000), .ZN(new_n1004));
  AOI21_X1  g0804(.A(KEYINPUT111), .B1(new_n1004), .B2(new_n983), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n1003), .A2(new_n1005), .B1(new_n722), .B2(new_n989), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1004), .A2(new_n983), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT111), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n722), .A2(new_n989), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n1009), .A2(new_n1010), .A3(new_n998), .A4(new_n1002), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n728), .B(KEYINPUT41), .Z(new_n1012));
  OAI21_X1  g0812(.A(new_n725), .B1(new_n721), .B2(new_n724), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n711), .B(new_n1013), .ZN(new_n1014));
  AND2_X1   g0814(.A1(new_n1014), .A2(new_n779), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n725), .A2(new_n723), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n989), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT113), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT44), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n1016), .B(new_n989), .C1(new_n1018), .C2(new_n1019), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n1016), .A2(new_n989), .ZN(new_n1026));
  XOR2_X1   g0826(.A(KEYINPUT112), .B(KEYINPUT45), .Z(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1026), .B(new_n1028), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1025), .A2(new_n1029), .A3(new_n722), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n722), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1026), .B(new_n1027), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n1021), .A2(new_n1022), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1031), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1015), .A2(new_n1030), .A3(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1012), .B1(new_n1035), .B2(new_n779), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n782), .A2(G1), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1006), .B(new_n1011), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n842), .B1(new_n207), .B2(new_n336), .ZN(new_n1039));
  AND2_X1   g0839(.A1(new_n236), .A2(new_n843), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n784), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(G317), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n798), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT46), .ZN(new_n1044));
  NOR3_X1   g0844(.A1(new_n871), .A2(new_n1044), .A3(new_n615), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n1043), .B(new_n1045), .C1(G97), .C2(new_n823), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1044), .B1(new_n806), .B2(new_n615), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1047), .B(new_n350), .C1(new_n322), .C2(new_n808), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n804), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n865), .A2(G294), .B1(new_n1049), .B2(G303), .ZN(new_n1050));
  INV_X1    g0850(.A(G311), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1050), .B1(new_n1051), .B2(new_n812), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n1048), .B(new_n1052), .C1(G283), .C2(new_n821), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n254), .B1(new_n806), .B2(new_n356), .C1(new_n810), .C2(new_n799), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n820), .A2(new_n202), .B1(new_n298), .B2(new_n822), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n1054), .B(new_n1055), .C1(G137), .C2(new_n826), .ZN(new_n1056));
  INV_X1    g0856(.A(G150), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n812), .A2(new_n867), .B1(new_n804), .B2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n808), .A2(new_n357), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT114), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n1046), .A2(new_n1053), .B1(new_n1056), .B2(new_n1061), .ZN(new_n1062));
  OR2_X1    g0862(.A1(new_n1062), .A2(KEYINPUT47), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n792), .B1(new_n1062), .B2(KEYINPUT47), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1041), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n982), .B2(new_n851), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1038), .A2(new_n1066), .ZN(G387));
  NOR2_X1   g0867(.A1(new_n1015), .A2(new_n729), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n779), .B2(new_n1014), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1014), .A2(new_n1037), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n847), .A2(new_n731), .B1(new_n322), .B2(new_n727), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n233), .A2(new_n553), .ZN(new_n1072));
  AOI211_X1 g0872(.A(G45), .B(new_n731), .C1(G68), .C2(G77), .ZN(new_n1073));
  AND3_X1   g0873(.A1(new_n371), .A2(KEYINPUT50), .A3(new_n202), .ZN(new_n1074));
  AOI21_X1  g0874(.A(KEYINPUT50), .B1(new_n371), .B2(new_n202), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1073), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n843), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1071), .B1(new_n1072), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n787), .B1(new_n1078), .B2(new_n842), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(G322), .A2(new_n813), .B1(new_n1049), .B2(G317), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n1080), .B1(new_n1051), .B2(new_n810), .C1(new_n820), .C2(new_n876), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  OR2_X1    g0882(.A1(new_n1082), .A2(KEYINPUT48), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1082), .A2(KEYINPUT48), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n806), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n1085), .A2(G294), .B1(new_n833), .B2(G283), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1083), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  OR2_X1    g0888(.A1(new_n1088), .A2(KEYINPUT49), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n350), .B1(new_n798), .B2(new_n831), .C1(new_n615), .C2(new_n822), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(new_n1088), .B2(KEYINPUT49), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n820), .A2(new_n357), .B1(new_n276), .B2(new_n810), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT115), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(G97), .A2(new_n823), .B1(new_n826), .B2(G150), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n806), .A2(new_n298), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n804), .A2(new_n202), .ZN(new_n1096));
  AOI211_X1 g0896(.A(new_n1095), .B(new_n1096), .C1(G159), .C2(new_n813), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n833), .A2(new_n528), .ZN(new_n1098));
  AND4_X1   g0898(.A1(new_n481), .A2(new_n1094), .A3(new_n1097), .A4(new_n1098), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n1089), .A2(new_n1091), .B1(new_n1093), .B2(new_n1099), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n1079), .B1(new_n792), .B2(new_n1100), .C1(new_n721), .C2(new_n851), .ZN(new_n1101));
  AND2_X1   g0901(.A1(new_n1070), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1069), .A2(new_n1102), .ZN(G393));
  NAND2_X1  g0903(.A1(new_n1034), .A2(new_n1030), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT117), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1014), .A2(new_n779), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  AND2_X1   g0907(.A1(new_n1107), .A2(new_n728), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1035), .A2(new_n1105), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1104), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n989), .A2(new_n841), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n842), .B1(new_n220), .B2(new_n207), .ZN(new_n1115));
  AND2_X1   g0915(.A1(new_n244), .A2(new_n843), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n784), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(G150), .A2(new_n813), .B1(new_n1049), .B2(G159), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1118), .A2(KEYINPUT51), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(G87), .B2(new_n823), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n821), .A2(new_n371), .B1(KEYINPUT51), .B2(new_n1118), .ZN(new_n1121));
  OR2_X1    g0921(.A1(new_n798), .A2(new_n867), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n810), .A2(new_n202), .B1(new_n806), .B2(new_n357), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n350), .B(new_n1123), .C1(G77), .C2(new_n833), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .A4(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n254), .B1(new_n1085), .B2(G283), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n1126), .B1(new_n798), .B2(new_n828), .C1(new_n322), .C2(new_n822), .ZN(new_n1127));
  XOR2_X1   g0927(.A(new_n1127), .B(KEYINPUT116), .Z(new_n1128));
  OAI22_X1  g0928(.A1(new_n812), .A2(new_n1042), .B1(new_n804), .B2(new_n1051), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1129), .B(KEYINPUT52), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n865), .A2(G303), .B1(G116), .B2(new_n833), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n1130), .B(new_n1131), .C1(new_n877), .C2(new_n820), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1125), .B1(new_n1128), .B2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1117), .B1(new_n1133), .B2(new_n791), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n1113), .A2(new_n1037), .B1(new_n1114), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1112), .A2(new_n1135), .ZN(G390));
  OAI21_X1  g0936(.A(new_n784), .B1(new_n887), .B2(new_n371), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(KEYINPUT54), .B(G143), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n821), .A2(new_n1139), .B1(G50), .B2(new_n823), .ZN(new_n1140));
  INV_X1    g0940(.A(G132), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n254), .B1(new_n804), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(G137), .ZN(new_n1143));
  INV_X1    g0943(.A(G128), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n810), .A2(new_n1143), .B1(new_n812), .B2(new_n1144), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n1142), .B(new_n1145), .C1(G159), .C2(new_n833), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT53), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1147), .B1(new_n806), .B2(new_n1057), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1085), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n826), .A2(G125), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1140), .A2(new_n1146), .A3(new_n1150), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n357), .A2(new_n822), .B1(new_n798), .B2(new_n877), .ZN(new_n1152));
  XOR2_X1   g0952(.A(new_n1152), .B(KEYINPUT118), .Z(new_n1153));
  AOI22_X1  g0953(.A1(new_n821), .A2(G97), .B1(G87), .B2(new_n835), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n812), .A2(new_n874), .B1(new_n804), .B2(new_n615), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n254), .B(new_n1155), .C1(G107), .C2(new_n865), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1154), .B(new_n1156), .C1(new_n298), .C2(new_n808), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1151), .B1(new_n1153), .B2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1137), .B1(new_n1158), .B2(new_n791), .ZN(new_n1159));
  AOI21_X1  g0959(.A(KEYINPUT38), .B1(new_n927), .B2(new_n934), .ZN(new_n1160));
  NOR3_X1   g0960(.A1(new_n937), .A2(new_n940), .A3(new_n936), .ZN(new_n1161));
  OAI21_X1  g0961(.A(KEYINPUT39), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n954), .A2(new_n935), .A3(new_n955), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1159), .B1(new_n1164), .B2(new_n840), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n915), .A2(new_n916), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n944), .B1(new_n1166), .B2(new_n961), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n769), .A2(new_n719), .A3(new_n857), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n1168), .A2(new_n859), .B1(new_n918), .B2(new_n920), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n944), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n964), .A2(new_n1170), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n1167), .A2(new_n1164), .B1(new_n1169), .B2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n961), .A2(new_n962), .A3(G330), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1162), .B(new_n1163), .C1(new_n921), .C2(new_n944), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n858), .B1(new_n772), .B2(new_n857), .ZN(new_n1177));
  AND2_X1   g0977(.A1(new_n918), .A2(new_n920), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1170), .B(new_n964), .C1(new_n1177), .C2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1176), .A2(new_n1179), .A3(new_n1173), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1175), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1037), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1165), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1168), .A2(new_n859), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n753), .A2(G330), .A3(new_n755), .A4(new_n861), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1185), .A2(new_n918), .A3(new_n920), .ZN(new_n1186));
  AND3_X1   g0986(.A1(new_n1173), .A2(new_n1184), .A3(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1166), .B1(new_n1173), .B2(new_n1186), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n907), .B1(new_n771), .B2(new_n774), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n663), .A2(new_n413), .B1(new_n390), .B2(new_n403), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n310), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n316), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n972), .A2(new_n670), .A3(new_n975), .ZN(new_n1194));
  NOR3_X1   g0994(.A1(new_n1190), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1189), .A2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n729), .B1(new_n1181), .B2(new_n1196), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1175), .A2(new_n1195), .A3(new_n1189), .A4(new_n1180), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1183), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(G378));
  NAND2_X1  g1000(.A1(new_n1198), .A2(new_n1195), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT57), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n975), .B1(new_n966), .B2(new_n970), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1166), .A2(new_n942), .A3(new_n961), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n914), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1170), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n310), .A2(new_n316), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(KEYINPUT119), .B(KEYINPUT56), .ZN(new_n1209));
  AND2_X1   g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n292), .A2(new_n913), .ZN(new_n1212));
  XOR2_X1   g1012(.A(new_n1212), .B(KEYINPUT55), .Z(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  OR3_X1    g1014(.A1(new_n1210), .A2(new_n1211), .A3(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1214), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  NOR3_X1   g1017(.A1(new_n1206), .A2(new_n1207), .A3(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1217), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(new_n943), .B2(new_n958), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1203), .B1(new_n1218), .B2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n969), .B1(new_n968), .B2(new_n964), .ZN(new_n1222));
  AND4_X1   g1022(.A1(new_n969), .A2(new_n942), .A3(new_n961), .A4(new_n962), .ZN(new_n1223));
  OAI21_X1  g1023(.A(G330), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1217), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n943), .A2(new_n958), .A3(new_n1219), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1221), .A2(new_n1227), .ZN(new_n1228));
  AND3_X1   g1028(.A1(new_n1201), .A2(new_n1202), .A3(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1202), .B1(new_n1201), .B2(new_n1228), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n728), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1219), .A2(new_n839), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n784), .B1(new_n887), .B2(G50), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n821), .A2(new_n528), .B1(G58), .B2(new_n823), .ZN(new_n1234));
  NOR4_X1   g1034(.A1(new_n1095), .A2(new_n1059), .A3(new_n481), .A4(G41), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n812), .A2(new_n615), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n810), .A2(new_n220), .B1(new_n804), .B2(new_n322), .ZN(new_n1237));
  AOI211_X1 g1037(.A(new_n1236), .B(new_n1237), .C1(new_n826), .C2(G283), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1234), .A2(new_n1235), .A3(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT58), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n247), .B1(new_n350), .B2(new_n246), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n1239), .A2(new_n1240), .B1(new_n202), .B2(new_n1241), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n804), .A2(new_n1144), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n810), .A2(new_n1141), .B1(new_n806), .B2(new_n1138), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n1243), .B(new_n1244), .C1(G125), .C2(new_n813), .ZN(new_n1245));
  OAI221_X1 g1045(.A(new_n1245), .B1(new_n1143), .B2(new_n820), .C1(new_n1057), .C2(new_n808), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(KEYINPUT59), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n246), .B(new_n247), .C1(new_n822), .C2(new_n799), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1248), .B1(G124), .B2(new_n826), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1247), .A2(new_n1249), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1246), .A2(KEYINPUT59), .ZN(new_n1251));
  OAI221_X1 g1051(.A(new_n1242), .B1(new_n1240), .B2(new_n1239), .C1(new_n1250), .C2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1233), .B1(new_n1252), .B2(new_n791), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1232), .A2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1255), .B1(new_n1228), .B2(new_n1037), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1231), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT120), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(new_n1257), .B(new_n1258), .ZN(G375));
  OAI21_X1  g1059(.A(KEYINPUT121), .B1(new_n1189), .B2(new_n1195), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1012), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1173), .A2(new_n1184), .A3(new_n1186), .ZN(new_n1262));
  AND2_X1   g1062(.A1(new_n1173), .A2(new_n1186), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1262), .B1(new_n1263), .B2(new_n1166), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1194), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n911), .A2(new_n667), .A3(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT121), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1264), .A2(new_n1266), .A3(new_n1267), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1260), .A2(new_n1261), .A3(new_n1196), .A4(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1189), .A2(new_n1037), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n784), .B1(new_n887), .B2(G68), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(G58), .A2(new_n823), .B1(new_n826), .B2(G128), .ZN(new_n1272));
  OAI221_X1 g1072(.A(new_n1272), .B1(new_n1057), .B2(new_n820), .C1(new_n799), .C2(new_n871), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(new_n865), .A2(new_n1139), .B1(new_n813), .B2(G132), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n350), .B1(new_n833), .B2(G50), .ZN(new_n1275));
  OAI211_X1 g1075(.A(new_n1274), .B(new_n1275), .C1(new_n1143), .C2(new_n804), .ZN(new_n1276));
  AOI22_X1  g1076(.A1(G97), .A2(new_n835), .B1(new_n823), .B2(G77), .ZN(new_n1277));
  OAI221_X1 g1077(.A(new_n1277), .B1(new_n322), .B2(new_n820), .C1(new_n876), .C2(new_n798), .ZN(new_n1278));
  AOI22_X1  g1078(.A1(G294), .A2(new_n813), .B1(new_n1049), .B2(G283), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n254), .B1(new_n865), .B2(G116), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1279), .A2(new_n1098), .A3(new_n1280), .ZN(new_n1281));
  OAI22_X1  g1081(.A1(new_n1273), .A2(new_n1276), .B1(new_n1278), .B2(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1271), .B1(new_n1282), .B2(new_n791), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1283), .B1(new_n961), .B2(new_n840), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1270), .A2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1269), .A2(new_n1286), .ZN(G381));
  NOR2_X1   g1087(.A1(G375), .A2(G378), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1038), .A2(new_n1112), .A3(new_n1066), .A4(new_n1135), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  OR2_X1    g1090(.A1(G393), .A2(G396), .ZN(new_n1291));
  NOR3_X1   g1091(.A1(new_n1291), .A2(G384), .A3(G381), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1288), .A2(new_n1290), .A3(new_n1292), .ZN(G407));
  INV_X1    g1093(.A(G213), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1294), .A2(G343), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1288), .A2(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(G407), .A2(G213), .A3(new_n1296), .ZN(G409));
  NAND2_X1  g1097(.A1(G393), .A2(G396), .ZN(new_n1298));
  AND2_X1   g1098(.A1(new_n1291), .A2(new_n1298), .ZN(new_n1299));
  AOI22_X1  g1099(.A1(new_n1038), .A2(new_n1066), .B1(new_n1112), .B2(new_n1135), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1299), .B1(new_n1290), .B2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT61), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(G387), .A2(G390), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1291), .A2(new_n1298), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1303), .A2(new_n1289), .A3(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1301), .A2(new_n1302), .A3(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1201), .A2(new_n1261), .A3(new_n1228), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(new_n1256), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(new_n1199), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(KEYINPUT123), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT123), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1308), .A2(new_n1311), .A3(new_n1199), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1310), .A2(new_n1312), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1231), .A2(G378), .A3(new_n1256), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT122), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1231), .A2(KEYINPUT122), .A3(G378), .A4(new_n1256), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1313), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1264), .A2(new_n1266), .ZN(new_n1319));
  XNOR2_X1  g1119(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n1320));
  OAI211_X1 g1120(.A(new_n1260), .B(new_n1268), .C1(new_n1319), .C2(new_n1320), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1189), .A2(new_n1195), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n729), .B1(new_n1322), .B2(KEYINPUT60), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1321), .A2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(new_n1286), .ZN(new_n1325));
  OAI21_X1  g1125(.A(KEYINPUT125), .B1(new_n1325), .B2(new_n892), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT125), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(G384), .A2(new_n1327), .A3(new_n1286), .A4(new_n1324), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1325), .A2(new_n892), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1326), .A2(new_n1328), .A3(new_n1329), .ZN(new_n1330));
  NOR3_X1   g1130(.A1(new_n1318), .A2(new_n1295), .A3(new_n1330), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1306), .B1(new_n1331), .B2(KEYINPUT63), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1295), .A2(G2897), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1330), .A2(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1333), .ZN(new_n1335));
  NAND4_X1  g1135(.A1(new_n1326), .A2(new_n1328), .A3(new_n1329), .A4(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1334), .A2(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT126), .ZN(new_n1338));
  OAI211_X1 g1138(.A(new_n1337), .B(new_n1338), .C1(new_n1318), .C2(new_n1295), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1337), .B1(new_n1318), .B2(new_n1295), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1340), .A2(KEYINPUT126), .ZN(new_n1341));
  AND2_X1   g1141(.A1(new_n1310), .A2(new_n1312), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1256), .ZN(new_n1343));
  AND2_X1   g1143(.A1(new_n1221), .A2(new_n1227), .ZN(new_n1344));
  AND3_X1   g1144(.A1(new_n1176), .A2(new_n1179), .A3(new_n1173), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n1173), .B1(new_n1176), .B2(new_n1179), .ZN(new_n1346));
  NOR2_X1   g1146(.A1(new_n1345), .A2(new_n1346), .ZN(new_n1347));
  AOI21_X1  g1147(.A(new_n1266), .B1(new_n1347), .B2(new_n1319), .ZN(new_n1348));
  OAI21_X1  g1148(.A(KEYINPUT57), .B1(new_n1344), .B2(new_n1348), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1201), .A2(new_n1202), .A3(new_n1228), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1349), .A2(new_n1350), .ZN(new_n1351));
  AOI21_X1  g1151(.A(new_n1343), .B1(new_n1351), .B2(new_n728), .ZN(new_n1352));
  AOI21_X1  g1152(.A(KEYINPUT122), .B1(new_n1352), .B2(G378), .ZN(new_n1353));
  INV_X1    g1153(.A(new_n1317), .ZN(new_n1354));
  OAI21_X1  g1154(.A(new_n1342), .B1(new_n1353), .B2(new_n1354), .ZN(new_n1355));
  INV_X1    g1155(.A(new_n1295), .ZN(new_n1356));
  INV_X1    g1156(.A(new_n1330), .ZN(new_n1357));
  NAND3_X1  g1157(.A1(new_n1355), .A2(new_n1356), .A3(new_n1357), .ZN(new_n1358));
  INV_X1    g1158(.A(KEYINPUT63), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1358), .A2(new_n1359), .ZN(new_n1360));
  NAND4_X1  g1160(.A1(new_n1332), .A2(new_n1339), .A3(new_n1341), .A4(new_n1360), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1301), .A2(new_n1305), .ZN(new_n1362));
  INV_X1    g1162(.A(KEYINPUT62), .ZN(new_n1363));
  NAND4_X1  g1163(.A1(new_n1355), .A2(new_n1363), .A3(new_n1356), .A4(new_n1357), .ZN(new_n1364));
  XOR2_X1   g1164(.A(KEYINPUT127), .B(KEYINPUT61), .Z(new_n1365));
  NAND3_X1  g1165(.A1(new_n1364), .A2(new_n1340), .A3(new_n1365), .ZN(new_n1366));
  NOR2_X1   g1166(.A1(new_n1318), .A2(new_n1295), .ZN(new_n1367));
  AOI21_X1  g1167(.A(new_n1363), .B1(new_n1367), .B2(new_n1357), .ZN(new_n1368));
  OAI21_X1  g1168(.A(new_n1362), .B1(new_n1366), .B2(new_n1368), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1361), .A2(new_n1369), .ZN(G405));
  NAND2_X1  g1170(.A1(G375), .A2(new_n1199), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1372));
  AOI21_X1  g1172(.A(new_n1330), .B1(new_n1371), .B2(new_n1372), .ZN(new_n1373));
  INV_X1    g1173(.A(new_n1373), .ZN(new_n1374));
  NAND3_X1  g1174(.A1(new_n1371), .A2(new_n1372), .A3(new_n1330), .ZN(new_n1375));
  NAND4_X1  g1175(.A1(new_n1374), .A2(new_n1301), .A3(new_n1305), .A4(new_n1375), .ZN(new_n1376));
  INV_X1    g1176(.A(new_n1375), .ZN(new_n1377));
  OAI21_X1  g1177(.A(new_n1362), .B1(new_n1377), .B2(new_n1373), .ZN(new_n1378));
  NAND2_X1  g1178(.A1(new_n1376), .A2(new_n1378), .ZN(G402));
endmodule


