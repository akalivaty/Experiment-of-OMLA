

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U553 ( .A1(G2105), .A2(G2104), .ZN(n532) );
  AND2_X1 U554 ( .A1(n536), .A2(G2105), .ZN(n884) );
  NOR2_X2 U555 ( .A1(n747), .A2(n694), .ZN(n696) );
  NOR2_X1 U556 ( .A1(n728), .A2(n727), .ZN(n730) );
  NOR2_X1 U557 ( .A1(G2105), .A2(n536), .ZN(n610) );
  XNOR2_X2 U558 ( .A(n692), .B(n792), .ZN(n693) );
  AND2_X1 U559 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U560 ( .A(n718), .B(n717), .ZN(n722) );
  INV_X1 U561 ( .A(KEYINPUT95), .ZN(n717) );
  NOR2_X1 U562 ( .A1(n743), .A2(n526), .ZN(n744) );
  NOR2_X1 U563 ( .A1(G651), .A2(n656), .ZN(n655) );
  XNOR2_X1 U564 ( .A(n535), .B(KEYINPUT87), .ZN(n539) );
  NAND2_X1 U565 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U566 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U567 ( .A(n746), .B(n741), .Z(n523) );
  AND2_X1 U568 ( .A1(n815), .A2(n814), .ZN(n524) );
  XNOR2_X2 U569 ( .A(n561), .B(KEYINPUT65), .ZN(G160) );
  AND2_X1 U570 ( .A1(n538), .A2(n537), .ZN(n525) );
  AND2_X1 U571 ( .A1(G8), .A2(n742), .ZN(n526) );
  AND2_X1 U572 ( .A1(n780), .A2(n779), .ZN(n527) );
  NOR2_X1 U573 ( .A1(n774), .A2(n773), .ZN(n528) );
  AND2_X1 U574 ( .A1(n768), .A2(n956), .ZN(n529) );
  INV_X1 U575 ( .A(KEYINPUT26), .ZN(n695) );
  XNOR2_X1 U576 ( .A(n696), .B(n695), .ZN(n699) );
  INV_X1 U577 ( .A(KEYINPUT64), .ZN(n700) );
  INV_X1 U578 ( .A(KEYINPUT96), .ZN(n729) );
  INV_X1 U579 ( .A(KEYINPUT98), .ZN(n741) );
  NAND2_X1 U580 ( .A1(n523), .A2(n744), .ZN(n757) );
  INV_X1 U581 ( .A(n778), .ZN(n769) );
  INV_X1 U582 ( .A(KEYINPUT33), .ZN(n770) );
  INV_X1 U583 ( .A(n822), .ZN(n814) );
  INV_X1 U584 ( .A(KEYINPUT17), .ZN(n531) );
  NAND2_X1 U585 ( .A1(n573), .A2(n572), .ZN(n966) );
  AND2_X1 U586 ( .A1(n539), .A2(n525), .ZN(G164) );
  INV_X1 U587 ( .A(G2104), .ZN(n536) );
  NAND2_X1 U588 ( .A1(n610), .A2(G102), .ZN(n530) );
  XNOR2_X1 U589 ( .A(n530), .B(KEYINPUT86), .ZN(n534) );
  XNOR2_X2 U590 ( .A(n532), .B(n531), .ZN(n889) );
  NAND2_X1 U591 ( .A1(n889), .A2(G138), .ZN(n533) );
  NAND2_X1 U592 ( .A1(n534), .A2(n533), .ZN(n535) );
  NAND2_X1 U593 ( .A1(G126), .A2(n884), .ZN(n538) );
  AND2_X1 U594 ( .A1(G2105), .A2(G2104), .ZN(n885) );
  NAND2_X1 U595 ( .A1(G114), .A2(n885), .ZN(n537) );
  AND2_X1 U596 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U597 ( .A(G57), .ZN(G237) );
  INV_X1 U598 ( .A(G132), .ZN(G219) );
  INV_X1 U599 ( .A(G82), .ZN(G220) );
  XOR2_X1 U600 ( .A(G543), .B(KEYINPUT0), .Z(n656) );
  NAND2_X1 U601 ( .A1(G51), .A2(n655), .ZN(n542) );
  INV_X1 U602 ( .A(G651), .ZN(n546) );
  NOR2_X1 U603 ( .A1(G543), .A2(n546), .ZN(n540) );
  XOR2_X2 U604 ( .A(KEYINPUT1), .B(n540), .Z(n660) );
  NAND2_X1 U605 ( .A1(G63), .A2(n660), .ZN(n541) );
  NAND2_X1 U606 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U607 ( .A(n543), .B(KEYINPUT73), .ZN(n544) );
  XNOR2_X1 U608 ( .A(n544), .B(KEYINPUT6), .ZN(n552) );
  XNOR2_X1 U609 ( .A(KEYINPUT72), .B(KEYINPUT5), .ZN(n550) );
  NOR2_X1 U610 ( .A1(G651), .A2(G543), .ZN(n650) );
  NAND2_X1 U611 ( .A1(n650), .A2(G89), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n545), .B(KEYINPUT4), .ZN(n548) );
  NOR2_X1 U613 ( .A1(n656), .A2(n546), .ZN(n649) );
  NAND2_X1 U614 ( .A1(G76), .A2(n649), .ZN(n547) );
  NAND2_X1 U615 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(n551) );
  NAND2_X1 U617 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U618 ( .A(KEYINPUT7), .B(n553), .ZN(G168) );
  XOR2_X1 U619 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U620 ( .A1(n889), .A2(G137), .ZN(n555) );
  NAND2_X1 U621 ( .A1(G125), .A2(n884), .ZN(n554) );
  AND2_X1 U622 ( .A1(n555), .A2(n554), .ZN(n560) );
  NAND2_X1 U623 ( .A1(G101), .A2(n610), .ZN(n556) );
  XNOR2_X1 U624 ( .A(KEYINPUT23), .B(n556), .ZN(n558) );
  AND2_X1 U625 ( .A1(G113), .A2(n885), .ZN(n557) );
  NAND2_X1 U626 ( .A1(G7), .A2(G661), .ZN(n562) );
  XNOR2_X1 U627 ( .A(n562), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U628 ( .A(G223), .ZN(n834) );
  NAND2_X1 U629 ( .A1(n834), .A2(G567), .ZN(n563) );
  XOR2_X1 U630 ( .A(KEYINPUT11), .B(n563), .Z(G234) );
  NAND2_X1 U631 ( .A1(n660), .A2(G56), .ZN(n564) );
  XNOR2_X1 U632 ( .A(KEYINPUT14), .B(n564), .ZN(n570) );
  NAND2_X1 U633 ( .A1(n650), .A2(G81), .ZN(n565) );
  XNOR2_X1 U634 ( .A(n565), .B(KEYINPUT12), .ZN(n567) );
  NAND2_X1 U635 ( .A1(G68), .A2(n649), .ZN(n566) );
  NAND2_X1 U636 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U637 ( .A(KEYINPUT13), .B(n568), .ZN(n569) );
  NAND2_X1 U638 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U639 ( .A(n571), .B(KEYINPUT69), .ZN(n573) );
  NAND2_X1 U640 ( .A1(n655), .A2(G43), .ZN(n572) );
  INV_X1 U641 ( .A(G860), .ZN(n602) );
  OR2_X1 U642 ( .A1(n966), .A2(n602), .ZN(n574) );
  XNOR2_X1 U643 ( .A(KEYINPUT70), .B(n574), .ZN(G153) );
  NAND2_X1 U644 ( .A1(G77), .A2(n649), .ZN(n576) );
  NAND2_X1 U645 ( .A1(G90), .A2(n650), .ZN(n575) );
  NAND2_X1 U646 ( .A1(n576), .A2(n575), .ZN(n578) );
  XOR2_X1 U647 ( .A(KEYINPUT9), .B(KEYINPUT67), .Z(n577) );
  XNOR2_X1 U648 ( .A(n578), .B(n577), .ZN(n582) );
  NAND2_X1 U649 ( .A1(n655), .A2(G52), .ZN(n580) );
  NAND2_X1 U650 ( .A1(G64), .A2(n660), .ZN(n579) );
  AND2_X1 U651 ( .A1(n580), .A2(n579), .ZN(n581) );
  NAND2_X1 U652 ( .A1(n582), .A2(n581), .ZN(G301) );
  NAND2_X1 U653 ( .A1(G868), .A2(G301), .ZN(n592) );
  NAND2_X1 U654 ( .A1(n655), .A2(G54), .ZN(n589) );
  NAND2_X1 U655 ( .A1(G79), .A2(n649), .ZN(n584) );
  NAND2_X1 U656 ( .A1(G66), .A2(n660), .ZN(n583) );
  NAND2_X1 U657 ( .A1(n584), .A2(n583), .ZN(n587) );
  NAND2_X1 U658 ( .A1(G92), .A2(n650), .ZN(n585) );
  XNOR2_X1 U659 ( .A(KEYINPUT71), .B(n585), .ZN(n586) );
  NOR2_X1 U660 ( .A1(n587), .A2(n586), .ZN(n588) );
  NAND2_X1 U661 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U662 ( .A(KEYINPUT15), .B(n590), .Z(n904) );
  INV_X1 U663 ( .A(G868), .ZN(n674) );
  NAND2_X1 U664 ( .A1(n904), .A2(n674), .ZN(n591) );
  NAND2_X1 U665 ( .A1(n592), .A2(n591), .ZN(G284) );
  NAND2_X1 U666 ( .A1(G65), .A2(n660), .ZN(n594) );
  NAND2_X1 U667 ( .A1(G91), .A2(n650), .ZN(n593) );
  NAND2_X1 U668 ( .A1(n594), .A2(n593), .ZN(n597) );
  NAND2_X1 U669 ( .A1(n649), .A2(G78), .ZN(n595) );
  XOR2_X1 U670 ( .A(KEYINPUT68), .B(n595), .Z(n596) );
  NOR2_X1 U671 ( .A1(n597), .A2(n596), .ZN(n599) );
  NAND2_X1 U672 ( .A1(n655), .A2(G53), .ZN(n598) );
  NAND2_X1 U673 ( .A1(n599), .A2(n598), .ZN(G299) );
  NOR2_X1 U674 ( .A1(G286), .A2(n674), .ZN(n601) );
  NOR2_X1 U675 ( .A1(G868), .A2(G299), .ZN(n600) );
  NOR2_X1 U676 ( .A1(n601), .A2(n600), .ZN(G297) );
  NAND2_X1 U677 ( .A1(n602), .A2(G559), .ZN(n603) );
  INV_X1 U678 ( .A(n904), .ZN(n952) );
  NAND2_X1 U679 ( .A1(n603), .A2(n952), .ZN(n604) );
  XNOR2_X1 U680 ( .A(n604), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U681 ( .A1(G868), .A2(n966), .ZN(n607) );
  NAND2_X1 U682 ( .A1(G868), .A2(n952), .ZN(n605) );
  NOR2_X1 U683 ( .A1(G559), .A2(n605), .ZN(n606) );
  NOR2_X1 U684 ( .A1(n607), .A2(n606), .ZN(G282) );
  NAND2_X1 U685 ( .A1(G123), .A2(n884), .ZN(n608) );
  XNOR2_X1 U686 ( .A(n608), .B(KEYINPUT18), .ZN(n609) );
  XNOR2_X1 U687 ( .A(n609), .B(KEYINPUT74), .ZN(n612) );
  BUF_X1 U688 ( .A(n610), .Z(n892) );
  NAND2_X1 U689 ( .A1(G99), .A2(n892), .ZN(n611) );
  NAND2_X1 U690 ( .A1(n612), .A2(n611), .ZN(n616) );
  NAND2_X1 U691 ( .A1(G135), .A2(n889), .ZN(n614) );
  NAND2_X1 U692 ( .A1(G111), .A2(n885), .ZN(n613) );
  NAND2_X1 U693 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U694 ( .A1(n616), .A2(n615), .ZN(n1014) );
  XNOR2_X1 U695 ( .A(n1014), .B(G2096), .ZN(n618) );
  INV_X1 U696 ( .A(G2100), .ZN(n617) );
  NAND2_X1 U697 ( .A1(n618), .A2(n617), .ZN(G156) );
  NAND2_X1 U698 ( .A1(G93), .A2(n650), .ZN(n619) );
  XNOR2_X1 U699 ( .A(n619), .B(KEYINPUT76), .ZN(n621) );
  NAND2_X1 U700 ( .A1(n660), .A2(G67), .ZN(n620) );
  NAND2_X1 U701 ( .A1(n621), .A2(n620), .ZN(n625) );
  NAND2_X1 U702 ( .A1(G80), .A2(n649), .ZN(n623) );
  NAND2_X1 U703 ( .A1(G55), .A2(n655), .ZN(n622) );
  NAND2_X1 U704 ( .A1(n623), .A2(n622), .ZN(n624) );
  OR2_X1 U705 ( .A1(n625), .A2(n624), .ZN(n675) );
  NAND2_X1 U706 ( .A1(n952), .A2(G559), .ZN(n671) );
  XNOR2_X1 U707 ( .A(n966), .B(n671), .ZN(n626) );
  NOR2_X1 U708 ( .A1(G860), .A2(n626), .ZN(n627) );
  XOR2_X1 U709 ( .A(KEYINPUT75), .B(n627), .Z(n628) );
  XOR2_X1 U710 ( .A(n675), .B(n628), .Z(G145) );
  NAND2_X1 U711 ( .A1(n650), .A2(G86), .ZN(n637) );
  NAND2_X1 U712 ( .A1(G73), .A2(n649), .ZN(n629) );
  XNOR2_X1 U713 ( .A(n629), .B(KEYINPUT2), .ZN(n632) );
  NAND2_X1 U714 ( .A1(G48), .A2(n655), .ZN(n630) );
  XNOR2_X1 U715 ( .A(n630), .B(KEYINPUT78), .ZN(n631) );
  NAND2_X1 U716 ( .A1(n632), .A2(n631), .ZN(n635) );
  NAND2_X1 U717 ( .A1(G61), .A2(n660), .ZN(n633) );
  XNOR2_X1 U718 ( .A(KEYINPUT77), .B(n633), .ZN(n634) );
  NOR2_X1 U719 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U720 ( .A1(n637), .A2(n636), .ZN(n638) );
  XOR2_X1 U721 ( .A(KEYINPUT79), .B(n638), .Z(G305) );
  NAND2_X1 U722 ( .A1(G60), .A2(n660), .ZN(n640) );
  NAND2_X1 U723 ( .A1(G85), .A2(n650), .ZN(n639) );
  NAND2_X1 U724 ( .A1(n640), .A2(n639), .ZN(n644) );
  NAND2_X1 U725 ( .A1(G72), .A2(n649), .ZN(n642) );
  NAND2_X1 U726 ( .A1(G47), .A2(n655), .ZN(n641) );
  NAND2_X1 U727 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U728 ( .A1(n644), .A2(n643), .ZN(n645) );
  XOR2_X1 U729 ( .A(KEYINPUT66), .B(n645), .Z(G290) );
  NAND2_X1 U730 ( .A1(G50), .A2(n655), .ZN(n647) );
  NAND2_X1 U731 ( .A1(G62), .A2(n660), .ZN(n646) );
  NAND2_X1 U732 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U733 ( .A(KEYINPUT80), .B(n648), .ZN(n654) );
  NAND2_X1 U734 ( .A1(G75), .A2(n649), .ZN(n652) );
  NAND2_X1 U735 ( .A1(G88), .A2(n650), .ZN(n651) );
  NAND2_X1 U736 ( .A1(n652), .A2(n651), .ZN(n653) );
  NOR2_X1 U737 ( .A1(n654), .A2(n653), .ZN(G166) );
  NAND2_X1 U738 ( .A1(G49), .A2(n655), .ZN(n658) );
  NAND2_X1 U739 ( .A1(G87), .A2(n656), .ZN(n657) );
  NAND2_X1 U740 ( .A1(n658), .A2(n657), .ZN(n659) );
  NOR2_X1 U741 ( .A1(n660), .A2(n659), .ZN(n662) );
  NAND2_X1 U742 ( .A1(G651), .A2(G74), .ZN(n661) );
  NAND2_X1 U743 ( .A1(n662), .A2(n661), .ZN(G288) );
  XOR2_X1 U744 ( .A(KEYINPUT82), .B(KEYINPUT81), .Z(n664) );
  XNOR2_X1 U745 ( .A(G290), .B(KEYINPUT19), .ZN(n663) );
  XNOR2_X1 U746 ( .A(n664), .B(n663), .ZN(n668) );
  INV_X1 U747 ( .A(G299), .ZN(n955) );
  XNOR2_X1 U748 ( .A(G166), .B(n955), .ZN(n665) );
  XOR2_X1 U749 ( .A(n665), .B(n675), .Z(n666) );
  XNOR2_X1 U750 ( .A(n666), .B(n966), .ZN(n667) );
  XNOR2_X1 U751 ( .A(n668), .B(n667), .ZN(n669) );
  XNOR2_X1 U752 ( .A(n669), .B(G288), .ZN(n670) );
  XNOR2_X1 U753 ( .A(G305), .B(n670), .ZN(n905) );
  XNOR2_X1 U754 ( .A(n905), .B(n671), .ZN(n672) );
  NAND2_X1 U755 ( .A1(n672), .A2(G868), .ZN(n673) );
  XOR2_X1 U756 ( .A(KEYINPUT83), .B(n673), .Z(n677) );
  NAND2_X1 U757 ( .A1(n675), .A2(n674), .ZN(n676) );
  NAND2_X1 U758 ( .A1(n677), .A2(n676), .ZN(G295) );
  NAND2_X1 U759 ( .A1(G2084), .A2(G2078), .ZN(n678) );
  XOR2_X1 U760 ( .A(KEYINPUT20), .B(n678), .Z(n679) );
  NAND2_X1 U761 ( .A1(G2090), .A2(n679), .ZN(n680) );
  XNOR2_X1 U762 ( .A(KEYINPUT21), .B(n680), .ZN(n681) );
  NAND2_X1 U763 ( .A1(n681), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U764 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U765 ( .A1(G661), .A2(G483), .ZN(n689) );
  NOR2_X1 U766 ( .A1(G220), .A2(G219), .ZN(n682) );
  XOR2_X1 U767 ( .A(KEYINPUT22), .B(n682), .Z(n683) );
  NOR2_X1 U768 ( .A1(G218), .A2(n683), .ZN(n684) );
  NAND2_X1 U769 ( .A1(G96), .A2(n684), .ZN(n838) );
  NAND2_X1 U770 ( .A1(n838), .A2(G2106), .ZN(n688) );
  NAND2_X1 U771 ( .A1(G69), .A2(G120), .ZN(n685) );
  NOR2_X1 U772 ( .A1(G237), .A2(n685), .ZN(n686) );
  NAND2_X1 U773 ( .A1(G108), .A2(n686), .ZN(n839) );
  NAND2_X1 U774 ( .A1(n839), .A2(G567), .ZN(n687) );
  NAND2_X1 U775 ( .A1(n688), .A2(n687), .ZN(n840) );
  NOR2_X1 U776 ( .A1(n689), .A2(n840), .ZN(n690) );
  XNOR2_X1 U777 ( .A(n690), .B(KEYINPUT84), .ZN(n837) );
  NAND2_X1 U778 ( .A1(n837), .A2(G36), .ZN(n691) );
  XOR2_X1 U779 ( .A(KEYINPUT85), .B(n691), .Z(G176) );
  INV_X1 U780 ( .A(G166), .ZN(G303) );
  INV_X1 U781 ( .A(KEYINPUT92), .ZN(n692) );
  NAND2_X1 U782 ( .A1(G160), .A2(G40), .ZN(n792) );
  NOR2_X1 U783 ( .A1(G164), .A2(G1384), .ZN(n793) );
  NAND2_X2 U784 ( .A1(n693), .A2(n793), .ZN(n747) );
  INV_X1 U785 ( .A(G1996), .ZN(n694) );
  AND2_X1 U786 ( .A1(n747), .A2(G1341), .ZN(n697) );
  NOR2_X1 U787 ( .A1(n697), .A2(n966), .ZN(n698) );
  AND2_X1 U788 ( .A1(n699), .A2(n698), .ZN(n701) );
  XNOR2_X1 U789 ( .A(n701), .B(n700), .ZN(n708) );
  INV_X1 U790 ( .A(n708), .ZN(n702) );
  NAND2_X1 U791 ( .A1(n702), .A2(n952), .ZN(n707) );
  NAND2_X1 U792 ( .A1(n747), .A2(G1348), .ZN(n703) );
  XNOR2_X1 U793 ( .A(n703), .B(KEYINPUT94), .ZN(n705) );
  INV_X1 U794 ( .A(n747), .ZN(n711) );
  NAND2_X1 U795 ( .A1(n711), .A2(G2067), .ZN(n704) );
  NAND2_X1 U796 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U797 ( .A1(n707), .A2(n706), .ZN(n710) );
  NAND2_X1 U798 ( .A1(n708), .A2(n904), .ZN(n709) );
  NAND2_X1 U799 ( .A1(n710), .A2(n709), .ZN(n716) );
  NAND2_X1 U800 ( .A1(n711), .A2(G2072), .ZN(n712) );
  XNOR2_X1 U801 ( .A(n712), .B(KEYINPUT27), .ZN(n714) );
  AND2_X1 U802 ( .A1(G1956), .A2(n747), .ZN(n713) );
  NOR2_X1 U803 ( .A1(n714), .A2(n713), .ZN(n719) );
  NAND2_X1 U804 ( .A1(n955), .A2(n719), .ZN(n715) );
  NAND2_X1 U805 ( .A1(n716), .A2(n715), .ZN(n718) );
  OR2_X1 U806 ( .A1(n955), .A2(n719), .ZN(n720) );
  XNOR2_X1 U807 ( .A(KEYINPUT28), .B(n720), .ZN(n721) );
  NAND2_X1 U808 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U809 ( .A(n723), .B(KEYINPUT29), .ZN(n728) );
  XOR2_X1 U810 ( .A(G2078), .B(KEYINPUT25), .Z(n926) );
  NOR2_X1 U811 ( .A1(n926), .A2(n747), .ZN(n724) );
  XOR2_X1 U812 ( .A(KEYINPUT93), .B(n724), .Z(n726) );
  NOR2_X1 U813 ( .A1(n711), .A2(G1961), .ZN(n725) );
  NOR2_X1 U814 ( .A1(n726), .A2(n725), .ZN(n731) );
  NOR2_X1 U815 ( .A1(n731), .A2(G301), .ZN(n727) );
  XNOR2_X1 U816 ( .A(n730), .B(n729), .ZN(n740) );
  AND2_X1 U817 ( .A1(G301), .A2(n731), .ZN(n737) );
  NAND2_X1 U818 ( .A1(G8), .A2(n747), .ZN(n778) );
  NOR2_X1 U819 ( .A1(G1966), .A2(n778), .ZN(n743) );
  NOR2_X1 U820 ( .A1(G2084), .A2(n747), .ZN(n742) );
  NOR2_X1 U821 ( .A1(n743), .A2(n742), .ZN(n732) );
  NAND2_X1 U822 ( .A1(G8), .A2(n732), .ZN(n733) );
  XNOR2_X1 U823 ( .A(KEYINPUT30), .B(n733), .ZN(n734) );
  XOR2_X1 U824 ( .A(KEYINPUT97), .B(n734), .Z(n735) );
  NOR2_X1 U825 ( .A1(G168), .A2(n735), .ZN(n736) );
  NOR2_X1 U826 ( .A1(n737), .A2(n736), .ZN(n738) );
  XOR2_X1 U827 ( .A(KEYINPUT31), .B(n738), .Z(n739) );
  NAND2_X1 U828 ( .A1(n740), .A2(n739), .ZN(n746) );
  AND2_X1 U829 ( .A1(G286), .A2(G8), .ZN(n745) );
  NAND2_X1 U830 ( .A1(n746), .A2(n745), .ZN(n754) );
  INV_X1 U831 ( .A(G8), .ZN(n752) );
  NOR2_X1 U832 ( .A1(G1971), .A2(n778), .ZN(n749) );
  NOR2_X1 U833 ( .A1(G2090), .A2(n747), .ZN(n748) );
  NOR2_X1 U834 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U835 ( .A1(n750), .A2(G303), .ZN(n751) );
  OR2_X1 U836 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U837 ( .A(n755), .B(KEYINPUT32), .ZN(n756) );
  NAND2_X1 U838 ( .A1(n757), .A2(n756), .ZN(n767) );
  NOR2_X1 U839 ( .A1(G2090), .A2(G303), .ZN(n758) );
  XOR2_X1 U840 ( .A(KEYINPUT99), .B(n758), .Z(n759) );
  NAND2_X1 U841 ( .A1(G8), .A2(n759), .ZN(n760) );
  NAND2_X1 U842 ( .A1(n767), .A2(n760), .ZN(n761) );
  XNOR2_X1 U843 ( .A(n761), .B(KEYINPUT100), .ZN(n762) );
  NAND2_X1 U844 ( .A1(n762), .A2(n778), .ZN(n763) );
  XNOR2_X1 U845 ( .A(n763), .B(KEYINPUT101), .ZN(n764) );
  INV_X1 U846 ( .A(n764), .ZN(n781) );
  NOR2_X1 U847 ( .A1(G1971), .A2(G303), .ZN(n765) );
  NOR2_X1 U848 ( .A1(G1976), .A2(G288), .ZN(n959) );
  NOR2_X1 U849 ( .A1(n765), .A2(n959), .ZN(n766) );
  NAND2_X1 U850 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U851 ( .A1(G1976), .A2(G288), .ZN(n956) );
  NAND2_X1 U852 ( .A1(n529), .A2(n769), .ZN(n771) );
  NAND2_X1 U853 ( .A1(n771), .A2(n770), .ZN(n775) );
  XOR2_X1 U854 ( .A(G1981), .B(G305), .Z(n948) );
  INV_X1 U855 ( .A(n948), .ZN(n774) );
  NAND2_X1 U856 ( .A1(n959), .A2(KEYINPUT33), .ZN(n772) );
  NOR2_X1 U857 ( .A1(n778), .A2(n772), .ZN(n773) );
  NAND2_X1 U858 ( .A1(n775), .A2(n528), .ZN(n780) );
  NOR2_X1 U859 ( .A1(G1981), .A2(G305), .ZN(n776) );
  XOR2_X1 U860 ( .A(n776), .B(KEYINPUT24), .Z(n777) );
  OR2_X1 U861 ( .A1(n778), .A2(n777), .ZN(n779) );
  NAND2_X1 U862 ( .A1(n781), .A2(n527), .ZN(n816) );
  XOR2_X1 U863 ( .A(G290), .B(G1986), .Z(n961) );
  NAND2_X1 U864 ( .A1(G128), .A2(n884), .ZN(n783) );
  NAND2_X1 U865 ( .A1(G116), .A2(n885), .ZN(n782) );
  NAND2_X1 U866 ( .A1(n783), .A2(n782), .ZN(n784) );
  XNOR2_X1 U867 ( .A(n784), .B(KEYINPUT35), .ZN(n790) );
  NAND2_X1 U868 ( .A1(n892), .A2(G104), .ZN(n785) );
  XOR2_X1 U869 ( .A(KEYINPUT89), .B(n785), .Z(n787) );
  NAND2_X1 U870 ( .A1(n889), .A2(G140), .ZN(n786) );
  NAND2_X1 U871 ( .A1(n787), .A2(n786), .ZN(n788) );
  XOR2_X1 U872 ( .A(KEYINPUT34), .B(n788), .Z(n789) );
  NAND2_X1 U873 ( .A1(n790), .A2(n789), .ZN(n791) );
  XNOR2_X1 U874 ( .A(n791), .B(KEYINPUT36), .ZN(n900) );
  XOR2_X1 U875 ( .A(G2067), .B(KEYINPUT37), .Z(n817) );
  NAND2_X1 U876 ( .A1(n900), .A2(n817), .ZN(n818) );
  NAND2_X1 U877 ( .A1(n961), .A2(n818), .ZN(n795) );
  NOR2_X1 U878 ( .A1(n792), .A2(n793), .ZN(n794) );
  XNOR2_X1 U879 ( .A(n794), .B(KEYINPUT88), .ZN(n829) );
  NAND2_X1 U880 ( .A1(n795), .A2(n829), .ZN(n815) );
  NAND2_X1 U881 ( .A1(G131), .A2(n889), .ZN(n797) );
  NAND2_X1 U882 ( .A1(G119), .A2(n884), .ZN(n796) );
  NAND2_X1 U883 ( .A1(n797), .A2(n796), .ZN(n801) );
  NAND2_X1 U884 ( .A1(G95), .A2(n892), .ZN(n799) );
  NAND2_X1 U885 ( .A1(G107), .A2(n885), .ZN(n798) );
  NAND2_X1 U886 ( .A1(n799), .A2(n798), .ZN(n800) );
  OR2_X1 U887 ( .A1(n801), .A2(n800), .ZN(n871) );
  NAND2_X1 U888 ( .A1(G1991), .A2(n871), .ZN(n802) );
  XNOR2_X1 U889 ( .A(n802), .B(KEYINPUT90), .ZN(n811) );
  NAND2_X1 U890 ( .A1(G141), .A2(n889), .ZN(n804) );
  NAND2_X1 U891 ( .A1(G129), .A2(n884), .ZN(n803) );
  NAND2_X1 U892 ( .A1(n804), .A2(n803), .ZN(n807) );
  NAND2_X1 U893 ( .A1(n892), .A2(G105), .ZN(n805) );
  XOR2_X1 U894 ( .A(KEYINPUT38), .B(n805), .Z(n806) );
  NOR2_X1 U895 ( .A1(n807), .A2(n806), .ZN(n809) );
  NAND2_X1 U896 ( .A1(n885), .A2(G117), .ZN(n808) );
  NAND2_X1 U897 ( .A1(n809), .A2(n808), .ZN(n896) );
  NAND2_X1 U898 ( .A1(G1996), .A2(n896), .ZN(n810) );
  NAND2_X1 U899 ( .A1(n811), .A2(n810), .ZN(n812) );
  XNOR2_X1 U900 ( .A(KEYINPUT91), .B(n812), .ZN(n1012) );
  INV_X1 U901 ( .A(n829), .ZN(n813) );
  NOR2_X1 U902 ( .A1(n1012), .A2(n813), .ZN(n822) );
  NAND2_X1 U903 ( .A1(n816), .A2(n524), .ZN(n832) );
  NOR2_X1 U904 ( .A1(n900), .A2(n817), .ZN(n1028) );
  INV_X1 U905 ( .A(n818), .ZN(n1021) );
  NOR2_X1 U906 ( .A1(G1996), .A2(n896), .ZN(n1009) );
  NOR2_X1 U907 ( .A1(G1991), .A2(n871), .ZN(n1015) );
  NOR2_X1 U908 ( .A1(G290), .A2(G1986), .ZN(n819) );
  XNOR2_X1 U909 ( .A(KEYINPUT102), .B(n819), .ZN(n820) );
  NOR2_X1 U910 ( .A1(n1015), .A2(n820), .ZN(n821) );
  NOR2_X1 U911 ( .A1(n822), .A2(n821), .ZN(n823) );
  NOR2_X1 U912 ( .A1(n1009), .A2(n823), .ZN(n824) );
  XOR2_X1 U913 ( .A(KEYINPUT39), .B(n824), .Z(n825) );
  NOR2_X1 U914 ( .A1(n1021), .A2(n825), .ZN(n826) );
  XOR2_X1 U915 ( .A(KEYINPUT103), .B(n826), .Z(n827) );
  NOR2_X1 U916 ( .A1(n1028), .A2(n827), .ZN(n828) );
  XOR2_X1 U917 ( .A(KEYINPUT104), .B(n828), .Z(n830) );
  NAND2_X1 U918 ( .A1(n830), .A2(n829), .ZN(n831) );
  NAND2_X1 U919 ( .A1(n832), .A2(n831), .ZN(n833) );
  XNOR2_X1 U920 ( .A(n833), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U921 ( .A(G301), .ZN(G171) );
  NAND2_X1 U922 ( .A1(G2106), .A2(n834), .ZN(G217) );
  AND2_X1 U923 ( .A1(G15), .A2(G2), .ZN(n835) );
  NAND2_X1 U924 ( .A1(G661), .A2(n835), .ZN(G259) );
  NAND2_X1 U925 ( .A1(G3), .A2(G1), .ZN(n836) );
  NAND2_X1 U926 ( .A1(n837), .A2(n836), .ZN(G188) );
  INV_X1 U928 ( .A(G120), .ZN(G236) );
  INV_X1 U929 ( .A(G96), .ZN(G221) );
  INV_X1 U930 ( .A(G69), .ZN(G235) );
  NOR2_X1 U931 ( .A1(n839), .A2(n838), .ZN(G325) );
  INV_X1 U932 ( .A(G325), .ZN(G261) );
  INV_X1 U933 ( .A(n840), .ZN(G319) );
  XNOR2_X1 U934 ( .A(G1971), .B(G2474), .ZN(n850) );
  XOR2_X1 U935 ( .A(G1986), .B(G1956), .Z(n842) );
  XNOR2_X1 U936 ( .A(G1976), .B(G1961), .ZN(n841) );
  XNOR2_X1 U937 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U938 ( .A(G1991), .B(G1996), .Z(n844) );
  XNOR2_X1 U939 ( .A(G1981), .B(G1966), .ZN(n843) );
  XNOR2_X1 U940 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U941 ( .A(n846), .B(n845), .Z(n848) );
  XNOR2_X1 U942 ( .A(KEYINPUT108), .B(KEYINPUT41), .ZN(n847) );
  XNOR2_X1 U943 ( .A(n848), .B(n847), .ZN(n849) );
  XNOR2_X1 U944 ( .A(n850), .B(n849), .ZN(G229) );
  XOR2_X1 U945 ( .A(G2100), .B(KEYINPUT107), .Z(n852) );
  XNOR2_X1 U946 ( .A(KEYINPUT106), .B(G2678), .ZN(n851) );
  XNOR2_X1 U947 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U948 ( .A(KEYINPUT42), .B(G2090), .Z(n854) );
  XNOR2_X1 U949 ( .A(G2067), .B(G2072), .ZN(n853) );
  XNOR2_X1 U950 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U951 ( .A(n856), .B(n855), .Z(n858) );
  XNOR2_X1 U952 ( .A(KEYINPUT43), .B(G2096), .ZN(n857) );
  XNOR2_X1 U953 ( .A(n858), .B(n857), .ZN(n860) );
  XOR2_X1 U954 ( .A(G2084), .B(G2078), .Z(n859) );
  XNOR2_X1 U955 ( .A(n860), .B(n859), .ZN(G227) );
  NAND2_X1 U956 ( .A1(G124), .A2(n884), .ZN(n861) );
  XNOR2_X1 U957 ( .A(n861), .B(KEYINPUT44), .ZN(n863) );
  NAND2_X1 U958 ( .A1(n892), .A2(G100), .ZN(n862) );
  NAND2_X1 U959 ( .A1(n863), .A2(n862), .ZN(n867) );
  NAND2_X1 U960 ( .A1(G136), .A2(n889), .ZN(n865) );
  NAND2_X1 U961 ( .A1(G112), .A2(n885), .ZN(n864) );
  NAND2_X1 U962 ( .A1(n865), .A2(n864), .ZN(n866) );
  NOR2_X1 U963 ( .A1(n867), .A2(n866), .ZN(G162) );
  XOR2_X1 U964 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n869) );
  XNOR2_X1 U965 ( .A(KEYINPUT112), .B(KEYINPUT111), .ZN(n868) );
  XNOR2_X1 U966 ( .A(n869), .B(n868), .ZN(n870) );
  XNOR2_X1 U967 ( .A(n871), .B(n870), .ZN(n873) );
  XNOR2_X1 U968 ( .A(G164), .B(G160), .ZN(n872) );
  XNOR2_X1 U969 ( .A(n873), .B(n872), .ZN(n883) );
  NAND2_X1 U970 ( .A1(G130), .A2(n884), .ZN(n875) );
  NAND2_X1 U971 ( .A1(G118), .A2(n885), .ZN(n874) );
  NAND2_X1 U972 ( .A1(n875), .A2(n874), .ZN(n881) );
  NAND2_X1 U973 ( .A1(n889), .A2(G142), .ZN(n876) );
  XOR2_X1 U974 ( .A(KEYINPUT109), .B(n876), .Z(n878) );
  NAND2_X1 U975 ( .A1(n892), .A2(G106), .ZN(n877) );
  NAND2_X1 U976 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U977 ( .A(n879), .B(KEYINPUT45), .Z(n880) );
  NOR2_X1 U978 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U979 ( .A(n883), .B(n882), .Z(n902) );
  XNOR2_X1 U980 ( .A(n1014), .B(G162), .ZN(n898) );
  NAND2_X1 U981 ( .A1(G127), .A2(n884), .ZN(n887) );
  NAND2_X1 U982 ( .A1(G115), .A2(n885), .ZN(n886) );
  NAND2_X1 U983 ( .A1(n887), .A2(n886), .ZN(n888) );
  XNOR2_X1 U984 ( .A(n888), .B(KEYINPUT47), .ZN(n891) );
  NAND2_X1 U985 ( .A1(G139), .A2(n889), .ZN(n890) );
  NAND2_X1 U986 ( .A1(n891), .A2(n890), .ZN(n895) );
  NAND2_X1 U987 ( .A1(n892), .A2(G103), .ZN(n893) );
  XOR2_X1 U988 ( .A(KEYINPUT110), .B(n893), .Z(n894) );
  NOR2_X1 U989 ( .A1(n895), .A2(n894), .ZN(n1004) );
  XNOR2_X1 U990 ( .A(n896), .B(n1004), .ZN(n897) );
  XNOR2_X1 U991 ( .A(n898), .B(n897), .ZN(n899) );
  XNOR2_X1 U992 ( .A(n900), .B(n899), .ZN(n901) );
  XNOR2_X1 U993 ( .A(n902), .B(n901), .ZN(n903) );
  NOR2_X1 U994 ( .A1(G37), .A2(n903), .ZN(G395) );
  XNOR2_X1 U995 ( .A(G286), .B(n904), .ZN(n906) );
  XNOR2_X1 U996 ( .A(n906), .B(n905), .ZN(n907) );
  XNOR2_X1 U997 ( .A(n907), .B(G171), .ZN(n908) );
  NOR2_X1 U998 ( .A1(G37), .A2(n908), .ZN(G397) );
  XOR2_X1 U999 ( .A(KEYINPUT105), .B(G2427), .Z(n910) );
  XNOR2_X1 U1000 ( .A(G2435), .B(G2438), .ZN(n909) );
  XNOR2_X1 U1001 ( .A(n910), .B(n909), .ZN(n917) );
  XOR2_X1 U1002 ( .A(G2443), .B(G2430), .Z(n912) );
  XNOR2_X1 U1003 ( .A(G2454), .B(G2446), .ZN(n911) );
  XNOR2_X1 U1004 ( .A(n912), .B(n911), .ZN(n913) );
  XOR2_X1 U1005 ( .A(n913), .B(G2451), .Z(n915) );
  XNOR2_X1 U1006 ( .A(G1348), .B(G1341), .ZN(n914) );
  XNOR2_X1 U1007 ( .A(n915), .B(n914), .ZN(n916) );
  XNOR2_X1 U1008 ( .A(n917), .B(n916), .ZN(n918) );
  NAND2_X1 U1009 ( .A1(n918), .A2(G14), .ZN(n924) );
  NAND2_X1 U1010 ( .A1(G319), .A2(n924), .ZN(n921) );
  NOR2_X1 U1011 ( .A1(G229), .A2(G227), .ZN(n919) );
  XNOR2_X1 U1012 ( .A(KEYINPUT49), .B(n919), .ZN(n920) );
  NOR2_X1 U1013 ( .A1(n921), .A2(n920), .ZN(n923) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n922) );
  NAND2_X1 U1015 ( .A1(n923), .A2(n922), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  INV_X1 U1017 ( .A(G108), .ZN(G238) );
  INV_X1 U1018 ( .A(n924), .ZN(G401) );
  XOR2_X1 U1019 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n1036) );
  INV_X1 U1020 ( .A(KEYINPUT55), .ZN(n1030) );
  XOR2_X1 U1021 ( .A(KEYINPUT53), .B(KEYINPUT120), .Z(n938) );
  XNOR2_X1 U1022 ( .A(G2072), .B(KEYINPUT118), .ZN(n925) );
  XNOR2_X1 U1023 ( .A(n925), .B(G33), .ZN(n931) );
  XNOR2_X1 U1024 ( .A(n926), .B(G27), .ZN(n928) );
  XNOR2_X1 U1025 ( .A(G32), .B(G1996), .ZN(n927) );
  NOR2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1027 ( .A(KEYINPUT119), .B(n929), .ZN(n930) );
  NOR2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n936) );
  XOR2_X1 U1029 ( .A(G2067), .B(G26), .Z(n932) );
  NAND2_X1 U1030 ( .A1(n932), .A2(G28), .ZN(n934) );
  XNOR2_X1 U1031 ( .A(G25), .B(G1991), .ZN(n933) );
  NOR2_X1 U1032 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1033 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1034 ( .A(n938), .B(n937), .ZN(n940) );
  XNOR2_X1 U1035 ( .A(G35), .B(G2090), .ZN(n939) );
  NOR2_X1 U1036 ( .A1(n940), .A2(n939), .ZN(n943) );
  XOR2_X1 U1037 ( .A(G2084), .B(KEYINPUT54), .Z(n941) );
  XNOR2_X1 U1038 ( .A(G34), .B(n941), .ZN(n942) );
  NAND2_X1 U1039 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1040 ( .A(n1030), .B(n944), .ZN(n946) );
  INV_X1 U1041 ( .A(G29), .ZN(n945) );
  NAND2_X1 U1042 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1043 ( .A1(G11), .A2(n947), .ZN(n1002) );
  XNOR2_X1 U1044 ( .A(G16), .B(KEYINPUT56), .ZN(n972) );
  XNOR2_X1 U1045 ( .A(G1966), .B(G168), .ZN(n949) );
  NAND2_X1 U1046 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1047 ( .A(n950), .B(KEYINPUT57), .ZN(n970) );
  XNOR2_X1 U1048 ( .A(G303), .B(G1971), .ZN(n951) );
  XNOR2_X1 U1049 ( .A(n951), .B(KEYINPUT121), .ZN(n965) );
  XNOR2_X1 U1050 ( .A(G1348), .B(n952), .ZN(n954) );
  XNOR2_X1 U1051 ( .A(G171), .B(G1961), .ZN(n953) );
  NAND2_X1 U1052 ( .A1(n954), .A2(n953), .ZN(n963) );
  XNOR2_X1 U1053 ( .A(G1956), .B(n955), .ZN(n957) );
  NAND2_X1 U1054 ( .A1(n957), .A2(n956), .ZN(n958) );
  NOR2_X1 U1055 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n962) );
  NOR2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1058 ( .A1(n965), .A2(n964), .ZN(n968) );
  XNOR2_X1 U1059 ( .A(G1341), .B(n966), .ZN(n967) );
  NOR2_X1 U1060 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1061 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1062 ( .A1(n972), .A2(n971), .ZN(n1000) );
  INV_X1 U1063 ( .A(G16), .ZN(n998) );
  XOR2_X1 U1064 ( .A(G1966), .B(KEYINPUT124), .Z(n973) );
  XNOR2_X1 U1065 ( .A(G21), .B(n973), .ZN(n994) );
  XOR2_X1 U1066 ( .A(G1961), .B(G5), .Z(n985) );
  XOR2_X1 U1067 ( .A(KEYINPUT123), .B(G4), .Z(n975) );
  XNOR2_X1 U1068 ( .A(G1348), .B(KEYINPUT59), .ZN(n974) );
  XNOR2_X1 U1069 ( .A(n975), .B(n974), .ZN(n979) );
  XNOR2_X1 U1070 ( .A(G1341), .B(G19), .ZN(n977) );
  XNOR2_X1 U1071 ( .A(G1956), .B(G20), .ZN(n976) );
  NOR2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1073 ( .A1(n979), .A2(n978), .ZN(n982) );
  XNOR2_X1 U1074 ( .A(KEYINPUT122), .B(G1981), .ZN(n980) );
  XNOR2_X1 U1075 ( .A(G6), .B(n980), .ZN(n981) );
  NOR2_X1 U1076 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1077 ( .A(KEYINPUT60), .B(n983), .ZN(n984) );
  NAND2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n992) );
  XNOR2_X1 U1079 ( .A(G1976), .B(G23), .ZN(n987) );
  XNOR2_X1 U1080 ( .A(G1971), .B(G22), .ZN(n986) );
  NOR2_X1 U1081 ( .A1(n987), .A2(n986), .ZN(n989) );
  XOR2_X1 U1082 ( .A(G1986), .B(G24), .Z(n988) );
  NAND2_X1 U1083 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1084 ( .A(KEYINPUT58), .B(n990), .ZN(n991) );
  NOR2_X1 U1085 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1087 ( .A(n995), .B(KEYINPUT125), .ZN(n996) );
  XNOR2_X1 U1088 ( .A(KEYINPUT61), .B(n996), .ZN(n997) );
  NAND2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NOR2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1034) );
  XNOR2_X1 U1092 ( .A(G164), .B(G2078), .ZN(n1003) );
  XNOR2_X1 U1093 ( .A(n1003), .B(KEYINPUT117), .ZN(n1006) );
  XOR2_X1 U1094 ( .A(G2072), .B(n1004), .Z(n1005) );
  NOR2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1096 ( .A(KEYINPUT50), .B(n1007), .ZN(n1026) );
  XOR2_X1 U1097 ( .A(G2090), .B(G162), .Z(n1008) );
  NOR2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1099 ( .A(KEYINPUT51), .B(n1010), .Z(n1011) );
  NAND2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1024) );
  XNOR2_X1 U1101 ( .A(G160), .B(G2084), .ZN(n1013) );
  XNOR2_X1 U1102 ( .A(n1013), .B(KEYINPUT113), .ZN(n1018) );
  NOR2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1104 ( .A(KEYINPUT114), .B(n1016), .Z(n1017) );
  NOR2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1106 ( .A(n1019), .B(KEYINPUT115), .ZN(n1020) );
  NOR2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XOR2_X1 U1108 ( .A(KEYINPUT116), .B(n1022), .Z(n1023) );
  NOR2_X1 U1109 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1110 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1111 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1112 ( .A(KEYINPUT52), .B(n1029), .ZN(n1031) );
  NAND2_X1 U1113 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NAND2_X1 U1114 ( .A1(n1032), .A2(G29), .ZN(n1033) );
  NAND2_X1 U1115 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XNOR2_X1 U1116 ( .A(n1036), .B(n1035), .ZN(G311) );
  XNOR2_X1 U1117 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
endmodule

