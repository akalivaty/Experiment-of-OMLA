//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 1 0 1 1 1 0 1 0 1 0 0 1 1 1 0 0 0 0 1 1 1 1 0 1 1 0 0 0 1 1 1 0 0 0 1 0 1 1 1 1 1 1 1 1 1 1 1 0 0 1 1 0 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:03 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n770, new_n771,
    new_n772, new_n773, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n800, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050;
  INV_X1    g000(.A(G475), .ZN(new_n187));
  INV_X1    g001(.A(G131), .ZN(new_n188));
  INV_X1    g002(.A(G237), .ZN(new_n189));
  INV_X1    g003(.A(G953), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(G214), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT87), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(G143), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT87), .ZN(new_n196));
  NOR2_X1   g010(.A1(G237), .A2(G953), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(G214), .A3(new_n197), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n188), .B1(new_n194), .B2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT17), .ZN(new_n200));
  INV_X1    g014(.A(G140), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G125), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT16), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(KEYINPUT72), .A2(G125), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(new_n201), .ZN(new_n206));
  NAND3_X1  g020(.A1(KEYINPUT72), .A2(G125), .A3(G140), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n204), .B1(new_n208), .B2(new_n203), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G146), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n211), .B(new_n204), .C1(new_n208), .C2(new_n203), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n200), .A2(new_n210), .A3(new_n212), .ZN(new_n213));
  AND3_X1   g027(.A1(new_n194), .A2(new_n198), .A3(new_n188), .ZN(new_n214));
  NOR3_X1   g028(.A1(new_n214), .A2(new_n199), .A3(KEYINPUT17), .ZN(new_n215));
  OR2_X1    g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT93), .ZN(new_n217));
  XNOR2_X1  g031(.A(G113), .B(G122), .ZN(new_n218));
  INV_X1    g032(.A(G104), .ZN(new_n219));
  XNOR2_X1  g033(.A(new_n218), .B(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n196), .B1(G214), .B2(new_n197), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n191), .A2(new_n193), .ZN(new_n222));
  OAI211_X1 g036(.A(KEYINPUT18), .B(G131), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  XNOR2_X1  g037(.A(G125), .B(G140), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(new_n211), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n225), .B1(new_n211), .B2(new_n208), .ZN(new_n226));
  NAND2_X1  g040(.A1(KEYINPUT18), .A2(G131), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n194), .A2(new_n198), .A3(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n223), .A2(new_n226), .A3(new_n228), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n216), .A2(new_n217), .A3(new_n220), .A4(new_n229), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n220), .B(new_n229), .C1(new_n213), .C2(new_n215), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT93), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  AND2_X1   g047(.A1(new_n216), .A2(new_n229), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n233), .B1(new_n220), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G902), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n187), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT20), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n206), .A2(KEYINPUT19), .A3(new_n207), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(KEYINPUT89), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT89), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n206), .A2(new_n242), .A3(KEYINPUT19), .A4(new_n207), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G125), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G140), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT19), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n202), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT90), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT90), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n224), .A2(new_n250), .A3(new_n247), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n244), .A2(new_n252), .A3(new_n211), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT91), .ZN(new_n254));
  OAI21_X1  g068(.A(KEYINPUT88), .B1(new_n214), .B2(new_n199), .ZN(new_n255));
  OAI21_X1  g069(.A(G131), .B1(new_n221), .B2(new_n222), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT88), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n194), .A2(new_n198), .A3(new_n188), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n256), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT91), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n244), .A2(new_n252), .A3(new_n261), .A4(new_n211), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n254), .A2(new_n260), .A3(new_n210), .A4(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n220), .B1(new_n263), .B2(new_n229), .ZN(new_n264));
  AOI22_X1  g078(.A1(new_n264), .A2(KEYINPUT92), .B1(new_n230), .B2(new_n232), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n263), .A2(new_n229), .ZN(new_n266));
  INV_X1    g080(.A(new_n220), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT92), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n265), .A2(new_n270), .ZN(new_n271));
  NOR2_X1   g085(.A1(G475), .A2(G902), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n239), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n272), .ZN(new_n274));
  AOI211_X1 g088(.A(KEYINPUT20), .B(new_n274), .C1(new_n265), .C2(new_n270), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n238), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT94), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n266), .A2(KEYINPUT92), .A3(new_n267), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n233), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n264), .A2(KEYINPUT92), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n272), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(KEYINPUT20), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n271), .A2(new_n239), .A3(new_n272), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n285), .A2(KEYINPUT94), .A3(new_n238), .ZN(new_n286));
  INV_X1    g100(.A(G116), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(G122), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT95), .ZN(new_n289));
  XNOR2_X1  g103(.A(new_n288), .B(new_n289), .ZN(new_n290));
  OR2_X1    g104(.A1(new_n287), .A2(G122), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(G107), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n290), .A2(G107), .A3(new_n291), .ZN(new_n295));
  INV_X1    g109(.A(G134), .ZN(new_n296));
  AND2_X1   g110(.A1(KEYINPUT66), .A2(G128), .ZN(new_n297));
  NOR2_X1   g111(.A1(KEYINPUT66), .A2(G128), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G143), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT13), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n296), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n195), .A2(G128), .ZN(new_n303));
  AND3_X1   g117(.A1(new_n302), .A2(new_n300), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n302), .B1(new_n300), .B2(new_n303), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n294), .B(new_n295), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n291), .A2(KEYINPUT14), .A3(G107), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n294), .A2(new_n295), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n300), .A2(new_n303), .ZN(new_n309));
  XOR2_X1   g123(.A(KEYINPUT96), .B(G134), .Z(new_n310));
  XNOR2_X1  g124(.A(new_n309), .B(new_n310), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n290), .A2(KEYINPUT14), .A3(G107), .A4(new_n291), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n308), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n306), .A2(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT9), .B(G234), .ZN(new_n315));
  INV_X1    g129(.A(G217), .ZN(new_n316));
  NOR3_X1   g130(.A1(new_n315), .A2(new_n316), .A3(G953), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n314), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n306), .A2(new_n313), .A3(new_n317), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(new_n236), .ZN(new_n322));
  INV_X1    g136(.A(G478), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n323), .A2(KEYINPUT15), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  OAI211_X1 g139(.A(new_n321), .B(new_n236), .C1(KEYINPUT15), .C2(new_n323), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AOI211_X1 g141(.A(new_n236), .B(new_n190), .C1(G234), .C2(G237), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT21), .B(G898), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  OR2_X1    g144(.A1(KEYINPUT97), .A2(G952), .ZN(new_n331));
  NAND2_X1  g145(.A1(KEYINPUT97), .A2(G952), .ZN(new_n332));
  AOI21_X1  g146(.A(G953), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(G234), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n333), .B1(new_n334), .B2(new_n189), .ZN(new_n335));
  AND2_X1   g149(.A1(new_n330), .A2(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n327), .A2(new_n336), .ZN(new_n337));
  AND3_X1   g151(.A1(new_n278), .A2(new_n286), .A3(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(G221), .ZN(new_n339));
  INV_X1    g153(.A(new_n315), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n339), .B1(new_n340), .B2(new_n236), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n341), .B(KEYINPUT77), .ZN(new_n342));
  OAI21_X1  g156(.A(G214), .B1(G237), .B2(G902), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n211), .A2(G143), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n195), .A2(G146), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT1), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n347), .B1(G143), .B2(new_n211), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n346), .B1(new_n299), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(G128), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n350), .A2(KEYINPUT1), .ZN(new_n351));
  AND3_X1   g165(.A1(new_n195), .A2(KEYINPUT64), .A3(G146), .ZN(new_n352));
  AOI21_X1  g166(.A(KEYINPUT64), .B1(new_n195), .B2(G146), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n344), .B(new_n351), .C1(new_n352), .C2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n349), .A2(new_n354), .A3(new_n245), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n195), .A2(G146), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT64), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n357), .B1(new_n211), .B2(G143), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n195), .A2(KEYINPUT64), .A3(G146), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n356), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  AND2_X1   g174(.A1(KEYINPUT0), .A2(G128), .ZN(new_n361));
  NOR2_X1   g175(.A1(KEYINPUT0), .A2(G128), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI22_X1  g177(.A1(new_n360), .A2(new_n361), .B1(new_n363), .B2(new_n346), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n355), .B1(new_n364), .B2(new_n245), .ZN(new_n365));
  OAI21_X1  g179(.A(KEYINPUT86), .B1(new_n364), .B2(new_n245), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT7), .ZN(new_n367));
  INV_X1    g181(.A(G224), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n368), .A2(G953), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n365), .B(new_n366), .C1(new_n367), .C2(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n369), .A2(new_n367), .ZN(new_n371));
  OAI221_X1 g185(.A(new_n355), .B1(KEYINPUT86), .B2(new_n371), .C1(new_n364), .C2(new_n245), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n219), .A2(G107), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n219), .A2(G107), .ZN(new_n376));
  OAI21_X1  g190(.A(G101), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(KEYINPUT3), .B1(new_n219), .B2(G107), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT3), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n379), .A2(new_n293), .A3(G104), .ZN(new_n380));
  INV_X1    g194(.A(G101), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n378), .A2(new_n380), .A3(new_n381), .A4(new_n374), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n377), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT67), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n384), .B1(new_n287), .B2(G119), .ZN(new_n385));
  INV_X1    g199(.A(G119), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(KEYINPUT67), .A3(G116), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n287), .A2(G119), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n385), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(KEYINPUT2), .B(G113), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  OR2_X1    g205(.A1(new_n383), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT84), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT5), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n389), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n394), .A2(new_n386), .A3(G116), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(KEYINPUT83), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT83), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n398), .A2(new_n394), .A3(new_n386), .A4(G116), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n397), .A2(G113), .A3(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n393), .B1(new_n395), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n400), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n402), .B(KEYINPUT84), .C1(new_n394), .C2(new_n389), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n392), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  XOR2_X1   g218(.A(new_n389), .B(new_n390), .Z(new_n405));
  NAND3_X1  g219(.A1(new_n378), .A2(new_n380), .A3(new_n374), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(KEYINPUT78), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT78), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n378), .A2(new_n380), .A3(new_n408), .A4(new_n374), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n407), .A2(G101), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n382), .A2(KEYINPUT4), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n407), .A2(KEYINPUT4), .A3(G101), .A4(new_n409), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n405), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n404), .A2(new_n414), .ZN(new_n415));
  XNOR2_X1  g229(.A(G110), .B(G122), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n373), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT85), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n395), .B1(new_n418), .B2(new_n400), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n419), .B1(new_n418), .B2(new_n400), .ZN(new_n420));
  INV_X1    g234(.A(new_n392), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n383), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n391), .B1(new_n403), .B2(new_n401), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n422), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n416), .B(KEYINPUT8), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(G902), .B1(new_n417), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n403), .A2(new_n401), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n421), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n412), .A2(new_n413), .ZN(new_n431));
  INV_X1    g245(.A(new_n405), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n430), .A2(new_n433), .A3(new_n416), .ZN(new_n434));
  INV_X1    g248(.A(new_n416), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n435), .B1(new_n404), .B2(new_n414), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n434), .A2(new_n436), .A3(KEYINPUT6), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT6), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n438), .B(new_n435), .C1(new_n404), .C2(new_n414), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n365), .B(new_n369), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n437), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(G210), .B1(G237), .B2(G902), .ZN(new_n442));
  AND3_X1   g256(.A1(new_n428), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n442), .B1(new_n428), .B2(new_n441), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n343), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(G469), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT82), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT79), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n354), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n350), .B1(new_n344), .B2(KEYINPUT1), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n360), .A2(new_n450), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n358), .A2(new_n359), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n453), .A2(KEYINPUT79), .A3(new_n344), .A4(new_n351), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n454), .A2(new_n377), .A3(new_n382), .ZN(new_n455));
  NOR3_X1   g269(.A1(new_n452), .A2(KEYINPUT80), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT80), .ZN(new_n457));
  AND3_X1   g271(.A1(new_n454), .A2(new_n377), .A3(new_n382), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n354), .B(new_n448), .C1(new_n360), .C2(new_n450), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n457), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n349), .A2(new_n354), .ZN(new_n461));
  OAI22_X1  g275(.A1(new_n456), .A2(new_n460), .B1(new_n461), .B2(new_n423), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT11), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n463), .B1(new_n296), .B2(G137), .ZN(new_n464));
  INV_X1    g278(.A(G137), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n465), .A2(KEYINPUT11), .A3(G134), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n296), .A2(G137), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n464), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(G131), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n464), .A2(new_n466), .A3(new_n188), .A4(new_n467), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(KEYINPUT12), .B1(new_n462), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n423), .A2(new_n461), .ZN(new_n473));
  OAI21_X1  g287(.A(KEYINPUT80), .B1(new_n452), .B2(new_n455), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n458), .A2(new_n457), .A3(new_n459), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT12), .ZN(new_n477));
  INV_X1    g291(.A(new_n471), .ZN(new_n478));
  NOR3_X1   g292(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n472), .A2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT10), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n481), .B1(new_n456), .B2(new_n460), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n423), .A2(KEYINPUT10), .A3(new_n461), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n484), .B1(new_n431), .B2(new_n364), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n482), .A2(new_n485), .A3(new_n478), .ZN(new_n486));
  XNOR2_X1  g300(.A(G110), .B(G140), .ZN(new_n487));
  AND2_X1   g301(.A1(new_n190), .A2(G227), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n487), .B(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n447), .B1(new_n480), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n462), .A2(KEYINPUT12), .A3(new_n471), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n477), .B1(new_n476), .B2(new_n478), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n495), .A2(KEYINPUT82), .A3(new_n486), .A4(new_n490), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n431), .A2(new_n364), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(new_n483), .ZN(new_n499));
  AOI21_X1  g313(.A(KEYINPUT10), .B1(new_n474), .B2(new_n475), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n471), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(KEYINPUT81), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT81), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n503), .B(new_n471), .C1(new_n499), .C2(new_n500), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n490), .B1(new_n505), .B2(new_n486), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n446), .B(new_n236), .C1(new_n497), .C2(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n491), .B1(new_n502), .B2(new_n504), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n490), .B1(new_n495), .B2(new_n486), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(G469), .B1(new_n510), .B2(G902), .ZN(new_n511));
  AOI211_X1 g325(.A(new_n342), .B(new_n445), .C1(new_n507), .C2(new_n511), .ZN(new_n512));
  AND2_X1   g326(.A1(new_n338), .A2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT71), .ZN(new_n514));
  AND2_X1   g328(.A1(new_n514), .A2(KEYINPUT23), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n514), .A2(KEYINPUT23), .ZN(new_n516));
  OAI22_X1  g330(.A1(new_n515), .A2(new_n516), .B1(new_n386), .B2(G128), .ZN(new_n517));
  INV_X1    g331(.A(new_n298), .ZN(new_n518));
  NAND2_X1  g332(.A1(KEYINPUT66), .A2(G128), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n518), .A2(KEYINPUT23), .A3(G119), .A4(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(G110), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n350), .A2(G119), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n517), .A2(new_n520), .A3(new_n521), .A4(new_n523), .ZN(new_n524));
  XNOR2_X1  g338(.A(KEYINPUT24), .B(G110), .ZN(new_n525));
  NOR3_X1   g339(.A1(new_n297), .A2(new_n298), .A3(new_n386), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n525), .B1(new_n526), .B2(new_n522), .ZN(new_n527));
  AND3_X1   g341(.A1(new_n524), .A2(KEYINPUT74), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(KEYINPUT74), .B1(new_n524), .B2(new_n527), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n210), .B(new_n225), .C1(new_n528), .C2(new_n529), .ZN(new_n530));
  NOR3_X1   g344(.A1(new_n526), .A2(new_n522), .A3(new_n525), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n517), .A2(new_n523), .A3(new_n520), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n531), .B1(G110), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n210), .A2(new_n212), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT73), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n535), .B1(new_n533), .B2(new_n534), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n530), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  XOR2_X1   g352(.A(KEYINPUT22), .B(G137), .Z(new_n539));
  INV_X1    g353(.A(KEYINPUT75), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g355(.A(KEYINPUT22), .B(G137), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(KEYINPUT75), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT76), .ZN(new_n545));
  NOR3_X1   g359(.A1(new_n339), .A2(new_n334), .A3(G953), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT76), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n541), .A2(new_n547), .A3(new_n543), .ZN(new_n548));
  AND3_X1   g362(.A1(new_n545), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n546), .B1(new_n545), .B2(new_n548), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n538), .A2(new_n552), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n551), .B(new_n530), .C1(new_n536), .C2(new_n537), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n553), .A2(new_n236), .A3(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT25), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n553), .A2(KEYINPUT25), .A3(new_n554), .A4(new_n236), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n316), .B1(G234), .B2(new_n236), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n553), .A2(new_n554), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n560), .A2(G902), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT68), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n471), .A2(new_n364), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n296), .A2(G137), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n465), .A2(G134), .ZN(new_n570));
  OAI21_X1  g384(.A(G131), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  AND2_X1   g385(.A1(new_n470), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n461), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n405), .A2(new_n568), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n197), .A2(G210), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n575), .B(KEYINPUT27), .ZN(new_n576));
  XNOR2_X1  g390(.A(KEYINPUT26), .B(G101), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n576), .B(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT30), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n581), .B1(new_n568), .B2(new_n573), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n470), .A2(new_n571), .ZN(new_n583));
  AOI22_X1  g397(.A1(new_n583), .A2(KEYINPUT65), .B1(new_n349), .B2(new_n354), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT65), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n470), .A2(new_n571), .A3(new_n585), .ZN(new_n586));
  AOI22_X1  g400(.A1(new_n584), .A2(new_n586), .B1(new_n471), .B2(new_n364), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n582), .B1(new_n581), .B2(new_n587), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n567), .B(new_n580), .C1(new_n588), .C2(new_n405), .ZN(new_n589));
  AND2_X1   g403(.A1(new_n471), .A2(new_n364), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n583), .B1(new_n354), .B2(new_n349), .ZN(new_n591));
  OAI21_X1  g405(.A(KEYINPUT30), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n583), .A2(KEYINPUT65), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n593), .A2(new_n461), .A3(new_n586), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n594), .A2(new_n581), .A3(new_n568), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n405), .B1(new_n592), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(KEYINPUT68), .B1(new_n596), .B2(new_n579), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n589), .A2(new_n597), .A3(KEYINPUT31), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n592), .A2(new_n595), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n579), .B1(new_n599), .B2(new_n432), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT31), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT28), .ZN(new_n602));
  AOI22_X1  g416(.A1(new_n471), .A2(new_n364), .B1(new_n461), .B2(new_n572), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n602), .B1(new_n603), .B2(new_n405), .ZN(new_n604));
  AND4_X1   g418(.A1(new_n602), .A2(new_n405), .A3(new_n568), .A4(new_n573), .ZN(new_n605));
  OAI22_X1  g419(.A1(new_n604), .A2(new_n605), .B1(new_n405), .B2(new_n587), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT69), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n578), .B(new_n607), .ZN(new_n608));
  AOI22_X1  g422(.A1(new_n600), .A2(new_n601), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n598), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(G472), .A2(G902), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(KEYINPUT70), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT32), .ZN(new_n614));
  INV_X1    g428(.A(new_n611), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n615), .B1(new_n598), .B2(new_n609), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT70), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n613), .A2(new_n614), .A3(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n604), .A2(new_n605), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n603), .A2(new_n405), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n578), .A2(KEYINPUT29), .ZN(new_n623));
  AOI21_X1  g437(.A(G902), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n574), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n596), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n626), .A2(new_n578), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT29), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n628), .B1(new_n606), .B2(new_n608), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n624), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  AOI22_X1  g444(.A1(new_n616), .A2(KEYINPUT32), .B1(new_n630), .B2(G472), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n566), .B1(new_n619), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n513), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(G101), .ZN(G3));
  AOI21_X1  g448(.A(new_n342), .B1(new_n507), .B2(new_n511), .ZN(new_n635));
  INV_X1    g449(.A(new_n566), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n610), .A2(new_n236), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(G472), .ZN(new_n638));
  AND3_X1   g452(.A1(new_n613), .A2(new_n638), .A3(new_n618), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n635), .A2(new_n636), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(KEYINPUT98), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT98), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n635), .A2(new_n642), .A3(new_n636), .A4(new_n639), .ZN(new_n643));
  AND2_X1   g457(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n278), .A2(new_n286), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n317), .B1(new_n306), .B2(new_n313), .ZN(new_n646));
  OAI211_X1 g460(.A(new_n321), .B(KEYINPUT33), .C1(KEYINPUT99), .C2(new_n646), .ZN(new_n647));
  OAI21_X1  g461(.A(KEYINPUT33), .B1(new_n646), .B2(KEYINPUT99), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n648), .A2(new_n320), .A3(new_n319), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n647), .A2(new_n649), .A3(G478), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n323), .A2(new_n236), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  OAI211_X1 g466(.A(new_n650), .B(new_n652), .C1(G478), .C2(new_n322), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n445), .A2(new_n336), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n645), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(KEYINPUT100), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n653), .B1(new_n278), .B2(new_n286), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT100), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n658), .A2(new_n659), .A3(new_n655), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n644), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT101), .ZN(new_n663));
  XNOR2_X1  g477(.A(KEYINPUT34), .B(G104), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G6));
  INV_X1    g479(.A(new_n445), .ZN(new_n666));
  INV_X1    g480(.A(new_n336), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g482(.A(KEYINPUT102), .B1(new_n273), .B2(new_n275), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT102), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n283), .A2(new_n670), .A3(new_n284), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n669), .A2(new_n671), .A3(new_n238), .A4(new_n327), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n644), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT35), .B(G107), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G9));
  OR3_X1    g490(.A1(new_n538), .A2(KEYINPUT36), .A3(new_n552), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n538), .B1(new_n552), .B2(KEYINPUT36), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n564), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n561), .A2(new_n681), .ZN(new_n682));
  AND4_X1   g496(.A1(new_n613), .A2(new_n682), .A3(new_n618), .A4(new_n638), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n513), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g498(.A(KEYINPUT37), .B(G110), .Z(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G12));
  OR2_X1    g500(.A1(KEYINPUT103), .A2(G900), .ZN(new_n687));
  NAND2_X1  g501(.A1(KEYINPUT103), .A2(G900), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n328), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n335), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n672), .A2(new_n691), .ZN(new_n692));
  AOI22_X1  g506(.A1(new_n560), .A2(new_n559), .B1(new_n680), .B2(new_n564), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n693), .B1(new_n619), .B2(new_n631), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n512), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT104), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n512), .A2(new_n692), .A3(KEYINPUT104), .A4(new_n694), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G128), .ZN(G30));
  NOR2_X1   g514(.A1(new_n443), .A2(new_n444), .ZN(new_n701));
  OR2_X1    g515(.A1(new_n701), .A2(KEYINPUT38), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(KEYINPUT38), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  AND4_X1   g518(.A1(new_n343), .A2(new_n704), .A3(new_n327), .A4(new_n693), .ZN(new_n705));
  AND2_X1   g519(.A1(new_n705), .A2(new_n645), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n690), .B(KEYINPUT39), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n635), .A2(new_n707), .ZN(new_n708));
  OR2_X1    g522(.A1(new_n708), .A2(KEYINPUT40), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(KEYINPUT40), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n608), .B1(new_n625), .B2(new_n621), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT105), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI211_X1 g527(.A(new_n608), .B(KEYINPUT105), .C1(new_n625), .C2(new_n621), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n589), .A2(new_n597), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n236), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AOI22_X1  g531(.A1(new_n717), .A2(G472), .B1(new_n616), .B2(KEYINPUT32), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n619), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n706), .A2(new_n709), .A3(new_n710), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G143), .ZN(G45));
  AOI211_X1 g535(.A(new_n653), .B(new_n691), .C1(new_n278), .C2(new_n286), .ZN(new_n722));
  AND3_X1   g536(.A1(new_n722), .A2(new_n512), .A3(new_n694), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(new_n211), .ZN(G48));
  INV_X1    g538(.A(new_n507), .ZN(new_n725));
  INV_X1    g539(.A(new_n486), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n726), .B1(new_n502), .B2(new_n504), .ZN(new_n727));
  OAI211_X1 g541(.A(new_n492), .B(new_n496), .C1(new_n727), .C2(new_n490), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n446), .B1(new_n728), .B2(new_n236), .ZN(new_n729));
  NOR3_X1   g543(.A1(new_n725), .A2(new_n729), .A3(new_n341), .ZN(new_n730));
  AND2_X1   g544(.A1(new_n730), .A2(new_n632), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n661), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(KEYINPUT41), .B(G113), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n732), .B(new_n733), .ZN(G15));
  NAND3_X1  g548(.A1(new_n673), .A2(new_n730), .A3(new_n632), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G116), .ZN(G18));
  AOI21_X1  g550(.A(KEYINPUT94), .B1(new_n285), .B2(new_n238), .ZN(new_n737));
  AOI211_X1 g551(.A(new_n277), .B(new_n237), .C1(new_n283), .C2(new_n284), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n739), .A2(new_n694), .A3(new_n337), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n725), .A2(new_n729), .ZN(new_n741));
  INV_X1    g555(.A(new_n341), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n741), .A2(KEYINPUT106), .A3(new_n742), .A4(new_n666), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n236), .B1(new_n497), .B2(new_n506), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(G469), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n745), .A2(new_n507), .A3(new_n742), .A4(new_n666), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT106), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n740), .B1(new_n743), .B2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(new_n386), .ZN(G21));
  OAI211_X1 g564(.A(new_n327), .B(new_n343), .C1(new_n443), .C2(new_n444), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n752), .B1(new_n737), .B2(new_n738), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT108), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n645), .A2(KEYINPUT108), .A3(new_n752), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n745), .A2(new_n507), .A3(new_n742), .A4(new_n667), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n600), .A2(new_n601), .ZN(new_n759));
  AND2_X1   g573(.A1(new_n622), .A2(KEYINPUT107), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n608), .B1(new_n622), .B2(KEYINPUT107), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(new_n598), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n611), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n764), .A2(new_n638), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n636), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n758), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n757), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G122), .ZN(G24));
  AND2_X1   g583(.A1(new_n765), .A2(new_n682), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n722), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n743), .A2(new_n748), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G125), .ZN(G27));
  INV_X1    g588(.A(new_n444), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n428), .A2(new_n441), .A3(new_n442), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n775), .A2(new_n343), .A3(new_n776), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n777), .A2(new_n341), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(G469), .A2(G902), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(KEYINPUT109), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n782), .B1(new_n510), .B2(G469), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n507), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(KEYINPUT110), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT110), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n507), .A2(new_n783), .A3(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n779), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT42), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n788), .A2(new_n789), .A3(new_n632), .A4(new_n722), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n507), .A2(new_n786), .A3(new_n783), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n786), .B1(new_n507), .B2(new_n783), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n778), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n612), .A2(new_n614), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n566), .B1(new_n631), .B2(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n645), .A2(new_n795), .A3(new_n654), .A4(new_n690), .ZN(new_n796));
  OAI21_X1  g610(.A(KEYINPUT42), .B1(new_n793), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n790), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(new_n188), .ZN(G33));
  NAND2_X1  g613(.A1(new_n785), .A2(new_n787), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n800), .A2(new_n632), .A3(new_n692), .A4(new_n778), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G134), .ZN(G36));
  NAND2_X1  g616(.A1(new_n739), .A2(new_n654), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n803), .A2(KEYINPUT113), .A3(KEYINPUT43), .ZN(new_n804));
  AOI21_X1  g618(.A(KEYINPUT43), .B1(new_n803), .B2(KEYINPUT113), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n639), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n806), .A2(new_n807), .A3(new_n682), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(KEYINPUT44), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n510), .A2(KEYINPUT45), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT45), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n811), .B1(new_n508), .B2(new_n509), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n810), .A2(G469), .A3(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n813), .A2(KEYINPUT46), .A3(new_n781), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n507), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(KEYINPUT111), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT111), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n814), .A2(new_n817), .A3(new_n507), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n813), .A2(new_n781), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT46), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n816), .A2(new_n818), .A3(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n822), .A2(new_n341), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT112), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n823), .A2(new_n824), .A3(new_n707), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n823), .A2(new_n707), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(KEYINPUT112), .ZN(new_n827));
  XOR2_X1   g641(.A(new_n777), .B(KEYINPUT114), .Z(new_n828));
  NAND4_X1  g642(.A1(new_n809), .A2(new_n825), .A3(new_n827), .A4(new_n828), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(G137), .ZN(G39));
  INV_X1    g644(.A(KEYINPUT47), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n831), .B1(new_n822), .B2(new_n341), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n816), .A2(new_n818), .A3(new_n821), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n833), .A2(KEYINPUT47), .A3(new_n742), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(new_n777), .ZN(new_n836));
  AND4_X1   g650(.A1(new_n619), .A2(new_n836), .A3(new_n631), .A4(new_n566), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n835), .A2(new_n722), .A3(new_n837), .ZN(new_n838));
  XNOR2_X1  g652(.A(new_n838), .B(G140), .ZN(G42));
  XNOR2_X1  g653(.A(new_n741), .B(KEYINPUT49), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n719), .A2(new_n566), .ZN(new_n841));
  INV_X1    g655(.A(new_n342), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n654), .A2(new_n842), .A3(new_n343), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n704), .A2(new_n645), .A3(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n840), .A2(new_n841), .A3(new_n844), .ZN(new_n845));
  OR2_X1    g659(.A1(G952), .A2(G953), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n766), .A2(new_n335), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n804), .A2(new_n805), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n741), .A2(new_n742), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n850), .A2(new_n343), .A3(new_n704), .ZN(new_n851));
  AOI21_X1  g665(.A(KEYINPUT50), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n803), .A2(KEYINPUT113), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT43), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n803), .A2(KEYINPUT113), .A3(KEYINPUT43), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n855), .A2(new_n851), .A3(new_n856), .A4(new_n847), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT50), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g673(.A(KEYINPUT116), .B1(new_n852), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n741), .A2(new_n342), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n832), .A2(new_n834), .A3(new_n861), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n849), .A2(new_n828), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NOR4_X1   g678(.A1(new_n779), .A2(new_n725), .A3(new_n729), .A4(new_n335), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n806), .A2(new_n770), .A3(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n865), .A2(new_n739), .A3(new_n653), .A4(new_n841), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n849), .A2(KEYINPUT50), .A3(new_n851), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT116), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n857), .A2(new_n858), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n860), .A2(new_n864), .A3(new_n869), .A4(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT51), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n865), .A2(new_n658), .A3(new_n841), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(new_n333), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n878), .B1(new_n849), .B2(new_n772), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n855), .A2(new_n795), .A3(new_n856), .A4(new_n865), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n880), .A2(KEYINPUT48), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n880), .A2(KEYINPUT48), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n879), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n868), .B1(new_n862), .B2(new_n863), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n875), .B1(new_n870), .B2(new_n872), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n876), .A2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT53), .ZN(new_n888));
  AOI21_X1  g702(.A(KEYINPUT108), .B1(new_n645), .B2(new_n752), .ZN(new_n889));
  AOI211_X1 g703(.A(new_n754), .B(new_n751), .C1(new_n278), .C2(new_n286), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AND4_X1   g705(.A1(new_n561), .A2(new_n681), .A3(new_n742), .A4(new_n690), .ZN(new_n892));
  OAI211_X1 g706(.A(new_n719), .B(new_n892), .C1(new_n791), .C2(new_n792), .ZN(new_n893));
  OAI21_X1  g707(.A(KEYINPUT115), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n719), .A2(new_n892), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n895), .B1(new_n787), .B2(new_n785), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT115), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n757), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n894), .A2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT52), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n723), .B1(new_n772), .B2(new_n771), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n899), .A2(new_n900), .A3(new_n901), .A4(new_n699), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n338), .B(new_n512), .C1(new_n683), .C2(new_n632), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n903), .A2(new_n735), .ZN(new_n904));
  INV_X1    g718(.A(new_n740), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n772), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n904), .A2(new_n906), .A3(new_n768), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n739), .A2(new_n327), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n645), .A2(new_n654), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n668), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n910), .A2(new_n643), .A3(new_n641), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n732), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n907), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n800), .A2(new_n722), .A3(new_n770), .A4(new_n778), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n669), .A2(new_n238), .A3(new_n671), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n777), .A2(new_n327), .A3(new_n691), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n694), .A2(new_n635), .A3(new_n915), .A4(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n914), .A2(new_n801), .A3(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n798), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n902), .A2(new_n913), .A3(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(new_n723), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n699), .A2(new_n773), .A3(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n900), .B1(new_n923), .B2(new_n899), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n888), .B1(new_n920), .B2(new_n924), .ZN(new_n925));
  AOI22_X1  g739(.A1(new_n772), .A2(new_n905), .B1(new_n757), .B2(new_n767), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n926), .A2(new_n732), .A3(new_n904), .A4(new_n911), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n801), .A2(new_n917), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n928), .A2(new_n797), .A3(new_n790), .A4(new_n914), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n757), .A2(new_n896), .A3(new_n897), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n897), .B1(new_n757), .B2(new_n896), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(KEYINPUT52), .B1(new_n933), .B2(new_n922), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n930), .A2(new_n934), .A3(KEYINPUT53), .A4(new_n902), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n925), .A2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT54), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n925), .A2(KEYINPUT54), .A3(new_n935), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n887), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT117), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n846), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AOI211_X1 g756(.A(KEYINPUT117), .B(new_n887), .C1(new_n938), .C2(new_n939), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n845), .B1(new_n942), .B2(new_n943), .ZN(G75));
  AOI21_X1  g758(.A(new_n236), .B1(new_n925), .B2(new_n935), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(G210), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT56), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n437), .A2(new_n439), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(new_n440), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT55), .Z(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(KEYINPUT119), .Z(new_n951));
  NAND3_X1  g765(.A1(new_n946), .A2(new_n947), .A3(new_n951), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n190), .A2(G952), .ZN(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(KEYINPUT56), .B1(new_n945), .B2(G210), .ZN(new_n956));
  INV_X1    g770(.A(new_n950), .ZN(new_n957));
  OAI21_X1  g771(.A(KEYINPUT118), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n946), .A2(new_n947), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT118), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n959), .A2(new_n960), .A3(new_n950), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n955), .B1(new_n958), .B2(new_n961), .ZN(G51));
  XOR2_X1   g776(.A(new_n781), .B(KEYINPUT57), .Z(new_n963));
  NAND3_X1  g777(.A1(new_n938), .A2(new_n939), .A3(new_n963), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n728), .B(KEYINPUT120), .Z(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(new_n945), .ZN(new_n967));
  OR2_X1    g781(.A1(new_n967), .A2(new_n813), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n953), .B1(new_n966), .B2(new_n968), .ZN(G54));
  NAND3_X1  g783(.A1(new_n945), .A2(KEYINPUT58), .A3(G475), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n970), .A2(new_n270), .A3(new_n265), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n945), .A2(KEYINPUT58), .A3(G475), .A4(new_n271), .ZN(new_n972));
  AND3_X1   g786(.A1(new_n971), .A2(new_n954), .A3(new_n972), .ZN(G60));
  XNOR2_X1  g787(.A(new_n651), .B(KEYINPUT121), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n974), .B(KEYINPUT59), .Z(new_n975));
  NAND3_X1  g789(.A1(new_n938), .A2(new_n939), .A3(new_n975), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n647), .A2(new_n649), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n976), .A2(new_n977), .ZN(new_n979));
  NOR3_X1   g793(.A1(new_n978), .A2(new_n979), .A3(new_n953), .ZN(G63));
  XOR2_X1   g794(.A(KEYINPUT122), .B(KEYINPUT61), .Z(new_n981));
  NAND2_X1  g795(.A1(G217), .A2(G902), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n982), .B(KEYINPUT123), .Z(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(KEYINPUT60), .Z(new_n984));
  OAI21_X1  g798(.A(new_n900), .B1(new_n931), .B2(new_n932), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n985), .A2(new_n922), .ZN(new_n986));
  AOI211_X1 g800(.A(new_n766), .B(new_n758), .C1(new_n755), .C2(new_n756), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n903), .A2(new_n735), .ZN(new_n988));
  NOR3_X1   g802(.A1(new_n987), .A2(new_n988), .A3(new_n749), .ZN(new_n989));
  AOI22_X1  g803(.A1(new_n644), .A2(new_n910), .B1(new_n661), .B2(new_n731), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n919), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n986), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(KEYINPUT53), .B1(new_n992), .B2(new_n934), .ZN(new_n993));
  INV_X1    g807(.A(new_n935), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n984), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n954), .B1(new_n995), .B2(new_n679), .ZN(new_n996));
  INV_X1    g810(.A(new_n984), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n997), .B1(new_n925), .B2(new_n935), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n998), .A2(new_n563), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n981), .B1(new_n996), .B2(new_n999), .ZN(new_n1000));
  OAI21_X1  g814(.A(KEYINPUT61), .B1(new_n998), .B2(new_n563), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT124), .ZN(new_n1002));
  NOR3_X1   g816(.A1(new_n996), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(KEYINPUT61), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1004), .B1(new_n995), .B2(new_n562), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n953), .B1(new_n998), .B2(new_n680), .ZN(new_n1006));
  AOI21_X1  g820(.A(KEYINPUT124), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1000), .B1(new_n1003), .B2(new_n1007), .ZN(G66));
  OAI21_X1  g822(.A(G953), .B1(new_n329), .B2(new_n368), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n1009), .B(KEYINPUT125), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1010), .B1(new_n913), .B2(G953), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n948), .B1(G898), .B2(new_n190), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1011), .B(new_n1012), .ZN(G69));
  AOI21_X1  g827(.A(new_n190), .B1(G227), .B2(G900), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n244), .A2(new_n252), .ZN(new_n1015));
  XOR2_X1   g829(.A(new_n1015), .B(KEYINPUT126), .Z(new_n1016));
  XNOR2_X1  g830(.A(new_n599), .B(new_n1016), .ZN(new_n1017));
  NAND2_X1  g831(.A1(G900), .A2(G953), .ZN(new_n1018));
  NAND4_X1  g832(.A1(new_n827), .A2(new_n757), .A3(new_n795), .A4(new_n825), .ZN(new_n1019));
  INV_X1    g833(.A(new_n801), .ZN(new_n1020));
  NOR3_X1   g834(.A1(new_n922), .A2(new_n798), .A3(new_n1020), .ZN(new_n1021));
  NAND4_X1  g835(.A1(new_n829), .A2(new_n838), .A3(new_n1019), .A4(new_n1021), .ZN(new_n1022));
  OAI211_X1 g836(.A(new_n1017), .B(new_n1018), .C1(new_n1022), .C2(G953), .ZN(new_n1023));
  INV_X1    g837(.A(new_n1023), .ZN(new_n1024));
  INV_X1    g838(.A(KEYINPUT62), .ZN(new_n1025));
  INV_X1    g839(.A(new_n720), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1025), .B1(new_n1026), .B2(new_n922), .ZN(new_n1027));
  NAND3_X1  g841(.A1(new_n923), .A2(new_n720), .A3(KEYINPUT62), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n908), .A2(new_n909), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n708), .A2(new_n777), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n1030), .A2(new_n1031), .A3(new_n632), .ZN(new_n1032));
  NAND4_X1  g846(.A1(new_n829), .A2(new_n838), .A3(new_n1029), .A4(new_n1032), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n1017), .B1(new_n1033), .B2(new_n190), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n1014), .B1(new_n1024), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g849(.A(new_n1014), .ZN(new_n1036));
  AND2_X1   g850(.A1(new_n1033), .A2(new_n190), .ZN(new_n1037));
  OAI211_X1 g851(.A(new_n1023), .B(new_n1036), .C1(new_n1037), .C2(new_n1017), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1035), .A2(new_n1038), .ZN(G72));
  NAND2_X1  g853(.A1(G472), .A2(G902), .ZN(new_n1040));
  XOR2_X1   g854(.A(new_n1040), .B(KEYINPUT63), .Z(new_n1041));
  OAI21_X1  g855(.A(new_n1041), .B1(new_n1033), .B2(new_n927), .ZN(new_n1042));
  INV_X1    g856(.A(new_n626), .ZN(new_n1043));
  NAND3_X1  g857(.A1(new_n1042), .A2(new_n578), .A3(new_n1043), .ZN(new_n1044));
  OAI21_X1  g858(.A(new_n1041), .B1(new_n1022), .B2(new_n927), .ZN(new_n1045));
  INV_X1    g859(.A(new_n578), .ZN(new_n1046));
  NAND3_X1  g860(.A1(new_n1045), .A2(new_n1046), .A3(new_n626), .ZN(new_n1047));
  OAI21_X1  g861(.A(new_n1041), .B1(new_n716), .B2(new_n627), .ZN(new_n1048));
  XOR2_X1   g862(.A(new_n1048), .B(KEYINPUT127), .Z(new_n1049));
  AOI21_X1  g863(.A(new_n953), .B1(new_n936), .B2(new_n1049), .ZN(new_n1050));
  AND3_X1   g864(.A1(new_n1044), .A2(new_n1047), .A3(new_n1050), .ZN(G57));
endmodule


