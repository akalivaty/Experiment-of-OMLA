//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 0 1 0 1 1 0 0 0 1 0 0 1 1 0 0 0 1 1 0 0 1 1 1 1 1 0 0 0 0 0 1 1 0 0 1 0 1 1 0 0 0 0 1 0 0 1 1 1 0 1 1 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n768, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n867, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n968, new_n969,
    new_n970, new_n971, new_n973, new_n974, new_n975, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n991, new_n992, new_n993, new_n994,
    new_n996, new_n997;
  INV_X1    g000(.A(KEYINPUT3), .ZN(new_n202));
  XNOR2_X1  g001(.A(G197gat), .B(G204gat), .ZN(new_n203));
  INV_X1    g002(.A(G211gat), .ZN(new_n204));
  INV_X1    g003(.A(G218gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n203), .B1(KEYINPUT22), .B2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G211gat), .B(G218gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n207), .B(new_n208), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n202), .B1(new_n209), .B2(KEYINPUT29), .ZN(new_n210));
  INV_X1    g009(.A(G141gat), .ZN(new_n211));
  OAI21_X1  g010(.A(KEYINPUT76), .B1(new_n211), .B2(G148gat), .ZN(new_n212));
  OR3_X1    g011(.A1(new_n211), .A2(KEYINPUT76), .A3(G148gat), .ZN(new_n213));
  XOR2_X1   g012(.A(KEYINPUT75), .B(G141gat), .Z(new_n214));
  INV_X1    g013(.A(G148gat), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n212), .B(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(G155gat), .A2(G162gat), .ZN(new_n217));
  OR2_X1    g016(.A1(G155gat), .A2(G162gat), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n217), .B1(new_n218), .B2(KEYINPUT2), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n216), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(G141gat), .B(G148gat), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n217), .B(new_n218), .C1(new_n221), .C2(KEYINPUT2), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n210), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n209), .B(KEYINPUT72), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n220), .A2(new_n202), .A3(new_n222), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT29), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n224), .B1(new_n225), .B2(new_n229), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n230), .A2(G228gat), .A3(G233gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT81), .ZN(new_n232));
  INV_X1    g031(.A(new_n209), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n232), .B1(new_n229), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G228gat), .A2(G233gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n228), .A2(KEYINPUT81), .A3(new_n209), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n234), .A2(new_n235), .A3(new_n224), .A4(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT31), .B(G50gat), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  AND3_X1   g038(.A1(new_n231), .A2(new_n237), .A3(new_n239), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n239), .B1(new_n231), .B2(new_n237), .ZN(new_n241));
  XNOR2_X1  g040(.A(G78gat), .B(G106gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n242), .B(G22gat), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  OR3_X1    g043(.A1(new_n240), .A2(new_n241), .A3(new_n244), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n244), .B1(new_n240), .B2(new_n241), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(G226gat), .ZN(new_n249));
  INV_X1    g048(.A(G233gat), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(G183gat), .A2(G190gat), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(G169gat), .ZN(new_n255));
  INV_X1    g054(.A(G176gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NOR2_X1   g056(.A1(G169gat), .A2(G176gat), .ZN(new_n258));
  NOR3_X1   g057(.A1(new_n257), .A2(KEYINPUT26), .A3(new_n258), .ZN(new_n259));
  AOI211_X1 g058(.A(new_n254), .B(new_n259), .C1(KEYINPUT26), .C2(new_n258), .ZN(new_n260));
  XNOR2_X1  g059(.A(KEYINPUT27), .B(G183gat), .ZN(new_n261));
  INV_X1    g060(.A(G190gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(KEYINPUT66), .B(KEYINPUT28), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AND2_X1   g064(.A1(new_n265), .A2(KEYINPUT67), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT28), .ZN(new_n267));
  OAI22_X1  g066(.A1(new_n265), .A2(KEYINPUT67), .B1(new_n267), .B2(new_n263), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n260), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  OR2_X1    g068(.A1(G183gat), .A2(G190gat), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n270), .A2(KEYINPUT24), .A3(new_n253), .ZN(new_n271));
  OR2_X1    g070(.A1(new_n258), .A2(KEYINPUT23), .ZN(new_n272));
  OR2_X1    g071(.A1(new_n253), .A2(KEYINPUT24), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT65), .ZN(new_n275));
  OAI21_X1  g074(.A(KEYINPUT25), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n257), .B1(KEYINPUT23), .B2(new_n258), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n277), .A2(new_n271), .A3(new_n272), .A4(new_n273), .ZN(new_n278));
  AND2_X1   g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n276), .A2(new_n278), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n269), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT73), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n276), .B(new_n278), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n284), .A2(KEYINPUT73), .A3(new_n269), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n252), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n251), .A2(KEYINPUT29), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n281), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n233), .B1(new_n286), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n283), .A2(new_n287), .A3(new_n285), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n284), .A2(new_n251), .A3(new_n269), .ZN(new_n292));
  INV_X1    g091(.A(new_n225), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(G8gat), .B(G36gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(G64gat), .B(G92gat), .ZN(new_n296));
  XOR2_X1   g095(.A(new_n295), .B(new_n296), .Z(new_n297));
  NAND3_X1  g096(.A1(new_n290), .A2(new_n294), .A3(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT74), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT30), .ZN(new_n301));
  NAND4_X1  g100(.A1(new_n290), .A2(new_n294), .A3(KEYINPUT74), .A4(new_n297), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n297), .ZN(new_n304));
  INV_X1    g103(.A(new_n285), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT73), .B1(new_n284), .B2(new_n269), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n251), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n209), .B1(new_n307), .B2(new_n288), .ZN(new_n308));
  AND3_X1   g107(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n304), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n290), .A2(new_n294), .A3(KEYINPUT30), .A4(new_n297), .ZN(new_n311));
  AND2_X1   g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g111(.A(KEYINPUT82), .B1(new_n303), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n223), .A2(KEYINPUT3), .ZN(new_n315));
  XNOR2_X1  g114(.A(G113gat), .B(G120gat), .ZN(new_n316));
  INV_X1    g115(.A(G134gat), .ZN(new_n317));
  AND2_X1   g116(.A1(new_n317), .A2(G127gat), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT68), .ZN(new_n319));
  OAI22_X1  g118(.A1(new_n316), .A2(KEYINPUT1), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(G127gat), .B(G134gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n320), .B(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n315), .A2(new_n226), .A3(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT4), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n324), .B1(new_n223), .B2(new_n322), .ZN(new_n325));
  AND2_X1   g124(.A1(new_n320), .A2(new_n321), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n320), .A2(new_n321), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n328), .A2(KEYINPUT4), .A3(new_n220), .A4(new_n222), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n323), .A2(new_n325), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(G225gat), .A2(G233gat), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n328), .A2(new_n220), .A3(new_n222), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n223), .A2(new_n322), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT77), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n223), .A2(new_n322), .A3(KEYINPUT77), .ZN(new_n338));
  AND2_X1   g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n333), .B(KEYINPUT39), .C1(new_n339), .C2(new_n332), .ZN(new_n340));
  XOR2_X1   g139(.A(G1gat), .B(G29gat), .Z(new_n341));
  XNOR2_X1  g140(.A(G57gat), .B(G85gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n341), .B(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n343), .B(new_n344), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n340), .B(new_n345), .C1(KEYINPUT39), .C2(new_n333), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT40), .ZN(new_n347));
  OR2_X1    g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n337), .A2(new_n332), .A3(new_n338), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT5), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n323), .A2(new_n331), .A3(new_n325), .A4(new_n329), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT5), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n345), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n352), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n346), .A2(new_n347), .ZN(new_n358));
  AND3_X1   g157(.A1(new_n348), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n303), .A2(new_n312), .A3(KEYINPUT82), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n314), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(KEYINPUT84), .B(KEYINPUT38), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT37), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n290), .A2(new_n363), .A3(new_n294), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT85), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n290), .A2(new_n294), .A3(KEYINPUT85), .A4(new_n363), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n290), .A2(new_n294), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n297), .B1(new_n369), .B2(KEYINPUT37), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n362), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(KEYINPUT87), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT86), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n304), .A2(new_n362), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n307), .A2(new_n209), .A3(new_n288), .ZN(new_n375));
  AND2_X1   g174(.A1(new_n291), .A2(new_n292), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n375), .B1(new_n376), .B2(new_n293), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n374), .B1(new_n377), .B2(KEYINPUT37), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n373), .B1(new_n368), .B2(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n368), .A2(new_n373), .A3(new_n378), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n372), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(KEYINPUT79), .B(KEYINPUT6), .ZN(new_n383));
  OAI21_X1  g182(.A(KEYINPUT80), .B1(new_n357), .B2(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n354), .B1(new_n351), .B2(new_n350), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT80), .ZN(new_n386));
  INV_X1    g185(.A(new_n383), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n385), .A2(new_n386), .A3(new_n356), .A4(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n384), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT83), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n357), .A2(new_n383), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n385), .A2(new_n356), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n390), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n352), .A2(new_n355), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n345), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n395), .A2(KEYINPUT83), .A3(new_n357), .A4(new_n383), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n389), .B1(new_n393), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n300), .A2(new_n302), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n397), .B(new_n399), .C1(new_n371), .C2(KEYINPUT87), .ZN(new_n400));
  OAI211_X1 g199(.A(new_n248), .B(new_n361), .C1(new_n382), .C2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(G227gat), .A2(G233gat), .ZN(new_n402));
  XOR2_X1   g201(.A(new_n402), .B(KEYINPUT64), .Z(new_n403));
  NAND3_X1  g202(.A1(new_n284), .A2(new_n328), .A3(new_n269), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n328), .B1(new_n284), .B2(new_n269), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n403), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(KEYINPUT32), .ZN(new_n408));
  XNOR2_X1  g207(.A(G15gat), .B(G43gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(G71gat), .B(G99gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n409), .B(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  OAI21_X1  g211(.A(KEYINPUT33), .B1(new_n412), .B2(KEYINPUT70), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT70), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n411), .A2(new_n414), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n408), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n411), .B1(new_n407), .B2(KEYINPUT32), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT69), .ZN(new_n419));
  INV_X1    g218(.A(new_n403), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n281), .A2(new_n322), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n420), .B1(new_n421), .B2(new_n404), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n418), .B(new_n419), .C1(KEYINPUT33), .C2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT32), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n412), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n422), .A2(KEYINPUT33), .ZN(new_n426));
  OAI21_X1  g225(.A(KEYINPUT69), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n417), .B1(new_n423), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n421), .A2(new_n404), .ZN(new_n429));
  INV_X1    g228(.A(new_n402), .ZN(new_n430));
  OAI21_X1  g229(.A(KEYINPUT34), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT71), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n403), .A2(KEYINPUT34), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n432), .B1(new_n429), .B2(new_n434), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n421), .A2(KEYINPUT71), .A3(new_n404), .A4(new_n433), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n431), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  AND2_X1   g237(.A1(new_n428), .A2(new_n438), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n428), .A2(new_n438), .ZN(new_n440));
  OAI21_X1  g239(.A(KEYINPUT36), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n395), .A2(new_n357), .A3(new_n383), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n442), .A2(new_n388), .A3(new_n384), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n303), .A2(new_n312), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n247), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n423), .A2(new_n427), .ZN(new_n447));
  INV_X1    g246(.A(new_n417), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(new_n437), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT36), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n428), .A2(new_n438), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n441), .A2(new_n446), .A3(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n439), .A2(new_n440), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n444), .A2(new_n445), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n456), .A2(new_n457), .A3(new_n248), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT35), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n314), .A2(new_n360), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n397), .A2(KEYINPUT35), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n460), .A2(new_n461), .A3(new_n456), .A4(new_n248), .ZN(new_n462));
  AOI22_X1  g261(.A1(new_n401), .A2(new_n455), .B1(new_n459), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT96), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT18), .ZN(new_n465));
  INV_X1    g264(.A(G8gat), .ZN(new_n466));
  XNOR2_X1  g265(.A(G15gat), .B(G22gat), .ZN(new_n467));
  INV_X1    g266(.A(G1gat), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT16), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n467), .A2(G1gat), .ZN(new_n472));
  OAI211_X1 g271(.A(KEYINPUT93), .B(new_n466), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n472), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n466), .A2(KEYINPUT93), .ZN(new_n475));
  OR2_X1    g274(.A1(new_n466), .A2(KEYINPUT93), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n474), .A2(new_n470), .A3(new_n475), .A4(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT15), .ZN(new_n480));
  INV_X1    g279(.A(G43gat), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n481), .A2(G50gat), .ZN(new_n482));
  INV_X1    g281(.A(G50gat), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n483), .A2(G43gat), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n480), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n483), .A2(G43gat), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n481), .A2(G50gat), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n486), .A2(new_n487), .A3(KEYINPUT15), .ZN(new_n488));
  NAND2_X1  g287(.A1(KEYINPUT90), .A2(G29gat), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  NOR2_X1   g289(.A1(KEYINPUT90), .A2(G29gat), .ZN(new_n491));
  OAI21_X1  g290(.A(G36gat), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n485), .A2(new_n488), .A3(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT14), .ZN(new_n496));
  INV_X1    g295(.A(G29gat), .ZN(new_n497));
  INV_X1    g296(.A(G36gat), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT91), .ZN(new_n500));
  NOR2_X1   g299(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT91), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n501), .A2(new_n502), .A3(new_n498), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n495), .B1(new_n500), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g303(.A(KEYINPUT92), .B1(new_n493), .B2(new_n504), .ZN(new_n505));
  OR2_X1    g304(.A1(KEYINPUT90), .A2(G29gat), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n498), .B1(new_n506), .B2(new_n489), .ZN(new_n507));
  AOI21_X1  g306(.A(KEYINPUT15), .B1(new_n486), .B2(new_n487), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NOR4_X1   g308(.A1(KEYINPUT91), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n502), .B1(new_n501), .B2(new_n498), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n494), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT92), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n509), .A2(new_n512), .A3(new_n513), .A4(new_n488), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n505), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n507), .A2(new_n494), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n499), .A2(KEYINPUT15), .A3(new_n486), .A4(new_n487), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT17), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n518), .B1(new_n505), .B2(new_n514), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT17), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n479), .B1(new_n521), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n520), .A2(new_n479), .ZN(new_n526));
  NAND2_X1  g325(.A1(G229gat), .A2(G233gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n465), .B1(new_n525), .B2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT94), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n530), .B1(new_n522), .B2(new_n478), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(new_n526), .ZN(new_n532));
  XOR2_X1   g331(.A(new_n527), .B(KEYINPUT13), .Z(new_n533));
  NAND3_X1  g332(.A1(new_n520), .A2(new_n530), .A3(new_n479), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n523), .B1(new_n515), .B2(new_n519), .ZN(new_n536));
  AOI211_X1 g335(.A(KEYINPUT17), .B(new_n518), .C1(new_n505), .C2(new_n514), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n478), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  AOI22_X1  g337(.A1(new_n520), .A2(new_n479), .B1(G229gat), .B2(G233gat), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n538), .A2(KEYINPUT18), .A3(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n529), .A2(new_n535), .A3(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(G113gat), .B(G141gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(KEYINPUT88), .B(G197gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(KEYINPUT11), .B(G169gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  XOR2_X1   g345(.A(KEYINPUT89), .B(KEYINPUT12), .Z(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT95), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n529), .A2(new_n540), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n548), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AND2_X1   g352(.A1(new_n535), .A2(new_n548), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n554), .A2(KEYINPUT95), .A3(new_n529), .A4(new_n540), .ZN(new_n555));
  AOI221_X4 g354(.A(new_n464), .B1(new_n541), .B2(new_n549), .C1(new_n553), .C2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n553), .A2(new_n555), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n549), .ZN(new_n558));
  AOI21_X1  g357(.A(KEYINPUT96), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n463), .A2(new_n560), .ZN(new_n561));
  XOR2_X1   g360(.A(G183gat), .B(G211gat), .Z(new_n562));
  OR2_X1    g361(.A1(G57gat), .A2(G64gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(G57gat), .A2(G64gat), .ZN(new_n564));
  AND2_X1   g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT9), .ZN(new_n566));
  INV_X1    g365(.A(G71gat), .ZN(new_n567));
  INV_X1    g366(.A(G78gat), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  XOR2_X1   g368(.A(G71gat), .B(G78gat), .Z(new_n570));
  OAI211_X1 g369(.A(new_n565), .B(new_n569), .C1(new_n570), .C2(KEYINPUT97), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n569), .A2(new_n563), .A3(new_n564), .ZN(new_n572));
  XNOR2_X1  g371(.A(G71gat), .B(G78gat), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n563), .A2(KEYINPUT97), .A3(new_n564), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  AND2_X1   g375(.A1(G231gat), .A2(G233gat), .ZN(new_n577));
  OR3_X1    g376(.A1(new_n576), .A2(KEYINPUT21), .A3(new_n577), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n577), .B1(new_n576), .B2(KEYINPUT21), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(G127gat), .B(G155gat), .ZN(new_n581));
  XOR2_X1   g380(.A(new_n581), .B(KEYINPUT20), .Z(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n580), .A2(new_n582), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n562), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n585), .ZN(new_n587));
  INV_X1    g386(.A(new_n562), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n587), .A2(new_n588), .A3(new_n583), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n576), .A2(KEYINPUT21), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n478), .A2(new_n590), .ZN(new_n591));
  XOR2_X1   g390(.A(KEYINPUT98), .B(KEYINPUT19), .Z(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  AND3_X1   g392(.A1(new_n586), .A2(new_n589), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n593), .B1(new_n586), .B2(new_n589), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(G232gat), .A2(G233gat), .ZN(new_n597));
  XOR2_X1   g396(.A(new_n597), .B(KEYINPUT99), .Z(new_n598));
  INV_X1    g397(.A(KEYINPUT41), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT101), .ZN(new_n601));
  INV_X1    g400(.A(G85gat), .ZN(new_n602));
  INV_X1    g401(.A(G92gat), .ZN(new_n603));
  OAI21_X1  g402(.A(KEYINPUT7), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT7), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n605), .A2(G85gat), .A3(G92gat), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT100), .ZN(new_n608));
  NAND2_X1  g407(.A1(G99gat), .A2(G106gat), .ZN(new_n609));
  AOI22_X1  g408(.A1(KEYINPUT8), .A2(new_n609), .B1(new_n602), .B2(new_n603), .ZN(new_n610));
  AND3_X1   g409(.A1(new_n607), .A2(new_n608), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n608), .B1(new_n607), .B2(new_n610), .ZN(new_n612));
  XOR2_X1   g411(.A(G99gat), .B(G106gat), .Z(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NOR3_X1   g413(.A1(new_n611), .A2(new_n612), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n607), .A2(new_n610), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(KEYINPUT100), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n607), .A2(new_n608), .A3(new_n610), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n613), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n601), .B1(new_n615), .B2(new_n619), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n614), .B1(new_n611), .B2(new_n612), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n617), .A2(new_n613), .A3(new_n618), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n621), .A2(new_n622), .A3(KEYINPUT101), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n600), .B1(new_n625), .B2(new_n520), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n624), .B1(new_n536), .B2(new_n537), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(G190gat), .B(G218gat), .ZN(new_n629));
  XOR2_X1   g428(.A(new_n629), .B(KEYINPUT102), .Z(new_n630));
  NAND2_X1  g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n630), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n626), .A2(new_n632), .A3(new_n627), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n598), .A2(new_n599), .ZN(new_n635));
  XNOR2_X1  g434(.A(G134gat), .B(G162gat), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n635), .B(new_n636), .Z(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n631), .A2(new_n637), .A3(new_n633), .ZN(new_n640));
  NAND2_X1  g439(.A1(G230gat), .A2(G233gat), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT10), .ZN(new_n643));
  AOI22_X1  g442(.A1(new_n571), .A2(new_n575), .B1(KEYINPUT103), .B2(new_n616), .ZN(new_n644));
  AND3_X1   g443(.A1(new_n621), .A2(new_n644), .A3(new_n622), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n644), .B1(new_n622), .B2(new_n621), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n643), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n643), .B1(new_n571), .B2(new_n575), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n620), .A2(new_n623), .A3(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n642), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  NOR3_X1   g449(.A1(new_n645), .A2(new_n646), .A3(new_n641), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(G120gat), .B(G148gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(G176gat), .B(G204gat), .ZN(new_n654));
  XOR2_X1   g453(.A(new_n653), .B(new_n654), .Z(new_n655));
  NOR2_X1   g454(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n655), .ZN(new_n657));
  NOR3_X1   g456(.A1(new_n650), .A2(new_n651), .A3(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  AND4_X1   g458(.A1(new_n596), .A2(new_n639), .A3(new_n640), .A4(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n561), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n661), .A2(new_n443), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(new_n468), .ZN(G1324gat));
  NOR2_X1   g462(.A1(new_n661), .A2(new_n460), .ZN(new_n664));
  XOR2_X1   g463(.A(KEYINPUT16), .B(G8gat), .Z(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n666), .B1(new_n466), .B2(new_n664), .ZN(new_n667));
  MUX2_X1   g466(.A(new_n666), .B(new_n667), .S(KEYINPUT42), .Z(G1325gat));
  NAND2_X1  g467(.A1(new_n441), .A2(new_n453), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(G15gat), .B1(new_n661), .B2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n456), .ZN(new_n672));
  OR2_X1    g471(.A1(new_n672), .A2(G15gat), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n671), .B1(new_n661), .B2(new_n673), .ZN(G1326gat));
  NOR2_X1   g473(.A1(new_n661), .A2(new_n248), .ZN(new_n675));
  XOR2_X1   g474(.A(KEYINPUT43), .B(G22gat), .Z(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(G1327gat));
  NAND2_X1  g476(.A1(new_n401), .A2(new_n455), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n459), .A2(new_n462), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n560), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n639), .A2(new_n640), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n596), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(new_n659), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n680), .A2(new_n681), .A3(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NAND4_X1  g487(.A1(new_n688), .A2(new_n444), .A3(new_n506), .A4(new_n489), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT45), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT44), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n691), .B1(new_n463), .B2(new_n683), .ZN(new_n692));
  AND3_X1   g491(.A1(new_n303), .A2(new_n312), .A3(KEYINPUT82), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n693), .A2(new_n313), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n247), .B1(new_n694), .B2(new_n359), .ZN(new_n695));
  INV_X1    g494(.A(new_n379), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(new_n380), .ZN(new_n697));
  AOI211_X1 g496(.A(new_n389), .B(new_n398), .C1(new_n393), .C2(new_n396), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n368), .A2(new_n370), .ZN(new_n699));
  INV_X1    g498(.A(new_n362), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT87), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n697), .A2(new_n698), .A3(new_n703), .A4(new_n372), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n454), .B1(new_n695), .B2(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n450), .A2(new_n248), .A3(new_n452), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n706), .A2(KEYINPUT35), .A3(new_n397), .ZN(new_n707));
  AOI22_X1  g506(.A1(new_n707), .A2(new_n460), .B1(new_n458), .B2(KEYINPUT35), .ZN(new_n708));
  OAI211_X1 g507(.A(KEYINPUT44), .B(new_n682), .C1(new_n705), .C2(new_n708), .ZN(new_n709));
  AND2_X1   g508(.A1(new_n692), .A2(new_n709), .ZN(new_n710));
  AND3_X1   g509(.A1(new_n538), .A2(KEYINPUT18), .A3(new_n539), .ZN(new_n711));
  AOI21_X1  g510(.A(KEYINPUT18), .B1(new_n538), .B2(new_n539), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g512(.A(KEYINPUT95), .B1(new_n713), .B2(new_n554), .ZN(new_n714));
  NOR4_X1   g513(.A1(new_n552), .A2(new_n711), .A3(new_n712), .A4(new_n550), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n558), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n717), .A2(new_n685), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n710), .A2(new_n444), .A3(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(new_n491), .B2(new_n490), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n690), .A2(new_n720), .ZN(G1328gat));
  INV_X1    g520(.A(KEYINPUT46), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n460), .A2(G36gat), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n722), .B1(new_n688), .B2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n723), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n687), .A2(KEYINPUT46), .A3(new_n725), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n692), .A2(new_n694), .A3(new_n709), .A4(new_n718), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT104), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(G36gat), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n728), .A2(new_n729), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n727), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT105), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  OAI211_X1 g534(.A(new_n727), .B(KEYINPUT105), .C1(new_n731), .C2(new_n732), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(G1329gat));
  NAND4_X1  g536(.A1(new_n692), .A2(new_n669), .A3(new_n709), .A4(new_n718), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(G43gat), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n688), .A2(new_n481), .A3(new_n456), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  XOR2_X1   g540(.A(new_n741), .B(KEYINPUT47), .Z(G1330gat));
  OR2_X1    g541(.A1(new_n687), .A2(KEYINPUT106), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n687), .A2(KEYINPUT106), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n743), .A2(new_n483), .A3(new_n247), .A4(new_n744), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n692), .A2(new_n247), .A3(new_n709), .A4(new_n718), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(G50gat), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT48), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n748), .B(new_n749), .ZN(G1331gat));
  NOR4_X1   g549(.A1(new_n682), .A2(new_n716), .A3(new_n684), .A4(new_n659), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n680), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n752), .A2(new_n443), .ZN(new_n753));
  XOR2_X1   g552(.A(KEYINPUT107), .B(G57gat), .Z(new_n754));
  XNOR2_X1  g553(.A(new_n753), .B(new_n754), .ZN(G1332gat));
  NOR2_X1   g554(.A1(new_n752), .A2(new_n460), .ZN(new_n756));
  NOR2_X1   g555(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n757));
  AND2_X1   g556(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n756), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n759), .B1(new_n756), .B2(new_n757), .ZN(G1333gat));
  OAI21_X1  g559(.A(new_n567), .B1(new_n752), .B2(new_n672), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n680), .A2(G71gat), .A3(new_n669), .A4(new_n751), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT108), .ZN(new_n763));
  AND2_X1   g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n762), .A2(new_n763), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n761), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g566(.A1(new_n752), .A2(new_n248), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(new_n568), .ZN(G1335gat));
  NAND2_X1  g568(.A1(new_n717), .A2(new_n684), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(KEYINPUT109), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n682), .B(new_n771), .C1(new_n705), .C2(new_n708), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT51), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n772), .A2(new_n773), .ZN(new_n775));
  OR2_X1    g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(new_n659), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n776), .A2(new_n602), .A3(new_n444), .A4(new_n777), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n771), .A2(new_n777), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n710), .A2(new_n444), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(G85gat), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n778), .A2(new_n781), .ZN(G1336gat));
  INV_X1    g581(.A(KEYINPUT111), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n460), .A2(G92gat), .A3(new_n659), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n784), .B1(new_n774), .B2(new_n775), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n692), .A2(new_n694), .A3(new_n709), .A4(new_n779), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(G92gat), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT52), .ZN(new_n788));
  AND3_X1   g587(.A1(new_n785), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT110), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n772), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(new_n773), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n772), .A2(new_n790), .A3(KEYINPUT51), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n792), .A2(new_n793), .A3(new_n784), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n788), .B1(new_n794), .B2(new_n787), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n783), .B1(new_n789), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n785), .A2(new_n787), .A3(new_n788), .ZN(new_n797));
  AND3_X1   g596(.A1(new_n772), .A2(new_n790), .A3(KEYINPUT51), .ZN(new_n798));
  AOI21_X1  g597(.A(KEYINPUT51), .B1(new_n772), .B2(new_n790), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AOI22_X1  g599(.A1(new_n800), .A2(new_n784), .B1(G92gat), .B2(new_n786), .ZN(new_n801));
  OAI211_X1 g600(.A(KEYINPUT111), .B(new_n797), .C1(new_n801), .C2(new_n788), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n796), .A2(new_n802), .ZN(G1337gat));
  NOR3_X1   g602(.A1(new_n672), .A2(G99gat), .A3(new_n659), .ZN(new_n804));
  XOR2_X1   g603(.A(new_n804), .B(KEYINPUT113), .Z(new_n805));
  NAND2_X1  g604(.A1(new_n776), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n710), .A2(new_n669), .A3(new_n779), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT112), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(G99gat), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n807), .A2(new_n808), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n806), .B1(new_n810), .B2(new_n811), .ZN(G1338gat));
  NOR3_X1   g611(.A1(new_n248), .A2(G106gat), .A3(new_n659), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n813), .B1(new_n774), .B2(new_n775), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n692), .A2(new_n247), .A3(new_n709), .A4(new_n779), .ZN(new_n815));
  XOR2_X1   g614(.A(KEYINPUT114), .B(G106gat), .Z(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n818));
  AND3_X1   g617(.A1(new_n814), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n792), .A2(new_n793), .A3(new_n813), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n818), .B1(new_n820), .B2(new_n817), .ZN(new_n821));
  OAI21_X1  g620(.A(KEYINPUT115), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT115), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n814), .A2(new_n817), .A3(new_n818), .ZN(new_n824));
  AOI22_X1  g623(.A1(new_n800), .A2(new_n813), .B1(new_n815), .B2(new_n816), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n823), .B(new_n824), .C1(new_n825), .C2(new_n818), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n822), .A2(new_n826), .ZN(G1339gat));
  AND2_X1   g626(.A1(new_n660), .A2(new_n717), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n620), .A2(new_n623), .A3(new_n648), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n616), .A2(KEYINPUT103), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n576), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n831), .B1(new_n615), .B2(new_n619), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n621), .A2(new_n644), .A3(new_n622), .ZN(new_n833));
  AOI21_X1  g632(.A(KEYINPUT10), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n641), .B1(new_n829), .B2(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n647), .A2(new_n642), .A3(new_n649), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n835), .A2(new_n836), .A3(KEYINPUT54), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT54), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n655), .B1(new_n650), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n837), .A2(new_n839), .A3(KEYINPUT55), .ZN(new_n840));
  INV_X1    g639(.A(new_n658), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT55), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n837), .A2(new_n839), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n842), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n845), .A2(new_n716), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n527), .B1(new_n538), .B2(new_n526), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n533), .B1(new_n532), .B2(new_n534), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n546), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n777), .A2(new_n557), .A3(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n683), .B1(new_n846), .B2(new_n850), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n557), .A2(new_n849), .ZN(new_n852));
  AND3_X1   g651(.A1(new_n852), .A2(new_n845), .A3(new_n682), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(KEYINPUT116), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n852), .A2(new_n845), .A3(new_n682), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT116), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n851), .A2(new_n854), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n828), .B1(new_n858), .B2(new_n684), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n460), .A2(new_n444), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n859), .A2(new_n706), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(G113gat), .B1(new_n861), .B2(new_n716), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n681), .A2(G113gat), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n862), .B1(new_n861), .B2(new_n863), .ZN(G1340gat));
  NAND2_X1  g663(.A1(new_n861), .A2(new_n777), .ZN(new_n865));
  XNOR2_X1  g664(.A(new_n865), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g665(.A1(new_n861), .A2(new_n596), .ZN(new_n867));
  XNOR2_X1  g666(.A(new_n867), .B(G127gat), .ZN(G1342gat));
  AOI21_X1  g667(.A(new_n317), .B1(new_n861), .B2(new_n682), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n861), .A2(new_n317), .A3(new_n682), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n870), .A2(KEYINPUT117), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(KEYINPUT117), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n869), .B1(new_n873), .B2(KEYINPUT56), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT56), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n871), .A2(new_n875), .A3(new_n872), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n876), .A2(new_n877), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n874), .B1(new_n878), .B2(new_n879), .ZN(G1343gat));
  INV_X1    g679(.A(new_n214), .ZN(new_n881));
  INV_X1    g680(.A(new_n860), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(new_n670), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT57), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n248), .A2(new_n884), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n854), .A2(new_n857), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT119), .ZN(new_n887));
  AND3_X1   g686(.A1(new_n647), .A2(new_n642), .A3(new_n649), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n888), .A2(new_n650), .A3(new_n838), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n657), .B1(new_n835), .B2(KEYINPUT54), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n887), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n837), .A2(new_n839), .A3(KEYINPUT119), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n891), .A2(new_n843), .A3(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(new_n842), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n716), .A2(new_n464), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n557), .A2(KEYINPUT96), .A3(new_n558), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n683), .B1(new_n898), .B2(new_n850), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n596), .B1(new_n886), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n885), .B1(new_n900), .B2(new_n828), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n884), .B1(new_n859), .B2(new_n248), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n883), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n881), .B1(new_n903), .B2(new_n716), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n859), .A2(new_n248), .A3(new_n669), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(new_n882), .ZN(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n560), .A2(G141gat), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n904), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT58), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n881), .B1(new_n903), .B2(new_n681), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n907), .A2(new_n908), .ZN(new_n912));
  XOR2_X1   g711(.A(KEYINPUT120), .B(KEYINPUT58), .Z(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI22_X1  g713(.A1(new_n909), .A2(new_n910), .B1(new_n911), .B2(new_n914), .ZN(G1344gat));
  NAND3_X1  g714(.A1(new_n907), .A2(new_n215), .A3(new_n777), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT59), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT122), .ZN(new_n918));
  AOI21_X1  g717(.A(KEYINPUT55), .B1(new_n844), .B2(new_n887), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n842), .B1(new_n919), .B2(new_n892), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n920), .B1(new_n556), .B2(new_n559), .ZN(new_n921));
  INV_X1    g720(.A(new_n850), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n682), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n684), .B1(new_n923), .B2(new_n853), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n660), .A2(new_n896), .A3(new_n897), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT121), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n560), .A2(KEYINPUT121), .A3(new_n660), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n248), .B1(new_n924), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n918), .B1(new_n930), .B2(KEYINPUT57), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n927), .A2(new_n928), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n899), .A2(new_n855), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n932), .B1(new_n933), .B2(new_n684), .ZN(new_n934));
  OAI211_X1 g733(.A(KEYINPUT122), .B(new_n884), .C1(new_n934), .C2(new_n248), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n858), .A2(new_n684), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n885), .B1(new_n936), .B2(new_n828), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n931), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n883), .A2(new_n659), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n917), .B1(new_n940), .B2(G148gat), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n917), .A2(G148gat), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n942), .B1(new_n903), .B2(new_n777), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n916), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(KEYINPUT123), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT123), .ZN(new_n946));
  OAI211_X1 g745(.A(new_n946), .B(new_n916), .C1(new_n941), .C2(new_n943), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n945), .A2(new_n947), .ZN(G1345gat));
  INV_X1    g747(.A(new_n903), .ZN(new_n949));
  OAI21_X1  g748(.A(G155gat), .B1(new_n949), .B2(new_n684), .ZN(new_n950));
  OR2_X1    g749(.A1(new_n684), .A2(G155gat), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n950), .B1(new_n906), .B2(new_n951), .ZN(G1346gat));
  AOI21_X1  g751(.A(G162gat), .B1(new_n907), .B2(new_n682), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n682), .A2(G162gat), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n953), .B1(new_n903), .B2(new_n954), .ZN(G1347gat));
  NOR2_X1   g754(.A1(new_n859), .A2(new_n706), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n460), .A2(new_n444), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n957), .B(KEYINPUT125), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NOR3_X1   g758(.A1(new_n959), .A2(new_n255), .A3(new_n560), .ZN(new_n960));
  AND2_X1   g759(.A1(new_n956), .A2(new_n957), .ZN(new_n961));
  XOR2_X1   g760(.A(new_n961), .B(KEYINPUT124), .Z(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(new_n716), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n960), .B1(new_n963), .B2(new_n255), .ZN(G1348gat));
  NAND3_X1  g763(.A1(new_n962), .A2(new_n256), .A3(new_n777), .ZN(new_n965));
  OAI21_X1  g764(.A(G176gat), .B1(new_n959), .B2(new_n659), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(new_n966), .ZN(G1349gat));
  NAND3_X1  g766(.A1(new_n961), .A2(new_n261), .A3(new_n596), .ZN(new_n968));
  OAI21_X1  g767(.A(G183gat), .B1(new_n959), .B2(new_n684), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT126), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  XNOR2_X1  g770(.A(new_n971), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g771(.A1(new_n962), .A2(new_n262), .A3(new_n682), .ZN(new_n973));
  OAI21_X1  g772(.A(G190gat), .B1(new_n959), .B2(new_n683), .ZN(new_n974));
  XNOR2_X1  g773(.A(new_n974), .B(KEYINPUT61), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n973), .A2(new_n975), .ZN(G1351gat));
  NAND2_X1  g775(.A1(new_n958), .A2(new_n670), .ZN(new_n977));
  OR2_X1    g776(.A1(new_n977), .A2(KEYINPUT127), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n977), .A2(KEYINPUT127), .ZN(new_n979));
  AND3_X1   g778(.A1(new_n978), .A2(new_n938), .A3(new_n979), .ZN(new_n980));
  INV_X1    g779(.A(G197gat), .ZN(new_n981));
  NOR2_X1   g780(.A1(new_n560), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n905), .A2(new_n716), .A3(new_n957), .ZN(new_n983));
  AOI22_X1  g782(.A1(new_n980), .A2(new_n982), .B1(new_n981), .B2(new_n983), .ZN(G1352gat));
  NAND2_X1  g783(.A1(new_n980), .A2(new_n777), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n985), .A2(G204gat), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n905), .A2(new_n957), .ZN(new_n987));
  NOR3_X1   g786(.A1(new_n987), .A2(G204gat), .A3(new_n659), .ZN(new_n988));
  XNOR2_X1  g787(.A(new_n988), .B(KEYINPUT62), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n986), .A2(new_n989), .ZN(G1353gat));
  NAND4_X1  g789(.A1(new_n938), .A2(new_n670), .A3(new_n596), .A4(new_n958), .ZN(new_n991));
  AND3_X1   g790(.A1(new_n991), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n992));
  AOI21_X1  g791(.A(KEYINPUT63), .B1(new_n991), .B2(G211gat), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n596), .A2(new_n204), .ZN(new_n994));
  OAI22_X1  g793(.A1(new_n992), .A2(new_n993), .B1(new_n987), .B2(new_n994), .ZN(G1354gat));
  AOI21_X1  g794(.A(new_n205), .B1(new_n980), .B2(new_n682), .ZN(new_n996));
  NOR3_X1   g795(.A1(new_n987), .A2(G218gat), .A3(new_n683), .ZN(new_n997));
  OR2_X1    g796(.A1(new_n996), .A2(new_n997), .ZN(G1355gat));
endmodule


