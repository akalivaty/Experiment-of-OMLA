//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 1 1 1 0 0 0 0 1 1 1 0 1 1 1 0 1 1 0 1 1 1 0 0 0 0 0 0 1 0 0 1 0 1 1 1 0 1 1 0 0 1 0 0 0 0 0 0 1 1 1 0 0 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:01 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n551,
    new_n553, new_n554, new_n556, new_n557, new_n558, new_n559, new_n562,
    new_n563, new_n565, new_n566, new_n567, new_n568, new_n569, new_n571,
    new_n572, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n585, new_n586, new_n589, new_n591,
    new_n592, new_n593, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1128, new_n1129, new_n1130,
    new_n1131;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT65), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n462), .A2(new_n463), .A3(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(KEYINPUT67), .B1(new_n465), .B2(KEYINPUT3), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n467));
  OAI211_X1 g042(.A(new_n461), .B(new_n464), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G137), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n463), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G125), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n471), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(G101), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n465), .A2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n470), .B(new_n477), .C1(new_n478), .C2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G160));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n484));
  INV_X1    g059(.A(G136), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n484), .B1(new_n468), .B2(new_n485), .ZN(new_n486));
  OAI211_X1 g061(.A(G2105), .B(new_n464), .C1(new_n466), .C2(new_n467), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n486), .B1(G124), .B2(new_n488), .ZN(G162));
  INV_X1    g064(.A(G126), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n461), .A2(G114), .ZN(new_n491));
  OAI21_X1  g066(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n492));
  OAI22_X1  g067(.A1(new_n487), .A2(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n494), .A2(new_n461), .A3(G138), .ZN(new_n495));
  NOR3_X1   g070(.A1(new_n474), .A2(KEYINPUT68), .A3(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT68), .ZN(new_n497));
  XNOR2_X1  g072(.A(KEYINPUT3), .B(G2104), .ZN(new_n498));
  INV_X1    g073(.A(G138), .ZN(new_n499));
  NOR3_X1   g074(.A1(new_n499), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n497), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n496), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g077(.A(KEYINPUT4), .B1(new_n468), .B2(new_n499), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n493), .B1(new_n502), .B2(new_n503), .ZN(G164));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n510), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  OR2_X1    g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT6), .B(G651), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n514), .A2(G50), .A3(G543), .ZN(new_n515));
  XNOR2_X1  g090(.A(new_n515), .B(KEYINPUT69), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n510), .A2(new_n514), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G88), .ZN(new_n519));
  AND3_X1   g094(.A1(new_n516), .A2(KEYINPUT70), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g095(.A(KEYINPUT70), .B1(new_n516), .B2(new_n519), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n513), .B1(new_n520), .B2(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  NAND2_X1  g098(.A1(G76), .A2(G543), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT7), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT71), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n509), .B(new_n527), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n526), .B1(new_n528), .B2(G63), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n529), .A2(new_n512), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n525), .B1(new_n524), .B2(new_n512), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n514), .A2(G543), .ZN(new_n532));
  INV_X1    g107(.A(G51), .ZN(new_n533));
  XNOR2_X1  g108(.A(KEYINPUT72), .B(G89), .ZN(new_n534));
  OAI221_X1 g109(.A(new_n531), .B1(new_n532), .B2(new_n533), .C1(new_n517), .C2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n530), .A2(new_n535), .ZN(G168));
  AOI22_X1  g111(.A1(new_n528), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n512), .ZN(new_n538));
  INV_X1    g113(.A(G90), .ZN(new_n539));
  XNOR2_X1  g114(.A(KEYINPUT73), .B(G52), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n517), .A2(new_n539), .B1(new_n532), .B2(new_n540), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n538), .A2(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  AOI22_X1  g118(.A1(new_n528), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n544), .A2(new_n512), .ZN(new_n545));
  XOR2_X1   g120(.A(KEYINPUT74), .B(G81), .Z(new_n546));
  INV_X1    g121(.A(new_n532), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n518), .A2(new_n546), .B1(new_n547), .B2(G43), .ZN(new_n548));
  AND2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  AND3_X1   g125(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G36), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n551), .A2(new_n554), .ZN(G188));
  NAND2_X1  g130(.A1(new_n547), .A2(G53), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT9), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n518), .A2(G91), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n510), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n559));
  OAI211_X1 g134(.A(new_n557), .B(new_n558), .C1(new_n512), .C2(new_n559), .ZN(G299));
  INV_X1    g135(.A(G168), .ZN(G286));
  AOI22_X1  g136(.A1(new_n518), .A2(G87), .B1(G49), .B2(new_n547), .ZN(new_n562));
  OAI21_X1  g137(.A(G651), .B1(new_n528), .B2(G74), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(G288));
  AOI22_X1  g139(.A1(new_n510), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n565), .A2(new_n512), .ZN(new_n566));
  INV_X1    g141(.A(G86), .ZN(new_n567));
  INV_X1    g142(.A(G48), .ZN(new_n568));
  OAI22_X1  g143(.A1(new_n517), .A2(new_n567), .B1(new_n532), .B2(new_n568), .ZN(new_n569));
  OR2_X1    g144(.A1(new_n566), .A2(new_n569), .ZN(G305));
  AOI22_X1  g145(.A1(new_n518), .A2(G85), .B1(G47), .B2(new_n547), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n528), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n572), .B2(new_n512), .ZN(G290));
  NAND2_X1  g148(.A1(G301), .A2(G868), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n518), .A2(G92), .ZN(new_n575));
  XOR2_X1   g150(.A(new_n575), .B(KEYINPUT10), .Z(new_n576));
  NAND2_X1  g151(.A1(G79), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(G66), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n509), .B2(new_n578), .ZN(new_n579));
  AOI22_X1  g154(.A1(G54), .A2(new_n547), .B1(new_n579), .B2(G651), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n574), .B1(new_n582), .B2(G868), .ZN(G284));
  OAI21_X1  g158(.A(new_n574), .B1(new_n582), .B2(G868), .ZN(G321));
  INV_X1    g159(.A(G868), .ZN(new_n585));
  NAND2_X1  g160(.A1(G299), .A2(new_n585), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n586), .B1(new_n585), .B2(G168), .ZN(G297));
  XOR2_X1   g162(.A(G297), .B(KEYINPUT75), .Z(G280));
  INV_X1    g163(.A(G559), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n582), .B1(new_n589), .B2(G860), .ZN(G148));
  NAND2_X1  g165(.A1(new_n582), .A2(new_n589), .ZN(new_n591));
  XNOR2_X1  g166(.A(new_n591), .B(KEYINPUT76), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(G868), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n593), .B1(G868), .B2(new_n549), .ZN(G323));
  XNOR2_X1  g169(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g170(.A1(new_n474), .A2(new_n480), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n596), .B(KEYINPUT12), .ZN(new_n597));
  INV_X1    g172(.A(G2100), .ZN(new_n598));
  OAI22_X1  g173(.A1(new_n597), .A2(KEYINPUT13), .B1(KEYINPUT77), .B2(new_n598), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n599), .B1(KEYINPUT13), .B2(new_n597), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n598), .A2(KEYINPUT77), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n600), .B(new_n601), .ZN(new_n602));
  OR2_X1    g177(.A1(G99), .A2(G2105), .ZN(new_n603));
  OAI211_X1 g178(.A(new_n603), .B(G2104), .C1(G111), .C2(new_n461), .ZN(new_n604));
  INV_X1    g179(.A(G135), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n468), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n606), .B1(G123), .B2(new_n488), .ZN(new_n607));
  XNOR2_X1  g182(.A(KEYINPUT78), .B(G2096), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n607), .B(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n602), .A2(new_n609), .ZN(G156));
  INV_X1    g185(.A(KEYINPUT14), .ZN(new_n611));
  XNOR2_X1  g186(.A(KEYINPUT15), .B(G2430), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(G2435), .ZN(new_n613));
  XNOR2_X1  g188(.A(G2427), .B(G2438), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n611), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(new_n614), .B2(new_n613), .ZN(new_n616));
  XNOR2_X1  g191(.A(G2451), .B(G2454), .ZN(new_n617));
  XNOR2_X1  g192(.A(KEYINPUT16), .B(G1341), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  XNOR2_X1  g194(.A(G2443), .B(G2446), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G1348), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n619), .B(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(G14), .B1(new_n616), .B2(new_n622), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n623), .B1(new_n616), .B2(new_n622), .ZN(G401));
  XOR2_X1   g199(.A(G2084), .B(G2090), .Z(new_n625));
  INV_X1    g200(.A(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(G2067), .B(G2678), .Z(new_n627));
  NOR2_X1   g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(G2072), .B(G2078), .Z(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT18), .Z(new_n632));
  NAND2_X1  g207(.A1(new_n626), .A2(new_n627), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n633), .B1(KEYINPUT79), .B2(new_n630), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(KEYINPUT79), .B2(new_n630), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n629), .B(KEYINPUT17), .Z(new_n636));
  INV_X1    g211(.A(new_n628), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(new_n633), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n632), .B(new_n635), .C1(new_n636), .C2(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G2096), .B(G2100), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(G227));
  XOR2_X1   g216(.A(G1971), .B(G1976), .Z(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT80), .B(KEYINPUT19), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G1956), .B(G2474), .Z(new_n645));
  XOR2_X1   g220(.A(G1961), .B(G1966), .Z(new_n646));
  AND2_X1   g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AND2_X1   g222(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n648), .A2(KEYINPUT20), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n648), .A2(KEYINPUT20), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n645), .A2(new_n646), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n644), .A2(new_n651), .ZN(new_n652));
  OR3_X1    g227(.A1(new_n644), .A2(new_n647), .A3(new_n651), .ZN(new_n653));
  NAND4_X1  g228(.A1(new_n649), .A2(new_n650), .A3(new_n652), .A4(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G1991), .B(G1996), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT81), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n654), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G1981), .B(G1986), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(G229));
  INV_X1    g236(.A(G16), .ZN(new_n662));
  NOR2_X1   g237(.A1(G166), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n663), .B1(new_n662), .B2(G22), .ZN(new_n664));
  INV_X1    g239(.A(G1971), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n664), .A2(new_n665), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n662), .A2(G6), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n566), .A2(new_n569), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n668), .B1(new_n669), .B2(new_n662), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT32), .B(G1981), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n670), .A2(new_n671), .ZN(new_n673));
  INV_X1    g248(.A(G288), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n674), .A2(G16), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n675), .B1(G16), .B2(G23), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT33), .B(G1976), .Z(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  OAI211_X1 g253(.A(new_n672), .B(new_n673), .C1(new_n676), .C2(new_n678), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n679), .B1(new_n676), .B2(new_n678), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n666), .A2(new_n667), .A3(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(KEYINPUT34), .Z(new_n682));
  INV_X1    g257(.A(G29), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(G25), .ZN(new_n684));
  AND2_X1   g259(.A1(new_n488), .A2(G119), .ZN(new_n685));
  OR2_X1    g260(.A1(G95), .A2(G2105), .ZN(new_n686));
  OAI211_X1 g261(.A(new_n686), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n687));
  INV_X1    g262(.A(G131), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n687), .B1(new_n468), .B2(new_n688), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n684), .B1(new_n691), .B2(new_n683), .ZN(new_n692));
  XOR2_X1   g267(.A(KEYINPUT35), .B(G1991), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  MUX2_X1   g269(.A(G24), .B(G290), .S(G16), .Z(new_n695));
  OR2_X1    g270(.A1(new_n695), .A2(G1986), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(G1986), .ZN(new_n697));
  NAND4_X1  g272(.A1(new_n682), .A2(new_n694), .A3(new_n696), .A4(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(KEYINPUT36), .Z(new_n699));
  NAND2_X1  g274(.A1(new_n662), .A2(G5), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(G171), .B2(new_n662), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT96), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G1961), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT97), .Z(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT89), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n683), .A2(G26), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(G140), .ZN(new_n709));
  OR3_X1    g284(.A1(new_n468), .A2(KEYINPUT86), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n488), .A2(G128), .ZN(new_n711));
  OAI21_X1  g286(.A(KEYINPUT86), .B1(new_n468), .B2(new_n709), .ZN(new_n712));
  OR2_X1    g287(.A1(G104), .A2(G2105), .ZN(new_n713));
  OAI211_X1 g288(.A(new_n713), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n714));
  NAND4_X1  g289(.A1(new_n710), .A2(new_n711), .A3(new_n712), .A4(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G29), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n716), .A2(KEYINPUT87), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n716), .A2(KEYINPUT87), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n708), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(G2067), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT98), .ZN(new_n722));
  NAND3_X1  g297(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT26), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n723), .A2(new_n724), .ZN(new_n726));
  AOI22_X1  g301(.A1(new_n725), .A2(new_n726), .B1(G105), .B2(new_n479), .ZN(new_n727));
  INV_X1    g302(.A(G141), .ZN(new_n728));
  INV_X1    g303(.A(G129), .ZN(new_n729));
  OAI221_X1 g304(.A(new_n727), .B1(new_n468), .B2(new_n728), .C1(new_n729), .C2(new_n487), .ZN(new_n730));
  MUX2_X1   g305(.A(G32), .B(new_n730), .S(G29), .Z(new_n731));
  XOR2_X1   g306(.A(KEYINPUT27), .B(G1996), .Z(new_n732));
  INV_X1    g307(.A(KEYINPUT24), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n683), .B1(new_n733), .B2(G34), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT91), .ZN(new_n735));
  AOI22_X1  g310(.A1(new_n734), .A2(new_n735), .B1(new_n733), .B2(G34), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(new_n735), .B2(new_n734), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(new_n481), .B2(new_n683), .ZN(new_n738));
  INV_X1    g313(.A(G2084), .ZN(new_n739));
  AOI22_X1  g314(.A1(new_n731), .A2(new_n732), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(new_n702), .B2(G1961), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n704), .B(new_n721), .C1(new_n722), .C2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(G168), .A2(G16), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT93), .ZN(new_n744));
  INV_X1    g319(.A(G21), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n744), .B1(new_n662), .B2(new_n745), .ZN(new_n746));
  XOR2_X1   g321(.A(KEYINPUT94), .B(G1966), .Z(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n683), .A2(G35), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G162), .B2(new_n683), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT29), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(G2090), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n662), .A2(G19), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT83), .Z(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(new_n549), .B2(new_n662), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT84), .B(KEYINPUT85), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  OAI211_X1 g332(.A(new_n748), .B(new_n752), .C1(G1341), .C2(new_n757), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n741), .B2(new_n722), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT23), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n662), .A2(G20), .ZN(new_n761));
  AOI211_X1 g336(.A(new_n760), .B(new_n761), .C1(G299), .C2(G16), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n760), .B2(new_n761), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G1956), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n683), .A2(G27), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G164), .B2(new_n683), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G2078), .ZN(new_n767));
  INV_X1    g342(.A(G33), .ZN(new_n768));
  INV_X1    g343(.A(G2072), .ZN(new_n769));
  AOI22_X1  g344(.A1(new_n683), .A2(new_n768), .B1(new_n769), .B2(KEYINPUT92), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n479), .A2(G103), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT25), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G139), .B2(new_n469), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n498), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT90), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n461), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n775), .B2(new_n774), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n773), .A2(new_n777), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n770), .B1(new_n778), .B2(new_n683), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n769), .A2(KEYINPUT92), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n779), .B(new_n780), .Z(new_n781));
  NOR3_X1   g356(.A1(new_n764), .A2(new_n767), .A3(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n751), .A2(G2090), .ZN(new_n783));
  NOR2_X1   g358(.A1(G4), .A2(G16), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT82), .Z(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(new_n581), .B2(new_n662), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G1348), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n731), .A2(new_n732), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n738), .A2(new_n739), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n607), .A2(G29), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT31), .B(G11), .ZN(new_n791));
  INV_X1    g366(.A(G28), .ZN(new_n792));
  NOR3_X1   g367(.A1(new_n792), .A2(KEYINPUT95), .A3(KEYINPUT30), .ZN(new_n793));
  OAI21_X1  g368(.A(KEYINPUT95), .B1(new_n792), .B2(KEYINPUT30), .ZN(new_n794));
  AOI21_X1  g369(.A(G29), .B1(new_n792), .B2(KEYINPUT30), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  OAI211_X1 g371(.A(new_n790), .B(new_n791), .C1(new_n793), .C2(new_n796), .ZN(new_n797));
  NOR3_X1   g372(.A1(new_n788), .A2(new_n789), .A3(new_n797), .ZN(new_n798));
  OAI211_X1 g373(.A(new_n787), .B(new_n798), .C1(new_n746), .C2(new_n747), .ZN(new_n799));
  AOI211_X1 g374(.A(new_n783), .B(new_n799), .C1(G1341), .C2(new_n757), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n759), .A2(new_n782), .A3(new_n800), .ZN(new_n801));
  NOR3_X1   g376(.A1(new_n699), .A2(new_n742), .A3(new_n801), .ZN(G311));
  INV_X1    g377(.A(G311), .ZN(G150));
  XNOR2_X1  g378(.A(KEYINPUT101), .B(G860), .ZN(new_n804));
  AOI22_X1  g379(.A1(new_n518), .A2(G93), .B1(G55), .B2(new_n547), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n528), .A2(G67), .ZN(new_n806));
  NAND2_X1  g381(.A1(G80), .A2(G543), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n806), .A2(KEYINPUT99), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n808), .A2(G651), .ZN(new_n809));
  AOI21_X1  g384(.A(KEYINPUT99), .B1(new_n806), .B2(new_n807), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n805), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT100), .ZN(new_n812));
  AND2_X1   g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n549), .B1(new_n811), .B2(new_n812), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n813), .A2(new_n814), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n582), .A2(G559), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n804), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(new_n821), .B2(new_n820), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n811), .A2(new_n804), .ZN(new_n824));
  XOR2_X1   g399(.A(KEYINPUT102), .B(KEYINPUT37), .Z(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n823), .A2(new_n826), .ZN(G145));
  NAND2_X1  g402(.A1(new_n488), .A2(G130), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n469), .A2(G142), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n461), .A2(G118), .ZN(new_n830));
  OAI21_X1  g405(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n831));
  OAI211_X1 g406(.A(new_n828), .B(new_n829), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n690), .B(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT105), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(new_n597), .Z(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT106), .Z(new_n836));
  INV_X1    g411(.A(new_n493), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT103), .ZN(new_n838));
  AND3_X1   g413(.A1(new_n502), .A2(new_n838), .A3(new_n503), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n838), .B1(new_n502), .B2(new_n503), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n837), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(new_n730), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(new_n715), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT104), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n778), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n773), .A2(new_n777), .A3(KEYINPUT104), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n843), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(new_n845), .B2(new_n843), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n836), .B(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n481), .B(new_n607), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(G162), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(G37), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n851), .B1(new_n836), .B2(new_n848), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT107), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n848), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n848), .A2(new_n855), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(new_n835), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n854), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n852), .A2(new_n853), .A3(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g436(.A(G303), .B(new_n669), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n674), .B(G290), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n864), .B(KEYINPUT108), .Z(new_n865));
  NAND2_X1  g440(.A1(new_n862), .A2(new_n863), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n866), .B(KEYINPUT109), .Z(new_n867));
  NOR2_X1   g442(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT42), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n592), .B(new_n817), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n581), .B(G299), .Z(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n871), .B(KEYINPUT41), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n872), .B1(new_n870), .B2(new_n873), .ZN(new_n874));
  AND2_X1   g449(.A1(new_n869), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n869), .A2(new_n874), .ZN(new_n876));
  OAI21_X1  g451(.A(G868), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n811), .A2(new_n585), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(G331));
  INV_X1    g454(.A(KEYINPUT110), .ZN(new_n880));
  XNOR2_X1  g455(.A(G331), .B(new_n880), .ZN(G295));
  INV_X1    g456(.A(KEYINPUT44), .ZN(new_n882));
  INV_X1    g457(.A(new_n817), .ZN(new_n883));
  AOI21_X1  g458(.A(G171), .B1(G286), .B2(KEYINPUT112), .ZN(new_n884));
  NOR2_X1   g459(.A1(G286), .A2(KEYINPUT112), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n884), .B(new_n885), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n883), .A2(new_n886), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n887), .A2(new_n871), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n873), .B1(new_n887), .B2(new_n888), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n868), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(new_n853), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT113), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OR3_X1    g469(.A1(new_n889), .A2(new_n890), .A3(new_n868), .ZN(new_n895));
  XOR2_X1   g470(.A(KEYINPUT111), .B(KEYINPUT43), .Z(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n891), .A2(KEYINPUT113), .A3(new_n853), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n894), .A2(new_n895), .A3(new_n897), .A4(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n895), .A2(new_n891), .A3(new_n853), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(KEYINPUT43), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n882), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n900), .A2(new_n896), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n894), .A2(new_n895), .A3(new_n898), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n903), .B1(new_n904), .B2(new_n896), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n902), .B1(new_n882), .B2(new_n905), .ZN(G397));
  INV_X1    g481(.A(G1384), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n841), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT45), .ZN(new_n909));
  NAND2_X1  g484(.A1(G160), .A2(G40), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  AND3_X1   g486(.A1(new_n908), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  XOR2_X1   g487(.A(new_n912), .B(KEYINPUT114), .Z(new_n913));
  OR2_X1    g488(.A1(new_n691), .A2(new_n693), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n715), .B(new_n720), .ZN(new_n915));
  INV_X1    g490(.A(G1996), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n730), .B(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n691), .A2(new_n693), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n914), .A2(new_n915), .A3(new_n917), .A4(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(G290), .B(G1986), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n913), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT122), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT51), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT50), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n494), .B1(new_n469), .B2(G138), .ZN(new_n925));
  OAI21_X1  g500(.A(KEYINPUT68), .B1(new_n474), .B2(new_n495), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n498), .A2(new_n497), .A3(new_n500), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(KEYINPUT103), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n502), .A2(new_n838), .A3(new_n503), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n493), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NOR3_X1   g506(.A1(new_n931), .A2(KEYINPUT115), .A3(G1384), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT115), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n933), .B1(new_n841), .B2(new_n907), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n924), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT116), .ZN(new_n936));
  NOR2_X1   g511(.A1(G164), .A2(G1384), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n936), .B1(new_n937), .B2(new_n924), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n837), .B1(new_n925), .B2(new_n928), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(new_n907), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n940), .A2(KEYINPUT116), .A3(KEYINPUT50), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n938), .A2(new_n941), .A3(new_n911), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  XOR2_X1   g518(.A(KEYINPUT118), .B(G2084), .Z(new_n944));
  NAND3_X1  g519(.A1(new_n935), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(KEYINPUT119), .ZN(new_n946));
  OAI21_X1  g521(.A(KEYINPUT115), .B1(new_n931), .B2(G1384), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n841), .A2(new_n933), .A3(new_n907), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n942), .B1(new_n949), .B2(new_n924), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT119), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n950), .A2(new_n951), .A3(new_n944), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n947), .A2(new_n909), .A3(new_n948), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n910), .B1(KEYINPUT45), .B2(new_n937), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n747), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n946), .A2(new_n952), .A3(new_n957), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n923), .B(G8), .C1(new_n958), .C2(G286), .ZN(new_n959));
  INV_X1    g534(.A(G8), .ZN(new_n960));
  NOR2_X1   g535(.A1(G168), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n958), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  AOI211_X1 g538(.A(new_n923), .B(new_n961), .C1(new_n958), .C2(G8), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n922), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n958), .A2(G8), .ZN(new_n966));
  OAI211_X1 g541(.A(new_n966), .B(KEYINPUT51), .C1(new_n960), .C2(G168), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n967), .A2(KEYINPUT122), .A3(new_n962), .A4(new_n959), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(KEYINPUT62), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT62), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n965), .A2(new_n968), .A3(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT52), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n910), .B1(new_n947), .B2(new_n948), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n974), .A2(new_n960), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n674), .A2(G1976), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n973), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n974), .ZN(new_n979));
  NAND2_X1  g554(.A1(G305), .A2(G1981), .ZN(new_n980));
  INV_X1    g555(.A(G1981), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n669), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n983), .B(KEYINPUT49), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n979), .A2(new_n984), .A3(G8), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n973), .B1(new_n674), .B2(G1976), .ZN(new_n986));
  NOR4_X1   g561(.A1(new_n974), .A2(new_n960), .A3(new_n976), .A4(new_n986), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n978), .A2(new_n985), .A3(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G2090), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n950), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n841), .A2(KEYINPUT45), .A3(new_n907), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n940), .A2(new_n909), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n991), .A2(new_n911), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(new_n665), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n960), .B1(new_n990), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT55), .ZN(new_n996));
  NOR3_X1   g571(.A1(G166), .A2(new_n996), .A3(new_n960), .ZN(new_n997));
  AOI21_X1  g572(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n995), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n947), .A2(KEYINPUT50), .A3(new_n948), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT117), .B1(new_n937), .B2(new_n924), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT117), .ZN(new_n1004));
  NOR4_X1   g579(.A1(G164), .A2(new_n1004), .A3(KEYINPUT50), .A4(G1384), .ZN(new_n1005));
  NOR3_X1   g580(.A1(new_n1003), .A2(new_n910), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1002), .A2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n994), .B1(new_n1007), .B2(G2090), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(G8), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(new_n999), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n988), .A2(new_n1001), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(G1961), .ZN(new_n1012));
  AOI21_X1  g587(.A(KEYINPUT50), .B1(new_n947), .B2(new_n948), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1012), .B1(new_n1013), .B2(new_n942), .ZN(new_n1014));
  INV_X1    g589(.A(G2078), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n991), .A2(new_n1015), .A3(new_n911), .A4(new_n992), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT53), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n953), .A2(KEYINPUT53), .A3(new_n1015), .A4(new_n954), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1014), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(G171), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1011), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n970), .A2(new_n972), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n975), .A2(new_n984), .ZN(new_n1024));
  NOR2_X1   g599(.A1(G288), .A2(G1976), .ZN(new_n1025));
  AOI22_X1  g600(.A1(new_n1024), .A2(new_n1025), .B1(new_n981), .B2(new_n669), .ZN(new_n1026));
  INV_X1    g601(.A(new_n975), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1001), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1028), .B1(new_n1029), .B2(new_n988), .ZN(new_n1030));
  XNOR2_X1  g605(.A(KEYINPUT120), .B(KEYINPUT63), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  AND3_X1   g607(.A1(new_n988), .A2(new_n1001), .A3(new_n1010), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n958), .A2(G8), .A3(G168), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1032), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n988), .A2(new_n1001), .ZN(new_n1037));
  OAI21_X1  g612(.A(KEYINPUT63), .B1(new_n995), .B2(new_n1000), .ZN(new_n1038));
  NOR3_X1   g613(.A1(new_n1037), .A2(new_n1038), .A3(new_n1034), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1030), .B1(new_n1036), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT125), .ZN(new_n1041));
  XNOR2_X1  g616(.A(KEYINPUT123), .B(KEYINPUT54), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1017), .B1(new_n908), .B2(new_n909), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1043), .A2(new_n1015), .A3(new_n911), .A4(new_n991), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1014), .A2(G301), .A3(new_n1018), .A4(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(KEYINPUT124), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(new_n1021), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1045), .A2(KEYINPUT124), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1041), .B(new_n1042), .C1(new_n1047), .C2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1042), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(KEYINPUT125), .ZN(new_n1051));
  XNOR2_X1  g626(.A(G299), .B(KEYINPUT57), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(G1956), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1007), .A2(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g630(.A(KEYINPUT56), .B(G2072), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n993), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1053), .B1(new_n1055), .B2(new_n1059), .ZN(new_n1060));
  AOI211_X1 g635(.A(G2067), .B(new_n910), .C1(new_n947), .C2(new_n948), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n935), .A2(new_n943), .ZN(new_n1062));
  INV_X1    g637(.A(G1348), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1061), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1064), .A2(new_n581), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1055), .A2(new_n1053), .A3(new_n1059), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1060), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT61), .ZN(new_n1068));
  AOI21_X1  g643(.A(G1956), .B1(new_n1002), .B2(new_n1006), .ZN(new_n1069));
  NOR3_X1   g644(.A1(new_n1069), .A2(new_n1058), .A3(new_n1052), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1068), .B1(new_n1060), .B2(new_n1070), .ZN(new_n1071));
  XNOR2_X1  g646(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n1072));
  XNOR2_X1  g647(.A(new_n1072), .B(G1341), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n974), .A2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n993), .A2(G1996), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n549), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(KEYINPUT59), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT59), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1079), .B(new_n549), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1071), .A2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1052), .B1(new_n1069), .B2(new_n1058), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1066), .A2(KEYINPUT61), .A3(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT60), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n581), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n581), .A2(new_n1085), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1086), .B1(new_n1064), .B2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1063), .B1(new_n1013), .B2(new_n942), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n974), .A2(new_n720), .ZN(new_n1090));
  AND4_X1   g665(.A1(KEYINPUT60), .A2(new_n1089), .A3(new_n582), .A4(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1084), .B1(new_n1088), .B2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1067), .B1(new_n1082), .B2(new_n1092), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n1014), .A2(new_n1018), .A3(new_n1044), .ZN(new_n1094));
  OAI21_X1  g669(.A(KEYINPUT54), .B1(new_n1094), .B2(G301), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1020), .A2(G171), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1097), .A2(new_n1011), .ZN(new_n1098));
  AND4_X1   g673(.A1(new_n1049), .A2(new_n1051), .A3(new_n1093), .A4(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1040), .B1(new_n1099), .B2(new_n969), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1023), .B1(new_n1100), .B2(KEYINPUT126), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1030), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1039), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1031), .B1(new_n1011), .B2(new_n1034), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1102), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n969), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1051), .A2(new_n1093), .A3(new_n1098), .A4(new_n1049), .ZN(new_n1107));
  OAI211_X1 g682(.A(KEYINPUT126), .B(new_n1105), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n921), .B1(new_n1101), .B2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g685(.A1(G290), .A2(G1986), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n913), .A2(new_n1111), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1112), .A2(KEYINPUT48), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1112), .A2(KEYINPUT48), .ZN(new_n1114));
  AOI211_X1 g689(.A(new_n1113), .B(new_n1114), .C1(new_n913), .C2(new_n919), .ZN(new_n1115));
  AND2_X1   g690(.A1(new_n913), .A2(new_n916), .ZN(new_n1116));
  OR2_X1    g691(.A1(new_n1116), .A2(KEYINPUT46), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(KEYINPUT46), .ZN(new_n1118));
  INV_X1    g693(.A(new_n915), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n913), .B1(new_n730), .B2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1117), .A2(new_n1118), .A3(new_n1120), .ZN(new_n1121));
  XOR2_X1   g696(.A(new_n1121), .B(KEYINPUT47), .Z(new_n1122));
  NAND2_X1  g697(.A1(new_n915), .A2(new_n917), .ZN(new_n1123));
  OAI22_X1  g698(.A1(new_n1123), .A2(new_n918), .B1(G2067), .B2(new_n715), .ZN(new_n1124));
  AOI211_X1 g699(.A(new_n1115), .B(new_n1122), .C1(new_n913), .C2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1110), .A2(new_n1125), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g701(.A(G319), .ZN(new_n1128));
  NOR4_X1   g702(.A1(G229), .A2(new_n1128), .A3(G401), .A4(G227), .ZN(new_n1129));
  XNOR2_X1  g703(.A(new_n1129), .B(KEYINPUT127), .ZN(new_n1130));
  NAND2_X1  g704(.A1(new_n860), .A2(new_n1130), .ZN(new_n1131));
  NOR2_X1   g705(.A1(new_n905), .A2(new_n1131), .ZN(G308));
  OR2_X1    g706(.A1(new_n905), .A2(new_n1131), .ZN(G225));
endmodule


