//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 0 0 0 1 0 0 0 0 1 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 1 0 0 1 1 0 1 1 0 1 0 1 1 0 1 1 1 0 0 0 0 1 0 0 1 0 0 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n771, new_n772, new_n773, new_n774, new_n776, new_n777, new_n778,
    new_n779, new_n781, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n861, new_n862, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n979, new_n980, new_n981,
    new_n982;
  OAI21_X1  g000(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT14), .ZN(new_n203));
  INV_X1    g002(.A(G29gat), .ZN(new_n204));
  INV_X1    g003(.A(G36gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n203), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n206), .A2(KEYINPUT89), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT89), .ZN(new_n208));
  NOR2_X1   g007(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n208), .B1(new_n209), .B2(new_n205), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n202), .B1(new_n207), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT90), .ZN(new_n212));
  AOI22_X1  g011(.A1(new_n211), .A2(new_n212), .B1(G29gat), .B2(G36gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n213), .B1(new_n212), .B2(new_n211), .ZN(new_n214));
  INV_X1    g013(.A(G50gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G43gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT15), .ZN(new_n217));
  INV_X1    g016(.A(G43gat), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n217), .B1(new_n218), .B2(G50gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n214), .A2(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n219), .B1(G29gat), .B2(G36gat), .ZN(new_n221));
  AND2_X1   g020(.A1(new_n206), .A2(KEYINPUT92), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n206), .A2(KEYINPUT92), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n202), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT91), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n225), .B1(new_n215), .B2(G43gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n218), .A2(KEYINPUT91), .A3(G50gat), .ZN(new_n227));
  AND3_X1   g026(.A1(new_n226), .A2(new_n216), .A3(new_n227), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n221), .B(new_n224), .C1(KEYINPUT15), .C2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n220), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G15gat), .B(G22gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT16), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n231), .B1(new_n232), .B2(G1gat), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n233), .B1(G1gat), .B2(new_n231), .ZN(new_n234));
  INV_X1    g033(.A(G8gat), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n234), .B(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n230), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT93), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n230), .A2(KEYINPUT93), .A3(new_n237), .ZN(new_n241));
  INV_X1    g040(.A(new_n230), .ZN(new_n242));
  AOI22_X1  g041(.A1(new_n240), .A2(new_n241), .B1(new_n242), .B2(new_n236), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT96), .ZN(new_n244));
  NAND2_X1  g043(.A1(G229gat), .A2(G233gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n245), .B(KEYINPUT95), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n246), .B(KEYINPUT13), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  OR3_X1    g047(.A1(new_n243), .A2(new_n244), .A3(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n244), .B1(new_n243), .B2(new_n248), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n242), .A2(KEYINPUT17), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT17), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n230), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n252), .A2(new_n236), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n240), .A2(new_n241), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n255), .A2(new_n256), .A3(new_n245), .ZN(new_n257));
  AND3_X1   g056(.A1(new_n257), .A2(KEYINPUT94), .A3(KEYINPUT18), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT18), .B1(new_n257), .B2(KEYINPUT94), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n251), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n261));
  XNOR2_X1  g060(.A(G113gat), .B(G141gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n261), .B(new_n262), .ZN(new_n263));
  XOR2_X1   g062(.A(G169gat), .B(G197gat), .Z(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  XOR2_X1   g064(.A(new_n265), .B(KEYINPUT12), .Z(new_n266));
  NAND2_X1  g065(.A1(new_n260), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n266), .ZN(new_n268));
  OAI211_X1 g067(.A(new_n251), .B(new_n268), .C1(new_n258), .C2(new_n259), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT65), .ZN(new_n272));
  INV_X1    g071(.A(G183gat), .ZN(new_n273));
  INV_X1    g072(.A(G190gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n276));
  AOI21_X1  g075(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n275), .B(new_n276), .C1(new_n277), .C2(KEYINPUT64), .ZN(new_n278));
  AND2_X1   g077(.A1(new_n277), .A2(KEYINPUT64), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n272), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NOR2_X1   g079(.A1(G183gat), .A2(G190gat), .ZN(new_n281));
  AND2_X1   g080(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n281), .B1(new_n282), .B2(G190gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(G183gat), .A2(G190gat), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT24), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT64), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n277), .A2(KEYINPUT64), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n283), .A2(new_n288), .A3(KEYINPUT65), .A4(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(G169gat), .A2(G176gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT23), .ZN(new_n292));
  NAND2_X1  g091(.A1(G169gat), .A2(G176gat), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT23), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n294), .B1(G169gat), .B2(G176gat), .ZN(new_n295));
  AND3_X1   g094(.A1(new_n292), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n280), .A2(new_n290), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(KEYINPUT25), .ZN(new_n298));
  OAI21_X1  g097(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT66), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT66), .ZN(new_n301));
  OAI211_X1 g100(.A(new_n301), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n300), .A2(new_n302), .A3(new_n293), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT67), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT67), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n300), .A2(new_n305), .A3(new_n302), .A4(new_n293), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT26), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n304), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n273), .A2(KEYINPUT27), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT27), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(G183gat), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n310), .A2(new_n312), .A3(new_n274), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT28), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(KEYINPUT27), .B(G183gat), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n316), .A2(KEYINPUT28), .A3(new_n274), .ZN(new_n317));
  AOI22_X1  g116(.A1(new_n315), .A2(new_n317), .B1(G183gat), .B2(G190gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n309), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT25), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n286), .A2(new_n275), .A3(new_n276), .ZN(new_n321));
  AND3_X1   g120(.A1(new_n296), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n298), .A2(new_n319), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(G226gat), .A2(G233gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n325), .B(KEYINPUT72), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(G211gat), .A2(G218gat), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT22), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NOR2_X1   g129(.A1(G197gat), .A2(G204gat), .ZN(new_n331));
  AND2_X1   g130(.A1(G197gat), .A2(G204gat), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  XOR2_X1   g132(.A(G211gat), .B(G218gat), .Z(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(G211gat), .B(G218gat), .ZN(new_n336));
  XNOR2_X1  g135(.A(G197gat), .B(G204gat), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n336), .A2(new_n337), .A3(new_n330), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n327), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT73), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT29), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n324), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n342), .B1(new_n344), .B2(new_n325), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n322), .B1(new_n297), .B2(KEYINPUT25), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT29), .B1(new_n346), .B2(new_n319), .ZN(new_n347));
  INV_X1    g146(.A(new_n325), .ZN(new_n348));
  NOR3_X1   g147(.A1(new_n347), .A2(KEYINPUT73), .A3(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n341), .B1(new_n345), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n324), .A2(new_n348), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n351), .B1(new_n347), .B2(new_n326), .ZN(new_n352));
  INV_X1    g151(.A(new_n339), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(G8gat), .B(G36gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n355), .B(G64gat), .ZN(new_n356));
  INV_X1    g155(.A(G92gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n356), .B(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT30), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n350), .A2(new_n354), .A3(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n358), .B(KEYINPUT74), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n344), .A2(new_n342), .A3(new_n325), .ZN(new_n364));
  OAI21_X1  g163(.A(KEYINPUT73), .B1(new_n347), .B2(new_n348), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n340), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n326), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n344), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n339), .B1(new_n368), .B2(new_n351), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n363), .B1(new_n366), .B2(new_n369), .ZN(new_n370));
  AND2_X1   g169(.A1(new_n362), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n350), .A2(new_n354), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n360), .B1(new_n372), .B2(new_n359), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(G1gat), .B(G29gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n375), .B(KEYINPUT0), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n376), .B(G57gat), .ZN(new_n377));
  INV_X1    g176(.A(G85gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n377), .B(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT5), .ZN(new_n380));
  INV_X1    g179(.A(G113gat), .ZN(new_n381));
  INV_X1    g180(.A(G120gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT1), .ZN(new_n384));
  NAND2_X1  g183(.A1(G113gat), .A2(G120gat), .ZN(new_n385));
  AND3_X1   g184(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(G127gat), .A2(G134gat), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NOR2_X1   g187(.A1(G127gat), .A2(G134gat), .ZN(new_n389));
  OAI22_X1  g188(.A1(new_n388), .A2(new_n389), .B1(KEYINPUT68), .B2(KEYINPUT1), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n386), .A2(new_n390), .ZN(new_n391));
  NOR2_X1   g190(.A1(KEYINPUT68), .A2(KEYINPUT1), .ZN(new_n392));
  INV_X1    g191(.A(G127gat), .ZN(new_n393));
  INV_X1    g192(.A(G134gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n392), .B1(new_n395), .B2(new_n387), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT75), .ZN(new_n399));
  NAND2_X1  g198(.A1(G155gat), .A2(G162gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT2), .ZN(new_n401));
  INV_X1    g200(.A(G148gat), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n402), .A2(G141gat), .ZN(new_n403));
  INV_X1    g202(.A(G141gat), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n404), .A2(G148gat), .ZN(new_n405));
  OAI211_X1 g204(.A(new_n399), .B(new_n401), .C1(new_n403), .C2(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(G155gat), .B(G162gat), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n404), .A2(G148gat), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n402), .A2(G141gat), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT75), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n407), .B1(new_n412), .B2(new_n401), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n391), .B(new_n398), .C1(new_n409), .C2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n406), .A2(new_n408), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n412), .A2(new_n407), .A3(new_n401), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n386), .A2(new_n390), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n396), .A2(new_n397), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n415), .B(new_n416), .C1(new_n417), .C2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n414), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(G225gat), .A2(G233gat), .ZN(new_n421));
  XOR2_X1   g220(.A(new_n421), .B(KEYINPUT77), .Z(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT78), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n419), .A2(KEYINPUT4), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n391), .A2(new_n398), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT4), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n428), .A2(new_n429), .A3(new_n415), .A4(new_n416), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(KEYINPUT3), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n417), .A2(new_n418), .ZN(new_n434));
  XNOR2_X1  g233(.A(KEYINPUT76), .B(KEYINPUT3), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n415), .A2(new_n416), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n433), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n431), .A2(new_n422), .A3(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n380), .B1(new_n426), .B2(new_n438), .ZN(new_n439));
  AND2_X1   g238(.A1(new_n436), .A2(new_n434), .ZN(new_n440));
  AOI22_X1  g239(.A1(new_n433), .A2(new_n440), .B1(new_n427), .B2(new_n430), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n420), .A2(KEYINPUT78), .A3(new_n423), .ZN(new_n442));
  AOI22_X1  g241(.A1(new_n441), .A2(new_n422), .B1(new_n442), .B2(KEYINPUT5), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n379), .B1(new_n439), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n379), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n442), .A2(KEYINPUT5), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(new_n438), .ZN(new_n447));
  AOI21_X1  g246(.A(KEYINPUT78), .B1(new_n420), .B2(new_n423), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n448), .B1(new_n441), .B2(new_n422), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n445), .B(new_n447), .C1(new_n449), .C2(new_n380), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT6), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n444), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n439), .A2(new_n443), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n453), .A2(KEYINPUT6), .A3(new_n445), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n374), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(G227gat), .ZN(new_n458));
  INV_X1    g257(.A(G233gat), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n324), .A2(new_n428), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n346), .A2(new_n434), .A3(new_n319), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT34), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI211_X1 g264(.A(KEYINPUT34), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(G15gat), .B(G43gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(G71gat), .B(G99gat), .ZN(new_n470));
  XOR2_X1   g269(.A(new_n469), .B(new_n470), .Z(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n461), .A2(new_n460), .A3(new_n462), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT69), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT69), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n461), .A2(new_n475), .A3(new_n460), .A4(new_n462), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT32), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(KEYINPUT33), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n472), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  OR2_X1    g279(.A1(new_n471), .A2(KEYINPUT70), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT33), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n482), .B1(new_n471), .B2(KEYINPUT70), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n478), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n485), .B1(new_n474), .B2(new_n476), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n468), .B1(new_n480), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n477), .A2(new_n484), .ZN(new_n488));
  AOI22_X1  g287(.A1(new_n474), .A2(new_n476), .B1(new_n478), .B2(KEYINPUT33), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n488), .B(new_n467), .C1(new_n489), .C2(new_n472), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(G228gat), .A2(G233gat), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n333), .A2(new_n334), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n336), .B1(new_n330), .B2(new_n337), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n343), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  AOI22_X1  g295(.A1(new_n496), .A2(new_n435), .B1(new_n415), .B2(new_n416), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n339), .B1(new_n436), .B2(new_n343), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n493), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT80), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  OAI211_X1 g300(.A(KEYINPUT80), .B(new_n493), .C1(new_n497), .C2(new_n498), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT3), .ZN(new_n504));
  AOI21_X1  g303(.A(KEYINPUT29), .B1(new_n335), .B2(new_n338), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n504), .B1(new_n505), .B2(KEYINPUT81), .ZN(new_n506));
  AND3_X1   g305(.A1(new_n339), .A2(KEYINPUT81), .A3(new_n343), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n432), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT82), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT82), .ZN(new_n510));
  OAI211_X1 g309(.A(new_n510), .B(new_n432), .C1(new_n506), .C2(new_n507), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n498), .A2(new_n493), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n509), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(G22gat), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n503), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n514), .B1(new_n503), .B2(new_n513), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT83), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n503), .A2(new_n513), .A3(KEYINPUT83), .A4(new_n514), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(G78gat), .B(G106gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(KEYINPUT31), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(G50gat), .ZN(new_n523));
  XOR2_X1   g322(.A(new_n523), .B(KEYINPUT79), .Z(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n520), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n503), .A2(new_n513), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(G22gat), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n528), .A2(new_n515), .A3(new_n523), .ZN(new_n529));
  AOI21_X1  g328(.A(KEYINPUT84), .B1(new_n526), .B2(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n524), .B1(new_n518), .B2(new_n519), .ZN(new_n531));
  INV_X1    g330(.A(new_n529), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT84), .ZN(new_n533));
  NOR3_X1   g332(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n457), .B(new_n492), .C1(new_n530), .C2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT35), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n526), .A2(KEYINPUT84), .A3(new_n529), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n533), .B1(new_n531), .B2(new_n532), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT87), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT35), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n371), .A2(new_n455), .A3(new_n373), .A4(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n542), .A2(new_n491), .ZN(new_n543));
  AND3_X1   g342(.A1(new_n539), .A2(new_n540), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n540), .B1(new_n539), .B2(new_n543), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n536), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT38), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n363), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT37), .ZN(new_n549));
  AOI22_X1  g348(.A1(new_n344), .A2(new_n367), .B1(new_n324), .B2(new_n348), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n549), .B1(new_n550), .B2(new_n339), .ZN(new_n551));
  AOI22_X1  g350(.A1(new_n364), .A2(new_n365), .B1(new_n324), .B2(new_n326), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n551), .B1(new_n552), .B2(new_n339), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n549), .B1(new_n366), .B2(new_n369), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n548), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n372), .A2(new_n359), .ZN(new_n556));
  NOR3_X1   g355(.A1(new_n555), .A2(new_n455), .A3(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n554), .ZN(new_n558));
  NOR3_X1   g357(.A1(new_n366), .A2(new_n369), .A3(new_n549), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n359), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(KEYINPUT38), .ZN(new_n561));
  AOI22_X1  g360(.A1(new_n537), .A2(new_n538), .B1(new_n557), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n431), .A2(new_n437), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(new_n423), .ZN(new_n564));
  OAI21_X1  g363(.A(KEYINPUT85), .B1(new_n420), .B2(new_n423), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT85), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n414), .A2(new_n419), .A3(new_n566), .A4(new_n422), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n564), .A2(KEYINPUT39), .A3(new_n565), .A4(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT39), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n563), .A2(new_n569), .A3(new_n423), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n568), .A2(KEYINPUT40), .A3(new_n379), .A4(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n565), .A2(KEYINPUT39), .A3(new_n567), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n422), .B1(new_n431), .B2(new_n437), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n570), .B(new_n379), .C1(new_n572), .C2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT40), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AND3_X1   g375(.A1(new_n571), .A2(new_n576), .A3(new_n450), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n362), .A2(new_n370), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n364), .A2(new_n365), .ZN(new_n579));
  AOI22_X1  g378(.A1(new_n579), .A2(new_n341), .B1(new_n353), .B2(new_n352), .ZN(new_n580));
  AOI21_X1  g379(.A(KEYINPUT30), .B1(new_n580), .B2(new_n358), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n577), .B1(new_n578), .B2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT86), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI211_X1 g383(.A(new_n577), .B(KEYINPUT86), .C1(new_n578), .C2(new_n581), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n562), .A2(new_n586), .ZN(new_n587));
  OAI211_X1 g386(.A(new_n537), .B(new_n538), .C1(new_n456), .C2(new_n374), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT71), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT36), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(KEYINPUT71), .A2(KEYINPUT36), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n491), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n487), .A2(new_n490), .A3(new_n589), .A4(new_n590), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n587), .A2(new_n588), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n271), .B1(new_n546), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(G85gat), .A2(G92gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT100), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT7), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT100), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n599), .B(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(KEYINPUT7), .ZN(new_n605));
  NAND2_X1  g404(.A1(G99gat), .A2(G106gat), .ZN(new_n606));
  AOI22_X1  g405(.A1(KEYINPUT8), .A2(new_n606), .B1(new_n378), .B2(new_n357), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n602), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  XOR2_X1   g407(.A(G99gat), .B(G106gat), .Z(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT101), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n252), .A2(new_n254), .A3(new_n611), .ZN(new_n612));
  AND2_X1   g411(.A1(G232gat), .A2(G233gat), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(KEYINPUT41), .ZN(new_n614));
  OAI211_X1 g413(.A(new_n612), .B(new_n614), .C1(new_n242), .C2(new_n611), .ZN(new_n615));
  XOR2_X1   g414(.A(G134gat), .B(G162gat), .Z(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n613), .A2(KEYINPUT41), .ZN(new_n618));
  XNOR2_X1  g417(.A(G190gat), .B(G218gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n617), .B(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  XOR2_X1   g421(.A(G57gat), .B(G64gat), .Z(new_n623));
  INV_X1    g422(.A(G71gat), .ZN(new_n624));
  INV_X1    g423(.A(G78gat), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n623), .B1(KEYINPUT9), .B2(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(G71gat), .B(G78gat), .ZN(new_n628));
  XOR2_X1   g427(.A(new_n627), .B(new_n628), .Z(new_n629));
  INV_X1    g428(.A(KEYINPUT21), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(G231gat), .A2(G233gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(KEYINPUT20), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n236), .B1(new_n629), .B2(new_n630), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(new_n273), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n634), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g436(.A(KEYINPUT97), .B(KEYINPUT19), .Z(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(KEYINPUT98), .ZN(new_n639));
  XNOR2_X1  g438(.A(G127gat), .B(G155gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XOR2_X1   g440(.A(KEYINPUT99), .B(G211gat), .Z(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n637), .B(new_n643), .Z(new_n644));
  NAND2_X1  g443(.A1(new_n622), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT102), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n629), .B1(new_n610), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n610), .A2(new_n646), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n649), .A2(KEYINPUT10), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT10), .ZN(new_n651));
  NOR3_X1   g450(.A1(new_n611), .A2(new_n651), .A3(new_n629), .ZN(new_n652));
  INV_X1    g451(.A(G230gat), .ZN(new_n653));
  OAI22_X1  g452(.A1(new_n650), .A2(new_n652), .B1(new_n653), .B2(new_n459), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n653), .A2(new_n459), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n649), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(G120gat), .B(G148gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(G176gat), .ZN(new_n658));
  XOR2_X1   g457(.A(new_n658), .B(G204gat), .Z(new_n659));
  NAND3_X1  g458(.A1(new_n654), .A2(new_n656), .A3(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n659), .B1(new_n654), .B2(new_n656), .ZN(new_n662));
  OAI21_X1  g461(.A(KEYINPUT103), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n662), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT103), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n664), .A2(new_n665), .A3(new_n660), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n645), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n598), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n669), .A2(new_n455), .ZN(new_n670));
  XOR2_X1   g469(.A(new_n670), .B(G1gat), .Z(G1324gat));
  INV_X1    g470(.A(new_n374), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g472(.A(KEYINPUT16), .B(G8gat), .Z(new_n674));
  AND2_X1   g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OR2_X1    g474(.A1(new_n675), .A2(KEYINPUT42), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(KEYINPUT42), .ZN(new_n677));
  OAI211_X1 g476(.A(new_n676), .B(new_n677), .C1(new_n235), .C2(new_n673), .ZN(G1325gat));
  OAI21_X1  g477(.A(G15gat), .B1(new_n669), .B2(new_n596), .ZN(new_n679));
  OR2_X1    g478(.A1(new_n491), .A2(G15gat), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n679), .B1(new_n669), .B2(new_n680), .ZN(G1326gat));
  NOR2_X1   g480(.A1(new_n669), .A2(new_n539), .ZN(new_n682));
  XOR2_X1   g481(.A(KEYINPUT43), .B(G22gat), .Z(new_n683));
  XNOR2_X1  g482(.A(new_n682), .B(new_n683), .ZN(G1327gat));
  OAI21_X1  g483(.A(new_n543), .B1(new_n530), .B2(new_n534), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(KEYINPUT87), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n539), .A2(new_n540), .A3(new_n543), .ZN(new_n687));
  AOI22_X1  g486(.A1(new_n686), .A2(new_n687), .B1(KEYINPUT35), .B2(new_n535), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n557), .A2(new_n561), .ZN(new_n689));
  AND3_X1   g488(.A1(new_n586), .A2(new_n539), .A3(new_n689), .ZN(new_n690));
  OAI211_X1 g489(.A(new_n594), .B(new_n593), .C1(new_n539), .C2(new_n457), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n621), .B1(new_n688), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(KEYINPUT104), .B1(new_n690), .B2(new_n691), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT104), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n587), .A2(new_n596), .A3(new_n695), .A4(new_n588), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n694), .A2(new_n546), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(KEYINPUT105), .B(KEYINPUT44), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n622), .A2(new_n698), .ZN(new_n699));
  AOI22_X1  g498(.A1(new_n693), .A2(KEYINPUT44), .B1(new_n697), .B2(new_n699), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n667), .A2(new_n644), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(new_n270), .ZN(new_n702));
  OAI21_X1  g501(.A(KEYINPUT106), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT106), .ZN(new_n704));
  INV_X1    g503(.A(new_n702), .ZN(new_n705));
  INV_X1    g504(.A(new_n699), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n686), .A2(new_n687), .ZN(new_n707));
  INV_X1    g506(.A(new_n691), .ZN(new_n708));
  AOI21_X1  g507(.A(KEYINPUT104), .B1(new_n562), .B2(new_n586), .ZN(new_n709));
  AOI22_X1  g508(.A1(new_n707), .A2(new_n536), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n706), .B1(new_n710), .B2(new_n694), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n546), .A2(new_n597), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n712), .B1(new_n713), .B2(new_n621), .ZN(new_n714));
  OAI211_X1 g513(.A(new_n704), .B(new_n705), .C1(new_n711), .C2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n703), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(G29gat), .B1(new_n716), .B2(new_n455), .ZN(new_n717));
  AND3_X1   g516(.A1(new_n598), .A2(new_n621), .A3(new_n701), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n718), .A2(new_n204), .A3(new_n456), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT45), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT107), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n717), .A2(KEYINPUT107), .A3(new_n720), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(G1328gat));
  OAI21_X1  g524(.A(G36gat), .B1(new_n716), .B2(new_n672), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n718), .A2(new_n205), .A3(new_n374), .ZN(new_n727));
  AND2_X1   g526(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n728));
  NOR2_X1   g527(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n726), .B(new_n730), .C1(new_n728), .C2(new_n727), .ZN(G1329gat));
  NOR2_X1   g530(.A1(new_n491), .A2(G43gat), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n718), .A2(new_n732), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n700), .A2(new_n596), .A3(new_n702), .ZN(new_n734));
  OAI211_X1 g533(.A(KEYINPUT47), .B(new_n733), .C1(new_n734), .C2(new_n218), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n703), .A2(new_n595), .A3(new_n715), .ZN(new_n736));
  AOI22_X1  g535(.A1(new_n736), .A2(G43gat), .B1(new_n718), .B2(new_n732), .ZN(new_n737));
  XNOR2_X1  g536(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n735), .B1(new_n737), .B2(new_n738), .ZN(G1330gat));
  INV_X1    g538(.A(new_n539), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n703), .A2(new_n740), .A3(new_n715), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(G50gat), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n539), .A2(G50gat), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n718), .A2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT48), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n742), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT111), .ZN(new_n749));
  OAI211_X1 g548(.A(new_n740), .B(new_n705), .C1(new_n711), .C2(new_n714), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT110), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n215), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n693), .A2(KEYINPUT44), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n697), .A2(new_n699), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n755), .A2(KEYINPUT110), .A3(new_n740), .A4(new_n705), .ZN(new_n756));
  AOI22_X1  g555(.A1(new_n752), .A2(new_n756), .B1(new_n718), .B2(new_n743), .ZN(new_n757));
  OAI211_X1 g556(.A(new_n748), .B(new_n749), .C1(new_n745), .C2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n750), .A2(new_n751), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n759), .A2(G50gat), .A3(new_n756), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n745), .B1(new_n760), .B2(new_n744), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n746), .B1(new_n741), .B2(G50gat), .ZN(new_n762));
  OAI21_X1  g561(.A(KEYINPUT111), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n758), .A2(new_n763), .ZN(G1331gat));
  INV_X1    g563(.A(new_n667), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n645), .A2(new_n270), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n697), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(new_n456), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g569(.A1(new_n767), .A2(new_n672), .ZN(new_n771));
  NOR2_X1   g570(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n772));
  AND2_X1   g571(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n771), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n774), .B1(new_n771), .B2(new_n772), .ZN(G1333gat));
  OAI21_X1  g574(.A(G71gat), .B1(new_n767), .B2(new_n596), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n492), .A2(new_n624), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n776), .B1(new_n767), .B2(new_n777), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(KEYINPUT112), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g579(.A1(new_n767), .A2(new_n539), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(new_n625), .ZN(G1335gat));
  INV_X1    g581(.A(new_n644), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n271), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n784), .A2(new_n765), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n755), .A2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(G85gat), .B1(new_n786), .B2(new_n455), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n784), .A2(new_n622), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n697), .A2(new_n788), .ZN(new_n789));
  OR2_X1    g588(.A1(new_n789), .A2(KEYINPUT51), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(KEYINPUT51), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n790), .A2(new_n667), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n456), .A2(new_n378), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n787), .B1(new_n792), .B2(new_n793), .ZN(G1336gat));
  NOR3_X1   g593(.A1(new_n792), .A2(G92gat), .A3(new_n672), .ZN(new_n795));
  INV_X1    g594(.A(new_n786), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n357), .B1(new_n796), .B2(new_n374), .ZN(new_n797));
  OR3_X1    g596(.A1(new_n795), .A2(new_n797), .A3(KEYINPUT52), .ZN(new_n798));
  OAI21_X1  g597(.A(KEYINPUT52), .B1(new_n795), .B2(new_n797), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(G1337gat));
  NAND3_X1  g599(.A1(new_n796), .A2(G99gat), .A3(new_n595), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n792), .A2(new_n491), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n801), .B1(new_n802), .B2(G99gat), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n803), .B(KEYINPUT113), .ZN(G1338gat));
  INV_X1    g603(.A(KEYINPUT53), .ZN(new_n805));
  OAI21_X1  g604(.A(G106gat), .B1(new_n786), .B2(new_n539), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT114), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n539), .A2(G106gat), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n790), .A2(new_n667), .A3(new_n791), .A4(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n806), .A2(new_n807), .A3(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n807), .B1(new_n806), .B2(new_n809), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n805), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n806), .A2(new_n809), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(KEYINPUT114), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n815), .A2(KEYINPUT53), .A3(new_n810), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n813), .A2(new_n816), .ZN(G1339gat));
  NOR3_X1   g616(.A1(new_n645), .A2(new_n667), .A3(new_n270), .ZN(new_n818));
  INV_X1    g617(.A(new_n648), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n819), .B(new_n647), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n651), .ZN(new_n821));
  INV_X1    g620(.A(new_n652), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n655), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n659), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n821), .A2(new_n655), .A3(new_n822), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n654), .A2(new_n826), .A3(KEYINPUT54), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n825), .A2(new_n827), .A3(KEYINPUT55), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n660), .ZN(new_n829));
  AOI21_X1  g628(.A(KEYINPUT55), .B1(new_n825), .B2(new_n827), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n243), .A2(new_n248), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n245), .B1(new_n255), .B2(new_n256), .ZN(new_n833));
  OAI211_X1 g632(.A(KEYINPUT115), .B(new_n265), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n265), .B1(new_n832), .B2(new_n833), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT115), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AND3_X1   g636(.A1(new_n269), .A2(new_n834), .A3(new_n837), .ZN(new_n838));
  AOI22_X1  g637(.A1(new_n270), .A2(new_n831), .B1(new_n667), .B2(new_n838), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n837), .A2(new_n834), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT116), .ZN(new_n841));
  AND3_X1   g640(.A1(new_n840), .A2(new_n841), .A3(new_n269), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n841), .B1(new_n840), .B2(new_n269), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n831), .A2(new_n621), .ZN(new_n845));
  OAI22_X1  g644(.A1(new_n839), .A2(new_n621), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n818), .B1(new_n846), .B2(new_n783), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n847), .A2(new_n740), .A3(new_n491), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n374), .A2(new_n455), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n850), .A2(new_n381), .A3(new_n271), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n847), .A2(new_n455), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n740), .A2(new_n491), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n854), .A2(new_n374), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n270), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n851), .B1(new_n856), .B2(new_n381), .ZN(G1340gat));
  NOR3_X1   g656(.A1(new_n850), .A2(new_n382), .A3(new_n765), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n855), .A2(new_n667), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n858), .B1(new_n859), .B2(new_n382), .ZN(G1341gat));
  NAND3_X1  g659(.A1(new_n855), .A2(new_n393), .A3(new_n644), .ZN(new_n861));
  OAI21_X1  g660(.A(G127gat), .B1(new_n850), .B2(new_n783), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(G1342gat));
  NOR2_X1   g662(.A1(new_n622), .A2(new_n374), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(new_n394), .ZN(new_n865));
  OR3_X1    g664(.A1(new_n854), .A2(KEYINPUT56), .A3(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(G134gat), .B1(new_n850), .B2(new_n622), .ZN(new_n867));
  OAI21_X1  g666(.A(KEYINPUT56), .B1(new_n854), .B2(new_n865), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(G1343gat));
  NOR2_X1   g668(.A1(new_n844), .A2(new_n845), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n831), .A2(new_n270), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n667), .A2(new_n838), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n621), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n783), .B1(new_n870), .B2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(new_n818), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT57), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n876), .A2(new_n877), .A3(new_n740), .ZN(new_n878));
  OAI21_X1  g677(.A(KEYINPUT57), .B1(new_n847), .B2(new_n539), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n596), .A2(new_n849), .ZN(new_n880));
  XNOR2_X1  g679(.A(new_n880), .B(KEYINPUT117), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n878), .A2(new_n879), .A3(new_n270), .A4(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(G141gat), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n595), .A2(new_n539), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n852), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n271), .A2(G141gat), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n885), .A2(new_n672), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n883), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(KEYINPUT58), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT58), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n883), .A2(new_n887), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n889), .A2(new_n891), .ZN(G1344gat));
  AND2_X1   g691(.A1(new_n885), .A2(new_n672), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n893), .A2(new_n402), .A3(new_n667), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT59), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n878), .A2(new_n879), .A3(new_n667), .A4(new_n881), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n895), .B1(new_n896), .B2(G148gat), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n896), .A2(new_n895), .A3(G148gat), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n894), .B1(new_n897), .B2(new_n898), .ZN(G1345gat));
  INV_X1    g698(.A(G155gat), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n893), .A2(new_n900), .A3(new_n644), .ZN(new_n901));
  AND4_X1   g700(.A1(new_n644), .A2(new_n878), .A3(new_n879), .A4(new_n881), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n901), .B1(new_n900), .B2(new_n902), .ZN(G1346gat));
  INV_X1    g702(.A(G162gat), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n878), .A2(new_n879), .A3(new_n621), .A4(new_n881), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT118), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n904), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n907), .B1(new_n906), .B2(new_n905), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n885), .A2(new_n904), .A3(new_n864), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(G1347gat));
  NOR3_X1   g709(.A1(new_n740), .A2(new_n672), .A3(new_n491), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n876), .A2(new_n455), .A3(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT119), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n876), .A2(KEYINPUT119), .A3(new_n455), .A4(new_n911), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n271), .A2(G169gat), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n672), .A2(new_n456), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n848), .A2(new_n270), .A3(new_n918), .ZN(new_n919));
  AND3_X1   g718(.A1(new_n919), .A2(KEYINPUT120), .A3(G169gat), .ZN(new_n920));
  AOI21_X1  g719(.A(KEYINPUT120), .B1(new_n919), .B2(G169gat), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n917), .B1(new_n920), .B2(new_n921), .ZN(G1348gat));
  NOR2_X1   g721(.A1(new_n765), .A2(G176gat), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n914), .A2(new_n915), .A3(new_n923), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n876), .A2(new_n853), .A3(new_n918), .ZN(new_n925));
  OAI21_X1  g724(.A(G176gat), .B1(new_n925), .B2(new_n765), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT121), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n924), .A2(KEYINPUT121), .A3(new_n926), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(G1349gat));
  OAI21_X1  g730(.A(G183gat), .B1(new_n925), .B2(new_n783), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n847), .A2(new_n456), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n933), .A2(new_n316), .A3(new_n644), .A4(new_n911), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n932), .A2(KEYINPUT123), .A3(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT60), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n936), .A2(KEYINPUT122), .ZN(new_n938));
  NAND4_X1  g737(.A1(new_n932), .A2(KEYINPUT123), .A3(new_n934), .A4(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n932), .A2(new_n934), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(KEYINPUT122), .ZN(new_n941));
  AND3_X1   g740(.A1(new_n937), .A2(new_n939), .A3(new_n941), .ZN(G1350gat));
  NAND4_X1  g741(.A1(new_n914), .A2(new_n274), .A3(new_n621), .A4(new_n915), .ZN(new_n943));
  NAND4_X1  g742(.A1(new_n876), .A2(new_n853), .A3(new_n621), .A4(new_n918), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(G190gat), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT124), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n944), .A2(KEYINPUT124), .A3(G190gat), .ZN(new_n948));
  XOR2_X1   g747(.A(KEYINPUT125), .B(KEYINPUT61), .Z(new_n949));
  NAND3_X1  g748(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n947), .A2(new_n948), .ZN(new_n951));
  OR2_X1    g750(.A1(KEYINPUT125), .A2(KEYINPUT61), .ZN(new_n952));
  OAI211_X1 g751(.A(new_n943), .B(new_n950), .C1(new_n951), .C2(new_n952), .ZN(G1351gat));
  NAND2_X1  g752(.A1(new_n878), .A2(new_n879), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(KEYINPUT126), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT126), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n878), .A2(new_n879), .A3(new_n956), .ZN(new_n957));
  NOR3_X1   g756(.A1(new_n595), .A2(new_n456), .A3(new_n672), .ZN(new_n958));
  INV_X1    g757(.A(G197gat), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n271), .A2(new_n959), .ZN(new_n960));
  NAND4_X1  g759(.A1(new_n955), .A2(new_n957), .A3(new_n958), .A4(new_n960), .ZN(new_n961));
  NAND4_X1  g760(.A1(new_n876), .A2(new_n455), .A3(new_n374), .A4(new_n884), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n959), .B1(new_n962), .B2(new_n271), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n961), .A2(new_n963), .ZN(G1352gat));
  NAND4_X1  g763(.A1(new_n955), .A2(new_n667), .A3(new_n957), .A4(new_n958), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(G204gat), .ZN(new_n966));
  NOR3_X1   g765(.A1(new_n962), .A2(G204gat), .A3(new_n765), .ZN(new_n967));
  XNOR2_X1  g766(.A(new_n967), .B(KEYINPUT62), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n966), .A2(new_n968), .ZN(G1353gat));
  NAND2_X1  g768(.A1(new_n958), .A2(new_n644), .ZN(new_n970));
  OAI21_X1  g769(.A(G211gat), .B1(new_n954), .B2(new_n970), .ZN(new_n971));
  OR2_X1    g770(.A1(new_n971), .A2(KEYINPUT63), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(KEYINPUT63), .ZN(new_n973));
  OR2_X1    g772(.A1(new_n783), .A2(G211gat), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n962), .A2(new_n974), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT127), .ZN(new_n976));
  XNOR2_X1  g775(.A(new_n975), .B(new_n976), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n972), .A2(new_n973), .A3(new_n977), .ZN(G1354gat));
  INV_X1    g777(.A(G218gat), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n622), .A2(new_n979), .ZN(new_n980));
  NAND4_X1  g779(.A1(new_n955), .A2(new_n957), .A3(new_n958), .A4(new_n980), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n979), .B1(new_n962), .B2(new_n622), .ZN(new_n982));
  AND2_X1   g781(.A1(new_n981), .A2(new_n982), .ZN(G1355gat));
endmodule


