//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 0 1 1 1 0 1 1 1 0 0 1 0 0 1 0 1 0 0 1 0 0 1 0 0 0 1 0 1 1 0 1 0 0 0 1 1 1 0 0 0 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:33 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n450, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n564,
    new_n565, new_n566, new_n567, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n630,
    new_n631, new_n634, new_n636, new_n637, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT65), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT66), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT67), .ZN(G217));
  NOR4_X1   g026(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n454), .A2(G567), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT68), .Z(new_n458));
  AOI21_X1  g033(.A(new_n458), .B1(new_n453), .B2(G2106), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  AND2_X1   g035(.A1(new_n460), .A2(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G101), .ZN(new_n462));
  NAND2_X1  g037(.A1(KEYINPUT69), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g040(.A1(KEYINPUT69), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(new_n460), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n462), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  XNOR2_X1  g045(.A(KEYINPUT3), .B(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G125), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n460), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n470), .A2(new_n474), .ZN(G160));
  AOI21_X1  g050(.A(new_n460), .B1(new_n465), .B2(new_n466), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n460), .A2(G112), .ZN(new_n478));
  OAI21_X1  g053(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n468), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n480), .B1(G136), .B2(new_n481), .ZN(new_n482));
  XOR2_X1   g057(.A(new_n482), .B(KEYINPUT70), .Z(G162));
  AND3_X1   g058(.A1(KEYINPUT69), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n484));
  AOI21_X1  g059(.A(KEYINPUT3), .B1(KEYINPUT69), .B2(G2104), .ZN(new_n485));
  OAI211_X1 g060(.A(G126), .B(G2105), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(KEYINPUT71), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT71), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n467), .A2(new_n488), .A3(G126), .A4(G2105), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n491), .B1(new_n492), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  INV_X1    g071(.A(G138), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n471), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n460), .A2(G138), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n501), .B1(new_n465), .B2(new_n466), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n496), .B1(new_n502), .B2(KEYINPUT72), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n498), .B1(new_n484), .B2(new_n485), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT72), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n500), .B1(new_n503), .B2(new_n506), .ZN(new_n507));
  OAI21_X1  g082(.A(KEYINPUT73), .B1(new_n495), .B2(new_n507), .ZN(new_n508));
  OAI211_X1 g083(.A(KEYINPUT72), .B(new_n498), .C1(new_n484), .C2(new_n485), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(KEYINPUT4), .ZN(new_n510));
  AOI21_X1  g085(.A(KEYINPUT72), .B1(new_n467), .B2(new_n498), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n499), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n493), .B1(new_n487), .B2(new_n489), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT73), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n508), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(G164));
  AND2_X1   g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  NOR2_X1   g093(.A1(KEYINPUT5), .A2(G543), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AND2_X1   g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n524), .A2(G88), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n518), .A2(new_n519), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n526), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n527));
  INV_X1    g102(.A(G651), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  OAI21_X1  g104(.A(G543), .B1(new_n521), .B2(new_n522), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  AOI211_X1 g106(.A(new_n525), .B(new_n529), .C1(G50), .C2(new_n531), .ZN(G166));
  XNOR2_X1  g107(.A(KEYINPUT75), .B(KEYINPUT7), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT76), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n534), .B(new_n535), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n521), .A2(new_n522), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n537), .A2(G89), .ZN(new_n538));
  AND2_X1   g113(.A1(G63), .A2(G651), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n526), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n536), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n530), .A2(KEYINPUT74), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT74), .ZN(new_n543));
  OAI211_X1 g118(.A(new_n543), .B(G543), .C1(new_n521), .C2(new_n522), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  AND2_X1   g120(.A1(new_n545), .A2(G51), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n541), .A2(new_n546), .ZN(G168));
  AND2_X1   g122(.A1(new_n545), .A2(G52), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n526), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n526), .A2(new_n537), .ZN(new_n550));
  INV_X1    g125(.A(G90), .ZN(new_n551));
  OAI22_X1  g126(.A1(new_n549), .A2(new_n528), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n548), .A2(new_n552), .ZN(G171));
  NAND2_X1  g128(.A1(G68), .A2(G543), .ZN(new_n554));
  INV_X1    g129(.A(G56), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n520), .B2(new_n555), .ZN(new_n556));
  AOI22_X1  g131(.A1(G651), .A2(new_n556), .B1(new_n524), .B2(G81), .ZN(new_n557));
  INV_X1    g132(.A(new_n545), .ZN(new_n558));
  INV_X1    g133(.A(G43), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(G153));
  NAND4_X1  g137(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT77), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND4_X1  g141(.A1(G319), .A2(G483), .A3(G661), .A4(new_n566), .ZN(new_n567));
  XOR2_X1   g142(.A(new_n567), .B(KEYINPUT78), .Z(G188));
  INV_X1    g143(.A(KEYINPUT80), .ZN(new_n569));
  INV_X1    g144(.A(G53), .ZN(new_n570));
  OR4_X1    g145(.A1(new_n569), .A2(new_n530), .A3(KEYINPUT9), .A4(new_n570), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n537), .A2(G53), .A3(G543), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n569), .B1(new_n572), .B2(KEYINPUT9), .ZN(new_n573));
  OAI21_X1  g148(.A(KEYINPUT9), .B1(new_n530), .B2(new_n570), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(KEYINPUT79), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT79), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n572), .A2(new_n576), .A3(KEYINPUT9), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n571), .A2(new_n573), .A3(new_n575), .A4(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT81), .ZN(new_n579));
  NAND2_X1  g154(.A1(G78), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G65), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n520), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(G651), .A2(new_n582), .B1(new_n524), .B2(G91), .ZN(new_n583));
  AND3_X1   g158(.A1(new_n578), .A2(new_n579), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n579), .B1(new_n578), .B2(new_n583), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n584), .A2(new_n585), .ZN(G299));
  INV_X1    g161(.A(G171), .ZN(G301));
  INV_X1    g162(.A(G168), .ZN(G286));
  XNOR2_X1  g163(.A(G166), .B(KEYINPUT82), .ZN(G303));
  NAND2_X1  g164(.A1(new_n524), .A2(G87), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n531), .A2(G49), .ZN(new_n591));
  OAI21_X1  g166(.A(G651), .B1(new_n526), .B2(G74), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(G288));
  NAND2_X1  g168(.A1(G73), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G61), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n520), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n594), .B1(new_n596), .B2(KEYINPUT83), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n596), .A2(KEYINPUT83), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n528), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT84), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n599), .ZN(new_n603));
  OAI211_X1 g178(.A(new_n601), .B(G651), .C1(new_n603), .C2(new_n597), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n524), .A2(G86), .B1(new_n531), .B2(G48), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(G305));
  AND2_X1   g183(.A1(new_n545), .A2(G47), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n526), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G85), .ZN(new_n611));
  OAI22_X1  g186(.A1(new_n610), .A2(new_n528), .B1(new_n550), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(G290));
  NAND2_X1  g189(.A1(G301), .A2(G868), .ZN(new_n615));
  AND3_X1   g190(.A1(new_n524), .A2(KEYINPUT10), .A3(G92), .ZN(new_n616));
  AOI21_X1  g191(.A(KEYINPUT10), .B1(new_n524), .B2(G92), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n526), .A2(G66), .ZN(new_n619));
  NAND2_X1  g194(.A1(G79), .A2(G543), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n528), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(G54), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n622), .B1(new_n542), .B2(new_n544), .ZN(new_n623));
  INV_X1    g198(.A(KEYINPUT85), .ZN(new_n624));
  OR3_X1    g199(.A1(new_n621), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n621), .B2(new_n623), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n618), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n615), .B1(new_n627), .B2(G868), .ZN(G321));
  XOR2_X1   g203(.A(G321), .B(KEYINPUT86), .Z(G284));
  INV_X1    g204(.A(G868), .ZN(new_n630));
  NAND2_X1  g205(.A1(G299), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(new_n630), .B2(G168), .ZN(G297));
  OAI21_X1  g207(.A(new_n631), .B1(new_n630), .B2(G168), .ZN(G280));
  XNOR2_X1  g208(.A(KEYINPUT87), .B(G559), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n627), .B1(G860), .B2(new_n634), .ZN(G148));
  NAND2_X1  g210(.A1(new_n560), .A2(new_n630), .ZN(new_n636));
  AND2_X1   g211(.A1(new_n627), .A2(new_n634), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n636), .B1(new_n637), .B2(new_n630), .ZN(G323));
  XNOR2_X1  g213(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g214(.A1(new_n471), .A2(new_n461), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT12), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT13), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2100), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n476), .A2(G123), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n460), .A2(G111), .ZN(new_n645));
  OAI21_X1  g220(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n646));
  INV_X1    g221(.A(G135), .ZN(new_n647));
  OAI221_X1 g222(.A(new_n644), .B1(new_n645), .B2(new_n646), .C1(new_n647), .C2(new_n468), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(G2096), .Z(new_n649));
  NAND2_X1  g224(.A1(new_n643), .A2(new_n649), .ZN(G156));
  XNOR2_X1  g225(.A(KEYINPUT15), .B(G2435), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT88), .B(G2438), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2427), .B(G2430), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n655), .A2(KEYINPUT14), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2451), .B(G2454), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT16), .ZN(new_n659));
  XOR2_X1   g234(.A(G1341), .B(G1348), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n657), .B(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2443), .B(G2446), .Z(new_n663));
  AND2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g239(.A(G14), .B1(new_n662), .B2(new_n663), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(G401));
  XNOR2_X1  g241(.A(G2072), .B(G2078), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT17), .Z(new_n668));
  XNOR2_X1  g243(.A(G2067), .B(G2678), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G2084), .B(G2090), .Z(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n673), .B1(new_n669), .B2(new_n667), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT89), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n672), .A2(new_n669), .A3(new_n667), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT18), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n673), .A2(new_n669), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n678), .B1(new_n668), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n676), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G2096), .B(G2100), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(G227));
  XOR2_X1   g259(.A(G1971), .B(G1976), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT19), .ZN(new_n686));
  XOR2_X1   g261(.A(G1956), .B(G2474), .Z(new_n687));
  XOR2_X1   g262(.A(G1961), .B(G1966), .Z(new_n688));
  AND2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n687), .A2(new_n688), .ZN(new_n690));
  NOR3_X1   g265(.A1(new_n686), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n686), .A2(new_n689), .ZN(new_n692));
  XOR2_X1   g267(.A(KEYINPUT90), .B(KEYINPUT20), .Z(new_n693));
  XOR2_X1   g268(.A(new_n692), .B(new_n693), .Z(new_n694));
  AOI211_X1 g269(.A(new_n691), .B(new_n694), .C1(new_n686), .C2(new_n690), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1991), .B(G1996), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1981), .B(G1986), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(G229));
  NAND2_X1  g276(.A1(new_n607), .A2(G16), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(G6), .B2(G16), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT32), .B(G1981), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  AND2_X1   g280(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n703), .A2(new_n705), .ZN(new_n707));
  INV_X1    g282(.A(G16), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G22), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G166), .B2(new_n708), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(G1971), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n708), .A2(G23), .ZN(new_n712));
  INV_X1    g287(.A(G288), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n712), .B1(new_n713), .B2(new_n708), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT33), .B(G1976), .Z(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  NOR4_X1   g291(.A1(new_n706), .A2(new_n707), .A3(new_n711), .A4(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT34), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT92), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n613), .A2(new_n708), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(new_n708), .B2(G24), .ZN(new_n722));
  INV_X1    g297(.A(G1986), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n481), .A2(G131), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n476), .A2(G119), .ZN(new_n726));
  OAI21_X1  g301(.A(KEYINPUT91), .B1(G95), .B2(G2105), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  NOR3_X1   g303(.A1(KEYINPUT91), .A2(G95), .A3(G2105), .ZN(new_n729));
  OAI221_X1 g304(.A(G2104), .B1(G107), .B2(new_n460), .C1(new_n728), .C2(new_n729), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n725), .A2(new_n726), .A3(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G29), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G25), .B2(G29), .ZN(new_n734));
  XOR2_X1   g309(.A(KEYINPUT35), .B(G1991), .Z(new_n735));
  NAND2_X1  g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n724), .A2(new_n736), .ZN(new_n737));
  OAI22_X1  g312(.A1(new_n722), .A2(new_n723), .B1(new_n734), .B2(new_n735), .ZN(new_n738));
  AOI211_X1 g313(.A(new_n737), .B(new_n738), .C1(new_n717), .C2(new_n718), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n720), .A2(new_n739), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT93), .B(KEYINPUT36), .Z(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  AOI22_X1  g317(.A1(new_n471), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n743));
  OR3_X1    g318(.A1(new_n743), .A2(KEYINPUT96), .A3(new_n460), .ZN(new_n744));
  OAI21_X1  g319(.A(KEYINPUT96), .B1(new_n743), .B2(new_n460), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n481), .A2(G139), .ZN(new_n746));
  XOR2_X1   g321(.A(KEYINPUT95), .B(KEYINPUT25), .Z(new_n747));
  NAND3_X1  g322(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NAND4_X1  g324(.A1(new_n744), .A2(new_n745), .A3(new_n746), .A4(new_n749), .ZN(new_n750));
  MUX2_X1   g325(.A(G33), .B(new_n750), .S(G29), .Z(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT97), .Z(new_n752));
  INV_X1    g327(.A(G2072), .ZN(new_n753));
  OR2_X1    g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n752), .A2(new_n753), .ZN(new_n755));
  INV_X1    g330(.A(G29), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT24), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n756), .B1(new_n757), .B2(G34), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n757), .B2(G34), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G160), .B2(G29), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n756), .A2(G32), .ZN(new_n761));
  NAND3_X1  g336(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT26), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n762), .A2(new_n763), .ZN(new_n765));
  AOI22_X1  g340(.A1(new_n764), .A2(new_n765), .B1(G105), .B2(new_n461), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n476), .A2(G129), .ZN(new_n767));
  INV_X1    g342(.A(G141), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n766), .B(new_n767), .C1(new_n768), .C2(new_n468), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n761), .B1(new_n769), .B2(G29), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT27), .B(G1996), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n760), .A2(G2084), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n754), .A2(new_n755), .A3(new_n772), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT98), .Z(new_n774));
  NAND2_X1  g349(.A1(new_n708), .A2(G19), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(new_n561), .B2(new_n708), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(G1341), .Z(new_n777));
  NOR2_X1   g352(.A1(G4), .A2(G16), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n627), .B2(G16), .ZN(new_n779));
  OR2_X1    g354(.A1(new_n779), .A2(G1348), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n779), .A2(G1348), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n756), .A2(G26), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT28), .Z(new_n783));
  NAND2_X1  g358(.A1(new_n481), .A2(G140), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n476), .A2(G128), .ZN(new_n785));
  OR2_X1    g360(.A1(G104), .A2(G2105), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n786), .B(G2104), .C1(G116), .C2(new_n460), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n784), .A2(new_n785), .A3(new_n787), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n783), .B1(new_n788), .B2(G29), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G2067), .ZN(new_n790));
  NAND4_X1  g365(.A1(new_n777), .A2(new_n780), .A3(new_n781), .A4(new_n790), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT94), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n756), .A2(G35), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G162), .B2(new_n756), .ZN(new_n794));
  XOR2_X1   g369(.A(KEYINPUT99), .B(KEYINPUT29), .Z(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n796), .A2(G2090), .ZN(new_n797));
  INV_X1    g372(.A(G2078), .ZN(new_n798));
  NAND2_X1  g373(.A1(G164), .A2(G29), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G27), .B2(G29), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n797), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(new_n798), .B2(new_n800), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n708), .A2(G20), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT23), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n578), .A2(new_n583), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n805), .A2(KEYINPUT81), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n578), .A2(new_n579), .A3(new_n583), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n804), .B1(new_n808), .B2(new_n708), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(G1956), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n796), .A2(G2090), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n708), .A2(G21), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G168), .B2(new_n708), .ZN(new_n813));
  INV_X1    g388(.A(G1966), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(KEYINPUT30), .B(G28), .ZN(new_n816));
  OR2_X1    g391(.A1(KEYINPUT31), .A2(G11), .ZN(new_n817));
  NAND2_X1  g392(.A1(KEYINPUT31), .A2(G11), .ZN(new_n818));
  AOI22_X1  g393(.A1(new_n816), .A2(new_n756), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(new_n648), .B2(new_n756), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n708), .A2(G5), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(G171), .B2(new_n708), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n820), .B1(new_n822), .B2(G1961), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n822), .A2(G1961), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n760), .A2(G2084), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n770), .A2(new_n771), .ZN(new_n826));
  NOR3_X1   g401(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NAND4_X1  g402(.A1(new_n811), .A2(new_n815), .A3(new_n823), .A4(new_n827), .ZN(new_n828));
  NOR3_X1   g403(.A1(new_n802), .A2(new_n810), .A3(new_n828), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n742), .A2(new_n774), .A3(new_n792), .A4(new_n829), .ZN(G150));
  INV_X1    g405(.A(G150), .ZN(G311));
  NAND2_X1  g406(.A1(G80), .A2(G543), .ZN(new_n832));
  INV_X1    g407(.A(G67), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n832), .B1(new_n520), .B2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT100), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n835), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n836), .A2(G651), .A3(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  AND2_X1   g414(.A1(new_n545), .A2(G55), .ZN(new_n840));
  AND2_X1   g415(.A1(new_n524), .A2(G93), .ZN(new_n841));
  OAI21_X1  g416(.A(KEYINPUT101), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AOI22_X1  g417(.A1(new_n545), .A2(G55), .B1(G93), .B2(new_n524), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT101), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n839), .B1(new_n842), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n560), .B1(new_n846), .B2(KEYINPUT102), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(KEYINPUT102), .B2(new_n846), .ZN(new_n848));
  OR3_X1    g423(.A1(new_n846), .A2(KEYINPUT102), .A3(new_n561), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(KEYINPUT38), .Z(new_n851));
  NAND2_X1  g426(.A1(new_n627), .A2(G559), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n851), .B(new_n852), .Z(new_n853));
  INV_X1    g428(.A(KEYINPUT39), .ZN(new_n854));
  AOI21_X1  g429(.A(G860), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n855), .B1(new_n854), .B2(new_n853), .ZN(new_n856));
  INV_X1    g431(.A(new_n846), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(G860), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(KEYINPUT37), .Z(new_n859));
  NAND2_X1  g434(.A1(new_n856), .A2(new_n859), .ZN(G145));
  XNOR2_X1  g435(.A(new_n750), .B(new_n769), .ZN(new_n861));
  AOI22_X1  g436(.A1(new_n481), .A2(G142), .B1(G130), .B2(new_n476), .ZN(new_n862));
  OAI21_X1  g437(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT103), .ZN(new_n864));
  INV_X1    g439(.A(G118), .ZN(new_n865));
  AOI22_X1  g440(.A1(new_n863), .A2(new_n864), .B1(new_n865), .B2(G2105), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n866), .B1(new_n864), .B2(new_n863), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n862), .A2(new_n867), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n868), .B(new_n641), .Z(new_n869));
  XNOR2_X1  g444(.A(new_n861), .B(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n512), .A2(new_n513), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(new_n788), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(new_n732), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n870), .B(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(G160), .B(new_n648), .ZN(new_n875));
  XNOR2_X1  g450(.A(G162), .B(new_n875), .ZN(new_n876));
  AND2_X1   g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n874), .A2(new_n876), .ZN(new_n878));
  NOR3_X1   g453(.A1(new_n877), .A2(new_n878), .A3(G37), .ZN(new_n879));
  XOR2_X1   g454(.A(new_n879), .B(KEYINPUT40), .Z(G395));
  NAND2_X1  g455(.A1(new_n857), .A2(new_n630), .ZN(new_n881));
  INV_X1    g456(.A(new_n627), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n808), .A2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT104), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n884), .B1(G299), .B2(new_n627), .ZN(new_n885));
  AND4_X1   g460(.A1(new_n884), .A2(new_n806), .A3(new_n627), .A4(new_n807), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n883), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT41), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT105), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n890), .B1(new_n885), .B2(new_n886), .ZN(new_n891));
  OAI21_X1  g466(.A(KEYINPUT104), .B1(new_n808), .B2(new_n882), .ZN(new_n892));
  NAND3_X1  g467(.A1(G299), .A2(new_n884), .A3(new_n627), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n892), .A2(new_n893), .A3(KEYINPUT105), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n891), .A2(new_n883), .A3(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n889), .B1(new_n895), .B2(new_n888), .ZN(new_n896));
  XOR2_X1   g471(.A(new_n850), .B(new_n637), .Z(new_n897));
  MUX2_X1   g472(.A(new_n896), .B(new_n895), .S(new_n897), .Z(new_n898));
  XNOR2_X1  g473(.A(new_n607), .B(G290), .ZN(new_n899));
  XNOR2_X1  g474(.A(G166), .B(new_n713), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n899), .B(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(KEYINPUT106), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(KEYINPUT42), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n898), .B(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n881), .B1(new_n904), .B2(new_n630), .ZN(G295));
  OAI21_X1  g480(.A(new_n881), .B1(new_n904), .B2(new_n630), .ZN(G331));
  NAND2_X1  g481(.A1(G168), .A2(G171), .ZN(new_n907));
  OAI21_X1  g482(.A(G301), .B1(new_n541), .B2(new_n546), .ZN(new_n908));
  AND2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n850), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n909), .A2(new_n848), .A3(new_n849), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n896), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n895), .ZN(new_n915));
  OAI21_X1  g490(.A(KEYINPUT107), .B1(new_n915), .B2(new_n913), .ZN(new_n916));
  INV_X1    g491(.A(new_n901), .ZN(new_n917));
  AND3_X1   g492(.A1(new_n909), .A2(new_n848), .A3(new_n849), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n909), .B1(new_n849), .B2(new_n848), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT107), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n920), .A2(new_n921), .A3(new_n895), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n914), .A2(new_n916), .A3(new_n917), .A4(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(G37), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n915), .B1(new_n920), .B2(new_n888), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n913), .A2(KEYINPUT41), .A3(new_n887), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n925), .A2(new_n901), .A3(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n923), .A2(new_n924), .A3(new_n927), .ZN(new_n928));
  OR2_X1    g503(.A1(new_n928), .A2(KEYINPUT43), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n914), .A2(new_n916), .A3(new_n922), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(new_n901), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n923), .A2(new_n924), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT43), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n929), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT110), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n928), .A2(KEYINPUT109), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT109), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n923), .A2(new_n927), .A3(new_n940), .A4(new_n924), .ZN(new_n941));
  AND4_X1   g516(.A1(new_n938), .A2(new_n939), .A3(KEYINPUT43), .A4(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT43), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n943), .B1(new_n928), .B2(KEYINPUT109), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n938), .B1(new_n944), .B2(new_n941), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n933), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n947), .A2(new_n943), .A3(new_n931), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(KEYINPUT108), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT108), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n947), .A2(new_n950), .A3(new_n943), .A4(new_n931), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n949), .A2(KEYINPUT44), .A3(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n937), .B1(new_n946), .B2(new_n952), .ZN(G397));
  XNOR2_X1  g528(.A(KEYINPUT111), .B(G1384), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n954), .B1(new_n512), .B2(new_n513), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n955), .A2(KEYINPUT45), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(G160), .A2(G40), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(G2067), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n788), .B(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n959), .B1(new_n769), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(G1996), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n959), .A2(new_n964), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n965), .A2(KEYINPUT46), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n965), .A2(KEYINPUT46), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n963), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  XOR2_X1   g543(.A(new_n968), .B(KEYINPUT47), .Z(new_n969));
  XNOR2_X1  g544(.A(new_n769), .B(new_n964), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n961), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n735), .ZN(new_n972));
  OAI22_X1  g547(.A1(new_n971), .A2(new_n972), .B1(G2067), .B2(new_n788), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n959), .ZN(new_n974));
  XOR2_X1   g549(.A(new_n974), .B(KEYINPUT126), .Z(new_n975));
  NOR2_X1   g550(.A1(G290), .A2(G1986), .ZN(new_n976));
  AOI21_X1  g551(.A(KEYINPUT48), .B1(new_n959), .B2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n959), .A2(KEYINPUT48), .A3(new_n976), .ZN(new_n978));
  INV_X1    g553(.A(new_n959), .ZN(new_n979));
  XOR2_X1   g554(.A(new_n731), .B(new_n735), .Z(new_n980));
  NOR2_X1   g555(.A1(new_n971), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n978), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n975), .B1(new_n977), .B2(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n969), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G1981), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n607), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(G1981), .B1(new_n602), .B2(new_n606), .ZN(new_n987));
  AND3_X1   g562(.A1(new_n986), .A2(KEYINPUT49), .A3(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT49), .B1(new_n986), .B2(new_n987), .ZN(new_n989));
  INV_X1    g564(.A(G1384), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n871), .A2(new_n990), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n991), .A2(new_n958), .ZN(new_n992));
  INV_X1    g567(.A(G8), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  OR3_X1    g570(.A1(new_n988), .A2(new_n989), .A3(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G1976), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n996), .A2(new_n997), .A3(new_n713), .ZN(new_n998));
  AND2_X1   g573(.A1(new_n998), .A2(new_n986), .ZN(new_n999));
  NAND2_X1  g574(.A1(G303), .A2(G8), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n1000), .B(KEYINPUT55), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(G1384), .B1(new_n512), .B2(new_n513), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT50), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n958), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(G1384), .B1(new_n508), .B2(new_n515), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1005), .B1(new_n1006), .B2(new_n1004), .ZN(new_n1007));
  OR2_X1    g582(.A1(new_n1007), .A2(G2090), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n958), .B1(new_n955), .B2(KEYINPUT45), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1009), .B1(new_n1006), .B2(KEYINPUT45), .ZN(new_n1010));
  XOR2_X1   g585(.A(KEYINPUT112), .B(G1971), .Z(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n993), .B1(new_n1008), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1002), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n713), .A2(G1976), .ZN(new_n1015));
  AOI21_X1  g590(.A(KEYINPUT52), .B1(G288), .B2(new_n997), .ZN(new_n1016));
  AND3_X1   g591(.A1(new_n994), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n994), .A2(new_n1015), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1017), .B1(KEYINPUT52), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n996), .A2(new_n1019), .ZN(new_n1020));
  OAI22_X1  g595(.A1(new_n999), .A2(new_n995), .B1(new_n1014), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT114), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1019), .ZN(new_n1023));
  NOR3_X1   g598(.A1(new_n988), .A2(new_n989), .A3(new_n995), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1022), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n996), .A2(KEYINPUT114), .A3(new_n1019), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  AND2_X1   g602(.A1(G160), .A2(G40), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1028), .B1(KEYINPUT45), .B2(new_n1003), .ZN(new_n1029));
  AOI22_X1  g604(.A1(KEYINPUT45), .A2(new_n1006), .B1(new_n1029), .B2(KEYINPUT115), .ZN(new_n1030));
  OR2_X1    g605(.A1(new_n1029), .A2(KEYINPUT115), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n814), .ZN(new_n1033));
  OR2_X1    g608(.A1(new_n1007), .A2(G2084), .ZN(new_n1034));
  AND2_X1   g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NOR3_X1   g610(.A1(new_n1035), .A2(new_n993), .A3(G286), .ZN(new_n1036));
  AND3_X1   g611(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n514), .B1(new_n512), .B2(new_n513), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1004), .B(new_n990), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(KEYINPUT113), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT113), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n516), .A2(new_n1041), .A3(new_n1004), .A4(new_n990), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1028), .B1(new_n1004), .B2(new_n1003), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1040), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1012), .B1(new_n1045), .B2(G2090), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(G8), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1001), .A2(new_n1047), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1027), .A2(new_n1036), .A3(new_n1048), .A4(new_n1014), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT63), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1001), .A2(KEYINPUT116), .ZN(new_n1052));
  OR2_X1    g627(.A1(new_n1052), .A2(new_n1013), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1020), .A2(new_n1050), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1052), .A2(new_n1013), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1053), .A2(new_n1036), .A3(new_n1054), .A4(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1021), .B1(new_n1051), .B2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1030), .A2(new_n798), .A3(new_n1031), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT124), .ZN(new_n1059));
  OR2_X1    g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1060), .A2(KEYINPUT53), .A3(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1028), .B1(new_n991), .B2(KEYINPUT50), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n990), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1063), .B1(KEYINPUT50), .B2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1065), .A2(G1961), .ZN(new_n1066));
  OR2_X1    g641(.A1(new_n1010), .A2(G2078), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT53), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1066), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(G301), .B1(new_n1062), .B2(new_n1069), .ZN(new_n1070));
  AND4_X1   g645(.A1(new_n1070), .A2(new_n1027), .A3(new_n1048), .A4(new_n1014), .ZN(new_n1071));
  OR2_X1    g646(.A1(new_n1035), .A2(new_n993), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1072), .A2(G168), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1033), .A2(G168), .A3(new_n1034), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1074), .B(G8), .C1(KEYINPUT123), .C2(KEYINPUT51), .ZN(new_n1075));
  NAND2_X1  g650(.A1(KEYINPUT123), .A2(KEYINPUT51), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1074), .A2(G8), .ZN(new_n1078));
  NOR2_X1   g653(.A1(KEYINPUT123), .A2(KEYINPUT51), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1077), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1073), .B1(new_n1075), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT62), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1071), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1080), .A2(new_n1075), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1084), .B1(G168), .B2(new_n1072), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1085), .A2(KEYINPUT62), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1057), .B1(new_n1083), .B2(new_n1086), .ZN(new_n1087));
  AND3_X1   g662(.A1(new_n1027), .A2(new_n1048), .A3(new_n1014), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT54), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n957), .A2(KEYINPUT53), .A3(new_n1009), .A4(new_n798), .ZN(new_n1090));
  XOR2_X1   g665(.A(new_n1090), .B(KEYINPUT125), .Z(new_n1091));
  NAND2_X1  g666(.A1(new_n1069), .A2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1092), .A2(G171), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1089), .B1(new_n1070), .B2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1062), .A2(G301), .A3(new_n1069), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1089), .B1(new_n1092), .B2(G171), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1085), .A2(new_n1088), .A3(new_n1094), .A4(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT60), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT118), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1064), .A2(KEYINPUT50), .ZN(new_n1101));
  AOI21_X1  g676(.A(G1348), .B1(new_n1101), .B2(new_n1005), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n992), .A2(new_n960), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1100), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  OAI211_X1 g680(.A(KEYINPUT118), .B(new_n1103), .C1(new_n1065), .C2(G1348), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1099), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(KEYINPUT121), .ZN(new_n1108));
  NOR3_X1   g683(.A1(new_n1102), .A2(new_n1100), .A3(new_n1104), .ZN(new_n1109));
  INV_X1    g684(.A(G1348), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1007), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT118), .B1(new_n1111), .B2(new_n1103), .ZN(new_n1112));
  OAI21_X1  g687(.A(KEYINPUT60), .B1(new_n1109), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT121), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n882), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NOR3_X1   g690(.A1(new_n1107), .A2(KEYINPUT121), .A3(new_n627), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1108), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1105), .A2(new_n1099), .A3(new_n1106), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(G1956), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1045), .A2(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g696(.A(KEYINPUT117), .B(KEYINPUT57), .ZN(new_n1122));
  XNOR2_X1  g697(.A(new_n805), .B(new_n1122), .ZN(new_n1123));
  XNOR2_X1  g698(.A(KEYINPUT56), .B(G2072), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1009), .B(new_n1124), .C1(new_n1006), .C2(KEYINPUT45), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1121), .A2(new_n1123), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1123), .B1(new_n1121), .B2(new_n1125), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT119), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1126), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1121), .A2(KEYINPUT119), .A3(new_n1123), .A4(new_n1125), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1129), .A2(KEYINPUT61), .A3(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1123), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1043), .B1(new_n1039), .B2(KEYINPUT113), .ZN(new_n1133));
  AOI21_X1  g708(.A(G1956), .B1(new_n1133), .B2(new_n1042), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1125), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1132), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(new_n1126), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT61), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n964), .B(new_n1009), .C1(new_n1006), .C2(KEYINPUT45), .ZN(new_n1139));
  INV_X1    g714(.A(new_n992), .ZN(new_n1140));
  XOR2_X1   g715(.A(KEYINPUT58), .B(G1341), .Z(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1139), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(new_n561), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(KEYINPUT59), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT59), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1143), .A2(new_n1146), .A3(new_n561), .ZN(new_n1147));
  AOI22_X1  g722(.A1(new_n1137), .A2(new_n1138), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1131), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(KEYINPUT120), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT120), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1131), .A2(new_n1151), .A3(new_n1148), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1119), .A2(new_n1150), .A3(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1136), .B1(new_n1154), .B2(new_n882), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(new_n1126), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1153), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1098), .B1(new_n1157), .B2(KEYINPUT122), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT122), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1153), .A2(new_n1159), .A3(new_n1156), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1087), .B1(new_n1158), .B2(new_n1160), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n613), .B(G1986), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n979), .B1(new_n1162), .B2(new_n981), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n984), .B1(new_n1161), .B2(new_n1163), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g739(.A(KEYINPUT127), .ZN(new_n1166));
  NAND2_X1  g740(.A1(new_n683), .A2(G319), .ZN(new_n1167));
  NOR4_X1   g741(.A1(G229), .A2(new_n879), .A3(G401), .A4(new_n1167), .ZN(new_n1168));
  AND3_X1   g742(.A1(new_n935), .A2(new_n1166), .A3(new_n1168), .ZN(new_n1169));
  AOI21_X1  g743(.A(new_n1166), .B1(new_n935), .B2(new_n1168), .ZN(new_n1170));
  NOR2_X1   g744(.A1(new_n1169), .A2(new_n1170), .ZN(G308));
  NAND2_X1  g745(.A1(new_n935), .A2(new_n1168), .ZN(G225));
endmodule


