//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 1 1 0 0 0 1 1 0 0 0 0 0 1 1 1 0 0 1 0 1 1 1 1 1 0 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 1 0 0 0 1 0 0 1 0 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:28 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n438, new_n449, new_n450, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n572, new_n573,
    new_n574, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n600, new_n601, new_n602, new_n603, new_n604, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n625, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n635, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n848, new_n849, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1228, new_n1229, new_n1230;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  OR2_X1    g011(.A1(new_n436), .A2(KEYINPUT66), .ZN(new_n437));
  NAND2_X1  g012(.A1(new_n436), .A2(KEYINPUT66), .ZN(new_n438));
  NAND2_X1  g013(.A1(new_n437), .A2(new_n438), .ZN(G220));
  INV_X1    g014(.A(G96), .ZN(G221));
  INV_X1    g015(.A(G69), .ZN(G235));
  XOR2_X1   g016(.A(KEYINPUT67), .B(G120), .Z(G236));
  INV_X1    g017(.A(G57), .ZN(G237));
  INV_X1    g018(.A(G108), .ZN(G238));
  NAND4_X1  g019(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g023(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n449));
  AND2_X1   g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n449), .B(new_n450), .ZN(G223));
  NAND2_X1  g026(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g027(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR3_X1   g028(.A1(G218), .A2(G221), .A3(G219), .ZN(new_n454));
  NAND3_X1  g029(.A1(new_n437), .A2(new_n454), .A3(new_n438), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT2), .ZN(new_n456));
  NOR4_X1   g031(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  AOI22_X1  g035(.A1(new_n456), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT69), .ZN(new_n462));
  XOR2_X1   g037(.A(new_n462), .B(KEYINPUT70), .Z(G319));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT72), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT72), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n465), .A2(new_n467), .A3(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  NAND4_X1  g046(.A1(new_n468), .A2(G137), .A3(new_n469), .A4(new_n471), .ZN(new_n472));
  AOI21_X1  g047(.A(G2105), .B1(new_n465), .B2(new_n467), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(KEYINPUT73), .A3(G101), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  AOI21_X1  g050(.A(KEYINPUT73), .B1(new_n473), .B2(G101), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n472), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n478));
  AND3_X1   g053(.A1(new_n471), .A2(new_n478), .A3(KEYINPUT71), .ZN(new_n479));
  AOI21_X1  g054(.A(KEYINPUT71), .B1(new_n471), .B2(new_n478), .ZN(new_n480));
  OAI21_X1  g055(.A(G125), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(G113), .A2(G2104), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n469), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n477), .A2(new_n483), .ZN(G160));
  NAND2_X1  g059(.A1(new_n468), .A2(new_n471), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n485), .A2(new_n469), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G124), .ZN(new_n489));
  OR2_X1    g064(.A1(G100), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G112), .C2(new_n469), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n487), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  NAND2_X1  g068(.A1(new_n471), .A2(new_n478), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT71), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n471), .A2(new_n478), .A3(KEYINPUT71), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G138), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n499), .A2(G2105), .ZN(new_n500));
  AOI21_X1  g075(.A(KEYINPUT4), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n468), .A2(G126), .A3(new_n471), .ZN(new_n502));
  NAND2_X1  g077(.A1(G114), .A2(G2104), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n469), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n505), .A2(new_n499), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n468), .A2(new_n471), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(G102), .A2(G2104), .ZN(new_n508));
  AOI21_X1  g083(.A(G2105), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NOR3_X1   g084(.A1(new_n501), .A2(new_n504), .A3(new_n509), .ZN(G164));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n515), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n514), .ZN(new_n519));
  NOR2_X1   g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  AND2_X1   g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  OAI22_X1  g097(.A1(new_n519), .A2(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G88), .ZN(new_n524));
  OAI21_X1  g099(.A(G543), .B1(new_n521), .B2(new_n522), .ZN(new_n525));
  INV_X1    g100(.A(G50), .ZN(new_n526));
  OAI22_X1  g101(.A1(new_n523), .A2(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n518), .A2(new_n527), .ZN(G166));
  NAND3_X1  g103(.A1(new_n515), .A2(G63), .A3(G651), .ZN(new_n529));
  OAI211_X1 g104(.A(G51), .B(G543), .C1(new_n521), .C2(new_n522), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT74), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n529), .A2(KEYINPUT74), .A3(new_n530), .ZN(new_n534));
  OR2_X1    g109(.A1(KEYINPUT6), .A2(G651), .ZN(new_n535));
  NAND2_X1  g110(.A1(KEYINPUT6), .A2(G651), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n535), .A2(new_n536), .B1(new_n513), .B2(new_n514), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(KEYINPUT7), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n538), .A2(KEYINPUT7), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n537), .A2(G89), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n533), .A2(new_n534), .A3(new_n541), .ZN(G286));
  INV_X1    g117(.A(G286), .ZN(G168));
  INV_X1    g118(.A(KEYINPUT75), .ZN(new_n544));
  INV_X1    g119(.A(G64), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n545), .B1(new_n513), .B2(new_n514), .ZN(new_n546));
  NAND2_X1  g121(.A1(G77), .A2(G543), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n544), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n519), .A2(new_n520), .ZN(new_n550));
  OAI211_X1 g125(.A(KEYINPUT75), .B(new_n547), .C1(new_n550), .C2(new_n545), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n549), .A2(new_n551), .A3(G651), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT76), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g129(.A1(new_n549), .A2(new_n551), .A3(KEYINPUT76), .A4(G651), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n512), .B1(new_n535), .B2(new_n536), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n537), .A2(G90), .B1(new_n556), .B2(G52), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n554), .A2(new_n555), .A3(new_n557), .ZN(G301));
  INV_X1    g133(.A(G301), .ZN(G171));
  AOI22_X1  g134(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n560), .A2(new_n517), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n537), .A2(G81), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n556), .A2(G43), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(KEYINPUT77), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n537), .A2(G81), .B1(new_n556), .B2(G43), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT77), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n561), .B1(new_n565), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G860), .ZN(G153));
  NAND4_X1  g145(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g146(.A1(G1), .A2(G3), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT8), .ZN(new_n573));
  NAND4_X1  g148(.A1(G319), .A2(G483), .A3(G661), .A4(new_n573), .ZN(new_n574));
  XOR2_X1   g149(.A(new_n574), .B(KEYINPUT78), .Z(G188));
  INV_X1    g150(.A(KEYINPUT80), .ZN(new_n576));
  NAND2_X1  g151(.A1(G78), .A2(G543), .ZN(new_n577));
  XNOR2_X1  g152(.A(KEYINPUT79), .B(G65), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n550), .B2(new_n578), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n579), .A2(G651), .B1(G91), .B2(new_n537), .ZN(new_n580));
  OAI211_X1 g155(.A(G53), .B(G543), .C1(new_n521), .C2(new_n522), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n581), .B(KEYINPUT9), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n576), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n580), .A2(new_n576), .A3(new_n582), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G299));
  INV_X1    g162(.A(G166), .ZN(G303));
  NAND2_X1  g163(.A1(new_n556), .A2(G49), .ZN(new_n589));
  OAI21_X1  g164(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(G87), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n523), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(KEYINPUT81), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n537), .A2(G87), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT81), .ZN(new_n596));
  NAND4_X1  g171(.A1(new_n595), .A2(new_n596), .A3(new_n590), .A4(new_n589), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(G288));
  AOI22_X1  g174(.A1(new_n537), .A2(G86), .B1(new_n556), .B2(G48), .ZN(new_n600));
  INV_X1    g175(.A(G61), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n601), .B1(new_n513), .B2(new_n514), .ZN(new_n602));
  AND2_X1   g177(.A1(G73), .A2(G543), .ZN(new_n603));
  OAI21_X1  g178(.A(G651), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n600), .A2(new_n604), .ZN(G305));
  AOI22_X1  g180(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n606), .A2(new_n517), .ZN(new_n607));
  INV_X1    g182(.A(G85), .ZN(new_n608));
  XOR2_X1   g183(.A(KEYINPUT82), .B(G47), .Z(new_n609));
  OAI22_X1  g184(.A1(new_n523), .A2(new_n608), .B1(new_n609), .B2(new_n525), .ZN(new_n610));
  OR3_X1    g185(.A1(new_n607), .A2(new_n610), .A3(KEYINPUT83), .ZN(new_n611));
  OAI21_X1  g186(.A(KEYINPUT83), .B1(new_n607), .B2(new_n610), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(G290));
  NAND2_X1  g188(.A1(G301), .A2(G868), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n556), .A2(G54), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n515), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(new_n517), .ZN(new_n617));
  INV_X1    g192(.A(G92), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n523), .A2(new_n618), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n619), .A2(KEYINPUT10), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(KEYINPUT10), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n617), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n614), .B1(G868), .B2(new_n622), .ZN(G284));
  XNOR2_X1  g198(.A(G284), .B(KEYINPUT84), .ZN(G321));
  NAND2_X1  g199(.A1(G286), .A2(G868), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(new_n586), .B2(G868), .ZN(G297));
  OAI21_X1  g201(.A(new_n625), .B1(new_n586), .B2(G868), .ZN(G280));
  INV_X1    g202(.A(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n622), .B1(new_n628), .B2(G860), .ZN(G148));
  NAND2_X1  g204(.A1(new_n620), .A2(new_n621), .ZN(new_n630));
  INV_X1    g205(.A(new_n617), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  OAI21_X1  g207(.A(G868), .B1(new_n632), .B2(G559), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(G868), .B2(new_n569), .ZN(G323));
  XOR2_X1   g209(.A(KEYINPUT85), .B(KEYINPUT11), .Z(new_n635));
  XNOR2_X1  g210(.A(G323), .B(new_n635), .ZN(G282));
  NAND2_X1  g211(.A1(new_n498), .A2(new_n473), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(KEYINPUT12), .ZN(new_n638));
  INV_X1    g213(.A(KEYINPUT12), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n498), .A2(new_n639), .A3(new_n473), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT13), .ZN(new_n642));
  INV_X1    g217(.A(G2100), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n486), .A2(G135), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n488), .A2(G123), .ZN(new_n647));
  OAI21_X1  g222(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n648), .A2(KEYINPUT87), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n648), .A2(KEYINPUT87), .ZN(new_n650));
  OR3_X1    g225(.A1(new_n469), .A2(KEYINPUT86), .A3(G111), .ZN(new_n651));
  OAI21_X1  g226(.A(KEYINPUT86), .B1(new_n469), .B2(G111), .ZN(new_n652));
  NAND4_X1  g227(.A1(new_n649), .A2(new_n650), .A3(new_n651), .A4(new_n652), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n646), .A2(new_n647), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(G2096), .Z(new_n655));
  NAND3_X1  g230(.A1(new_n644), .A2(new_n645), .A3(new_n655), .ZN(G156));
  XNOR2_X1  g231(.A(KEYINPUT15), .B(G2435), .ZN(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT88), .B(G2438), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2427), .B(G2430), .Z(new_n660));
  OR2_X1    g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n659), .A2(new_n660), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n661), .A2(KEYINPUT14), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2451), .B(G2454), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT16), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1341), .B(G1348), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n663), .B(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2443), .B(G2446), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  OAI21_X1  g246(.A(G14), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n672), .B1(new_n671), .B2(new_n669), .ZN(G401));
  XOR2_X1   g248(.A(G2072), .B(G2078), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT89), .ZN(new_n675));
  XOR2_X1   g250(.A(KEYINPUT90), .B(KEYINPUT18), .Z(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G2084), .B(G2090), .Z(new_n678));
  XNOR2_X1  g253(.A(G2067), .B(G2678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n675), .B1(new_n677), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n680), .A2(KEYINPUT17), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n678), .A2(new_n679), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n676), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n681), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G2096), .B(G2100), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(G227));
  XNOR2_X1  g262(.A(G1971), .B(G1976), .ZN(new_n688));
  INV_X1    g263(.A(KEYINPUT19), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(G1956), .B(G2474), .Z(new_n691));
  XOR2_X1   g266(.A(G1961), .B(G1966), .Z(new_n692));
  AND2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT20), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n691), .A2(new_n692), .ZN(new_n696));
  NOR3_X1   g271(.A1(new_n690), .A2(new_n693), .A3(new_n696), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(new_n690), .B2(new_n696), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(G1991), .B(G1996), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(G1981), .B(G1986), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(G229));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G6), .ZN(new_n708));
  INV_X1    g283(.A(G305), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n708), .B1(new_n709), .B2(new_n707), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT91), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT32), .B(G1981), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n711), .A2(new_n712), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n707), .A2(G22), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G166), .B2(new_n707), .ZN(new_n716));
  INV_X1    g291(.A(G1971), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n707), .A2(G23), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n591), .A2(new_n593), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n719), .B1(new_n720), .B2(new_n707), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT33), .B(G1976), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NAND4_X1  g298(.A1(new_n713), .A2(new_n714), .A3(new_n718), .A4(new_n723), .ZN(new_n724));
  AND2_X1   g299(.A1(new_n724), .A2(KEYINPUT34), .ZN(new_n725));
  MUX2_X1   g300(.A(G24), .B(G290), .S(G16), .Z(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(G1986), .ZN(new_n727));
  INV_X1    g302(.A(G29), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G25), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n486), .A2(G131), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n488), .A2(G119), .ZN(new_n731));
  OR2_X1    g306(.A1(G95), .A2(G2105), .ZN(new_n732));
  OAI211_X1 g307(.A(new_n732), .B(G2104), .C1(G107), .C2(new_n469), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n730), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n729), .B1(new_n735), .B2(new_n728), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT35), .B(G1991), .Z(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n736), .B(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n727), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(KEYINPUT34), .B2(new_n724), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT92), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n740), .B(KEYINPUT92), .C1(KEYINPUT34), .C2(new_n724), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n725), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT93), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n746), .A2(KEYINPUT36), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(KEYINPUT36), .ZN(new_n748));
  AND3_X1   g323(.A1(new_n745), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n745), .A2(new_n747), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n728), .A2(G32), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n468), .A2(new_n471), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n752), .A2(G141), .A3(new_n469), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n752), .A2(G129), .A3(G2105), .ZN(new_n754));
  NAND3_X1  g329(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT26), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n755), .A2(new_n756), .ZN(new_n758));
  AOI22_X1  g333(.A1(G105), .A2(new_n473), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n753), .A2(new_n754), .A3(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n751), .B1(new_n761), .B2(new_n728), .ZN(new_n762));
  XOR2_X1   g337(.A(KEYINPUT27), .B(G1996), .Z(new_n763));
  OR2_X1    g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(G2084), .ZN(new_n765));
  AND2_X1   g340(.A1(KEYINPUT24), .A2(G34), .ZN(new_n766));
  NOR2_X1   g341(.A1(KEYINPUT24), .A2(G34), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n728), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT96), .Z(new_n769));
  INV_X1    g344(.A(G160), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n769), .B1(new_n770), .B2(new_n728), .ZN(new_n771));
  NOR2_X1   g346(.A1(G168), .A2(new_n707), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(new_n707), .B2(G21), .ZN(new_n773));
  INV_X1    g348(.A(G1966), .ZN(new_n774));
  OAI221_X1 g349(.A(new_n764), .B1(new_n765), .B2(new_n771), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(G171), .A2(new_n707), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G5), .B2(new_n707), .ZN(new_n777));
  INV_X1    g352(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n775), .B1(G1961), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(G164), .A2(G29), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G27), .B2(G29), .ZN(new_n781));
  INV_X1    g356(.A(G2078), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  XOR2_X1   g358(.A(KEYINPUT31), .B(G11), .Z(new_n784));
  INV_X1    g359(.A(KEYINPUT30), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n728), .B1(new_n785), .B2(G28), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT98), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  AOI22_X1  g363(.A1(new_n786), .A2(new_n787), .B1(new_n785), .B2(G28), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n784), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(new_n654), .B2(new_n728), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n781), .A2(new_n782), .ZN(new_n792));
  AOI211_X1 g367(.A(new_n791), .B(new_n792), .C1(new_n774), .C2(new_n773), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n779), .A2(new_n783), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n728), .A2(G35), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT100), .Z(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G162), .B2(new_n728), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT29), .Z(new_n798));
  INV_X1    g373(.A(G2090), .ZN(new_n799));
  INV_X1    g374(.A(G2072), .ZN(new_n800));
  AND2_X1   g375(.A1(new_n728), .A2(G33), .ZN(new_n801));
  AND2_X1   g376(.A1(new_n498), .A2(G127), .ZN(new_n802));
  AND2_X1   g377(.A1(G115), .A2(G2104), .ZN(new_n803));
  OAI21_X1  g378(.A(G2105), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n752), .A2(G139), .A3(new_n469), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT25), .Z(new_n807));
  AND3_X1   g382(.A1(new_n805), .A2(KEYINPUT95), .A3(new_n807), .ZN(new_n808));
  AOI21_X1  g383(.A(KEYINPUT95), .B1(new_n805), .B2(new_n807), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n804), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n801), .B1(new_n810), .B2(G29), .ZN(new_n811));
  AOI22_X1  g386(.A1(new_n798), .A2(new_n799), .B1(new_n800), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n707), .A2(G20), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT23), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(new_n586), .B2(new_n707), .ZN(new_n815));
  INV_X1    g390(.A(G1956), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n812), .B(new_n817), .C1(new_n799), .C2(new_n798), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n794), .A2(new_n818), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n771), .A2(new_n765), .B1(new_n762), .B2(new_n763), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(new_n778), .B2(G1961), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT99), .Z(new_n822));
  NOR2_X1   g397(.A1(new_n811), .A2(new_n800), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT97), .Z(new_n824));
  NAND2_X1  g399(.A1(new_n707), .A2(G4), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(new_n622), .B2(new_n707), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(G1348), .Z(new_n827));
  NAND2_X1  g402(.A1(new_n569), .A2(G16), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(G16), .B2(G19), .ZN(new_n829));
  INV_X1    g404(.A(G1341), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n728), .A2(G26), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT28), .ZN(new_n833));
  NAND4_X1  g408(.A1(new_n468), .A2(G140), .A3(new_n469), .A4(new_n471), .ZN(new_n834));
  NAND4_X1  g409(.A1(new_n468), .A2(G128), .A3(G2105), .A4(new_n471), .ZN(new_n835));
  OR2_X1    g410(.A1(G104), .A2(G2105), .ZN(new_n836));
  OAI211_X1 g411(.A(new_n836), .B(G2104), .C1(G116), .C2(new_n469), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n834), .A2(new_n835), .A3(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n833), .B1(new_n839), .B2(new_n728), .ZN(new_n840));
  INV_X1    g415(.A(G2067), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n829), .A2(new_n830), .ZN(new_n843));
  NAND4_X1  g418(.A1(new_n827), .A2(new_n831), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT94), .ZN(new_n845));
  NAND4_X1  g420(.A1(new_n819), .A2(new_n822), .A3(new_n824), .A4(new_n845), .ZN(new_n846));
  NOR3_X1   g421(.A1(new_n749), .A2(new_n750), .A3(new_n846), .ZN(G311));
  NOR2_X1   g422(.A1(new_n750), .A2(new_n846), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n745), .A2(new_n747), .A3(new_n748), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(G150));
  AOI22_X1  g425(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n851), .A2(new_n517), .ZN(new_n852));
  INV_X1    g427(.A(G93), .ZN(new_n853));
  INV_X1    g428(.A(G55), .ZN(new_n854));
  OAI22_X1  g429(.A1(new_n523), .A2(new_n853), .B1(new_n525), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(G860), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(KEYINPUT37), .Z(new_n859));
  INV_X1    g434(.A(KEYINPUT39), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT101), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n569), .A2(new_n861), .ZN(new_n862));
  AOI211_X1 g437(.A(KEYINPUT101), .B(new_n561), .C1(new_n565), .C2(new_n568), .ZN(new_n863));
  NOR3_X1   g438(.A1(new_n862), .A2(new_n863), .A3(new_n857), .ZN(new_n864));
  INV_X1    g439(.A(new_n561), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n566), .A2(new_n567), .ZN(new_n866));
  AND3_X1   g441(.A1(new_n562), .A2(new_n567), .A3(new_n563), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n865), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(KEYINPUT101), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n569), .A2(new_n861), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n856), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(KEYINPUT38), .B1(new_n864), .B2(new_n871), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n632), .A2(new_n628), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n857), .B1(new_n862), .B2(new_n863), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT38), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n869), .A2(new_n870), .A3(new_n856), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  AND3_X1   g452(.A1(new_n872), .A2(new_n873), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n873), .B1(new_n872), .B2(new_n877), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n860), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT102), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n878), .A2(new_n879), .ZN(new_n882));
  AOI21_X1  g457(.A(G860), .B1(new_n882), .B2(KEYINPUT39), .ZN(new_n883));
  AND3_X1   g458(.A1(new_n881), .A2(KEYINPUT103), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(KEYINPUT103), .B1(new_n881), .B2(new_n883), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n859), .B1(new_n884), .B2(new_n885), .ZN(G145));
  INV_X1    g461(.A(KEYINPUT107), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n810), .A2(KEYINPUT105), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT105), .ZN(new_n889));
  OAI211_X1 g464(.A(new_n804), .B(new_n889), .C1(new_n808), .C2(new_n809), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n760), .A2(new_n839), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n838), .A2(new_n753), .A3(new_n754), .A4(new_n759), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n502), .A2(new_n503), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(G2105), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n507), .A2(new_n508), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(new_n469), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n500), .B1(new_n479), .B2(new_n480), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(new_n505), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n895), .A2(new_n897), .A3(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT104), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(G164), .A2(KEYINPUT104), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n893), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n893), .B1(new_n903), .B2(new_n902), .ZN(new_n906));
  OAI211_X1 g481(.A(new_n888), .B(new_n890), .C1(new_n905), .C2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n903), .A2(new_n902), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n908), .A2(new_n891), .A3(new_n892), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n909), .A2(KEYINPUT105), .A3(new_n810), .A4(new_n904), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n486), .A2(G142), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n488), .A2(G130), .ZN(new_n913));
  OR2_X1    g488(.A1(G106), .A2(G2105), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n914), .B(G2104), .C1(G118), .C2(new_n469), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n641), .A2(new_n912), .A3(new_n913), .A4(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n912), .A2(new_n913), .A3(new_n915), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n917), .A2(new_n638), .A3(new_n640), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n916), .A2(new_n918), .A3(new_n735), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n735), .B1(new_n916), .B2(new_n918), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(KEYINPUT106), .B1(new_n911), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT106), .ZN(new_n924));
  AOI211_X1 g499(.A(new_n924), .B(new_n921), .C1(new_n907), .C2(new_n910), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n887), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  NOR3_X1   g501(.A1(new_n905), .A2(new_n906), .A3(new_n888), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n888), .A2(new_n890), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n928), .B1(new_n909), .B2(new_n904), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n922), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(new_n924), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n911), .A2(KEYINPUT106), .A3(new_n922), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n931), .A2(KEYINPUT107), .A3(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n911), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(new_n921), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n926), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n492), .B(new_n654), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n937), .B(new_n770), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n931), .A2(new_n932), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n938), .B1(new_n934), .B2(new_n921), .ZN(new_n941));
  AOI21_X1  g516(.A(G37), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n939), .A2(KEYINPUT40), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(KEYINPUT40), .B1(new_n939), .B2(new_n942), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n943), .A2(new_n944), .ZN(G395));
  INV_X1    g520(.A(new_n585), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n632), .B1(new_n946), .B2(new_n583), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n584), .A2(new_n622), .A3(new_n585), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n632), .A2(G559), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n951), .B(KEYINPUT108), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n952), .B1(new_n864), .B2(new_n871), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT108), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n951), .B(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n955), .A2(new_n876), .A3(new_n874), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n950), .B1(new_n953), .B2(new_n956), .ZN(new_n957));
  OR2_X1    g532(.A1(new_n957), .A2(KEYINPUT109), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT42), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT113), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT112), .ZN(new_n961));
  NAND2_X1  g536(.A1(G303), .A2(new_n961), .ZN(new_n962));
  NOR3_X1   g537(.A1(new_n518), .A2(new_n527), .A3(new_n961), .ZN(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(G290), .A2(new_n962), .A3(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(G166), .A2(KEYINPUT112), .ZN(new_n966));
  OAI211_X1 g541(.A(new_n612), .B(new_n611), .C1(new_n966), .C2(new_n963), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n709), .B(new_n720), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n965), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n968), .B1(new_n965), .B2(new_n967), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n960), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n965), .A2(new_n967), .ZN(new_n973));
  INV_X1    g548(.A(new_n968), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n975), .A2(KEYINPUT113), .A3(new_n969), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n959), .B1(new_n972), .B2(new_n976), .ZN(new_n977));
  NOR3_X1   g552(.A1(new_n970), .A2(new_n971), .A3(KEYINPUT42), .ZN(new_n978));
  OR3_X1    g553(.A1(new_n977), .A2(KEYINPUT114), .A3(new_n978), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n953), .A2(new_n956), .ZN(new_n980));
  XOR2_X1   g555(.A(KEYINPUT111), .B(KEYINPUT41), .Z(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n950), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n947), .A2(new_n948), .A3(KEYINPUT110), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT41), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT110), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n586), .A2(new_n986), .A3(new_n632), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n984), .A2(new_n985), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n983), .A2(new_n988), .ZN(new_n989));
  AOI22_X1  g564(.A1(KEYINPUT109), .A2(new_n957), .B1(new_n980), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(KEYINPUT114), .B1(new_n977), .B2(new_n978), .ZN(new_n991));
  AND4_X1   g566(.A1(new_n958), .A2(new_n979), .A3(new_n990), .A4(new_n991), .ZN(new_n992));
  AOI22_X1  g567(.A1(new_n991), .A2(new_n979), .B1(new_n990), .B2(new_n958), .ZN(new_n993));
  OAI21_X1  g568(.A(G868), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n994), .B1(G868), .B2(new_n856), .ZN(G295));
  OAI21_X1  g570(.A(new_n994), .B1(G868), .B2(new_n856), .ZN(G331));
  NAND2_X1  g571(.A1(new_n972), .A2(new_n976), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT115), .ZN(new_n999));
  NAND2_X1  g574(.A1(G286), .A2(new_n999), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n533), .A2(KEYINPUT115), .A3(new_n541), .A4(new_n534), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(G171), .ZN(new_n1003));
  NAND3_X1  g578(.A1(G301), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1005), .B1(new_n864), .B2(new_n871), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n874), .A2(new_n876), .A3(new_n1004), .A4(new_n1003), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n950), .B1(new_n1008), .B2(new_n982), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n984), .A2(new_n987), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(KEYINPUT41), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1011), .B1(new_n1007), .B2(new_n1006), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n998), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT43), .ZN(new_n1014));
  INV_X1    g589(.A(G37), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1008), .A2(new_n989), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1006), .A2(new_n1007), .A3(new_n949), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1016), .A2(new_n997), .A3(new_n1017), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .A4(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT116), .ZN(new_n1020));
  AND2_X1   g595(.A1(new_n1018), .A2(new_n1015), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT116), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1021), .A2(new_n1022), .A3(new_n1014), .A4(new_n1013), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1018), .A2(new_n1015), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n997), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1025));
  OAI21_X1  g600(.A(KEYINPUT43), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1020), .A2(new_n1023), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT44), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1021), .A2(KEYINPUT43), .A3(new_n1013), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1014), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(KEYINPUT44), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1029), .A2(new_n1033), .ZN(G397));
  INV_X1    g609(.A(KEYINPUT45), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1035), .B1(G164), .B2(G1384), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n481), .A2(new_n482), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(G2105), .ZN(new_n1038));
  INV_X1    g613(.A(new_n476), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(new_n474), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1038), .A2(G40), .A3(new_n472), .A4(new_n1040), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1036), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1042), .A2(G1996), .A3(new_n760), .ZN(new_n1043));
  XOR2_X1   g618(.A(new_n1043), .B(KEYINPUT117), .Z(new_n1044));
  NOR2_X1   g619(.A1(new_n735), .A2(new_n737), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n734), .A2(new_n738), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1042), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g622(.A(new_n838), .B(new_n841), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1048), .B1(G1996), .B2(new_n760), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1042), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1044), .A2(new_n1047), .A3(new_n1050), .ZN(new_n1051));
  XNOR2_X1  g626(.A(G290), .B(G1986), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1051), .B1(new_n1042), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(G40), .ZN(new_n1054));
  NOR3_X1   g629(.A1(new_n477), .A2(new_n483), .A3(new_n1054), .ZN(new_n1055));
  AOI22_X1  g630(.A1(new_n469), .A2(new_n896), .B1(new_n898), .B2(new_n505), .ZN(new_n1056));
  AOI21_X1  g631(.A(G1384), .B1(new_n1056), .B2(new_n895), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT50), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1055), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G1384), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n900), .A2(new_n1058), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n816), .B1(new_n1059), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT121), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT57), .B1(new_n582), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT122), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n580), .A2(new_n1067), .A3(new_n582), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1067), .B1(new_n580), .B2(new_n582), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1066), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1070), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1072), .A2(new_n1065), .A3(new_n1068), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n900), .A2(KEYINPUT45), .A3(new_n1060), .ZN(new_n1075));
  XNOR2_X1  g650(.A(KEYINPUT56), .B(G2072), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1036), .A2(new_n1055), .A3(new_n1075), .A4(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1063), .A2(new_n1074), .A3(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n900), .A2(new_n1060), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1041), .B1(new_n1079), .B2(KEYINPUT50), .ZN(new_n1080));
  AOI21_X1  g655(.A(G1348), .B1(new_n1080), .B2(new_n1061), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1057), .A2(new_n1055), .A3(new_n841), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1084), .A2(new_n632), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1074), .B1(new_n1063), .B2(new_n1077), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1078), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT61), .ZN(new_n1088));
  AND3_X1   g663(.A1(new_n1063), .A2(new_n1074), .A3(new_n1077), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1088), .B1(new_n1089), .B2(new_n1086), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1074), .ZN(new_n1091));
  AOI21_X1  g666(.A(G1956), .B1(new_n1080), .B2(new_n1061), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1077), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1091), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1094), .A2(KEYINPUT61), .A3(new_n1078), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT60), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1059), .A2(new_n1062), .ZN(new_n1098));
  OAI211_X1 g673(.A(KEYINPUT60), .B(new_n1082), .C1(new_n1098), .C2(G1348), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1097), .A2(new_n1099), .A3(new_n622), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1084), .A2(KEYINPUT60), .A3(new_n632), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1090), .A2(new_n1095), .A3(new_n1100), .A4(new_n1101), .ZN(new_n1102));
  XNOR2_X1  g677(.A(KEYINPUT123), .B(G1996), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1036), .A2(new_n1055), .A3(new_n1075), .A4(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1057), .A2(new_n1055), .ZN(new_n1106));
  XOR2_X1   g681(.A(KEYINPUT58), .B(G1341), .Z(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n868), .B1(new_n1105), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT124), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT59), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1113), .B1(new_n1109), .B2(KEYINPUT124), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1110), .A2(new_n1111), .A3(new_n1113), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1087), .B1(new_n1102), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT51), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1055), .B1(new_n1057), .B2(KEYINPUT45), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1075), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n774), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1079), .A2(KEYINPUT50), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1123), .A2(new_n765), .A3(new_n1055), .A4(new_n1061), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1122), .A2(G168), .A3(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1119), .B1(new_n1125), .B2(G8), .ZN(new_n1126));
  AND2_X1   g701(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1127));
  OAI21_X1  g702(.A(KEYINPUT51), .B1(new_n1127), .B2(G168), .ZN(new_n1128));
  AND2_X1   g703(.A1(new_n1125), .A2(G8), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1126), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(G303), .A2(G8), .ZN(new_n1131));
  XNOR2_X1  g706(.A(new_n1131), .B(KEYINPUT55), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1036), .A2(new_n1055), .A3(new_n1075), .ZN(new_n1133));
  AOI22_X1  g708(.A1(new_n1098), .A2(new_n799), .B1(new_n717), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(G8), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1132), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1133), .A2(new_n717), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1080), .A2(new_n799), .A3(new_n1061), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1135), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1132), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n720), .A2(G1976), .ZN(new_n1142));
  OAI211_X1 g717(.A(G8), .B(new_n1142), .C1(new_n1079), .C2(new_n1041), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(KEYINPUT52), .ZN(new_n1144));
  INV_X1    g719(.A(G1981), .ZN(new_n1145));
  AND3_X1   g720(.A1(new_n600), .A2(new_n1145), .A3(new_n604), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1145), .B1(new_n600), .B2(new_n604), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT49), .ZN(new_n1148));
  OAI22_X1  g723(.A1(new_n1146), .A2(new_n1147), .B1(KEYINPUT118), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(KEYINPUT118), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  OAI211_X1 g726(.A(KEYINPUT118), .B(new_n1148), .C1(new_n1146), .C2(new_n1147), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1151), .A2(new_n1106), .A3(G8), .A4(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(G1976), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n594), .A2(new_n1154), .A3(new_n597), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT52), .ZN(new_n1156));
  AND2_X1   g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1157), .A2(new_n1106), .A3(G8), .A4(new_n1142), .ZN(new_n1158));
  AND3_X1   g733(.A1(new_n1144), .A2(new_n1153), .A3(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1136), .A2(new_n1141), .A3(new_n1159), .ZN(new_n1160));
  AND2_X1   g735(.A1(KEYINPUT125), .A2(G2078), .ZN(new_n1161));
  NOR2_X1   g736(.A1(KEYINPUT125), .A2(G2078), .ZN(new_n1162));
  OAI21_X1  g737(.A(KEYINPUT53), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  OR2_X1    g738(.A1(new_n1133), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT53), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1165), .B1(new_n1133), .B2(G2078), .ZN(new_n1166));
  INV_X1    g741(.A(G1961), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1167), .B1(new_n1059), .B2(new_n1062), .ZN(new_n1168));
  XOR2_X1   g743(.A(G301), .B(KEYINPUT54), .Z(new_n1169));
  NAND4_X1  g744(.A1(new_n1164), .A2(new_n1166), .A3(new_n1168), .A4(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1041), .B1(new_n1079), .B2(new_n1035), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n1171), .A2(KEYINPUT53), .A3(new_n782), .A4(new_n1075), .ZN(new_n1172));
  AND3_X1   g747(.A1(new_n1166), .A2(new_n1172), .A3(new_n1168), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1170), .B1(new_n1173), .B2(new_n1169), .ZN(new_n1174));
  NOR3_X1   g749(.A1(new_n1130), .A2(new_n1160), .A3(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1118), .A2(new_n1175), .ZN(new_n1176));
  AOI211_X1 g751(.A(new_n1135), .B(G286), .C1(new_n1122), .C2(new_n1124), .ZN(new_n1177));
  NAND4_X1  g752(.A1(new_n1136), .A2(new_n1141), .A3(new_n1159), .A4(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT120), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT63), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1178), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1153), .A2(new_n1154), .A3(new_n598), .ZN(new_n1182));
  INV_X1    g757(.A(new_n1146), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  OR2_X1    g759(.A1(new_n1184), .A2(KEYINPUT119), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1106), .A2(G8), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1186), .B1(new_n1184), .B2(KEYINPUT119), .ZN(new_n1187));
  AOI211_X1 g762(.A(new_n1135), .B(new_n1132), .C1(new_n1137), .C2(new_n1138), .ZN(new_n1188));
  AOI22_X1  g763(.A1(new_n1185), .A2(new_n1187), .B1(new_n1188), .B2(new_n1159), .ZN(new_n1189));
  AND2_X1   g764(.A1(new_n1181), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1176), .A2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1159), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1192));
  INV_X1    g767(.A(new_n1192), .ZN(new_n1193));
  NAND4_X1  g768(.A1(new_n1193), .A2(KEYINPUT63), .A3(new_n1141), .A4(new_n1177), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1178), .A2(new_n1180), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1194), .A2(new_n1195), .A3(KEYINPUT120), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1125), .A2(G8), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1197), .A2(KEYINPUT51), .ZN(new_n1198));
  AOI21_X1  g773(.A(G168), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1199));
  OAI211_X1 g774(.A(G8), .B(new_n1125), .C1(new_n1199), .C2(new_n1119), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT62), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1198), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1166), .A2(new_n1172), .A3(new_n1168), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1203), .A2(G171), .ZN(new_n1204));
  NOR3_X1   g779(.A1(new_n1192), .A2(new_n1204), .A3(new_n1188), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1201), .B1(new_n1198), .B2(new_n1200), .ZN(new_n1206));
  INV_X1    g781(.A(KEYINPUT126), .ZN(new_n1207));
  OAI211_X1 g782(.A(new_n1202), .B(new_n1205), .C1(new_n1206), .C2(new_n1207), .ZN(new_n1208));
  NOR3_X1   g783(.A1(new_n1130), .A2(KEYINPUT126), .A3(new_n1201), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n1196), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g785(.A(new_n1053), .B1(new_n1191), .B2(new_n1210), .ZN(new_n1211));
  OR3_X1    g786(.A1(new_n1036), .A2(G1996), .A3(new_n1041), .ZN(new_n1212));
  INV_X1    g787(.A(KEYINPUT46), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1048), .A2(new_n761), .ZN(new_n1214));
  AOI22_X1  g789(.A1(new_n1212), .A2(new_n1213), .B1(new_n1042), .B2(new_n1214), .ZN(new_n1215));
  OAI21_X1  g790(.A(new_n1215), .B1(new_n1213), .B2(new_n1212), .ZN(new_n1216));
  XNOR2_X1  g791(.A(KEYINPUT127), .B(KEYINPUT47), .ZN(new_n1217));
  XNOR2_X1  g792(.A(new_n1216), .B(new_n1217), .ZN(new_n1218));
  NOR2_X1   g793(.A1(G290), .A2(G1986), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n1042), .A2(new_n1219), .ZN(new_n1220));
  XOR2_X1   g795(.A(new_n1220), .B(KEYINPUT48), .Z(new_n1221));
  OAI21_X1  g796(.A(new_n1218), .B1(new_n1051), .B2(new_n1221), .ZN(new_n1222));
  NAND3_X1  g797(.A1(new_n1044), .A2(new_n1046), .A3(new_n1050), .ZN(new_n1223));
  OAI21_X1  g798(.A(new_n1223), .B1(G2067), .B2(new_n838), .ZN(new_n1224));
  AOI21_X1  g799(.A(new_n1222), .B1(new_n1042), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1211), .A2(new_n1225), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g801(.A1(G401), .A2(new_n462), .A3(G227), .ZN(new_n1228));
  NAND2_X1  g802(.A1(new_n705), .A2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g803(.A(new_n1229), .B1(new_n939), .B2(new_n942), .ZN(new_n1230));
  AND2_X1   g804(.A1(new_n1230), .A2(new_n1027), .ZN(G308));
  NAND2_X1  g805(.A1(new_n1230), .A2(new_n1027), .ZN(G225));
endmodule


