//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 0 0 0 0 0 0 1 0 0 1 1 0 1 1 0 1 0 0 0 0 1 1 1 1 0 0 0 1 1 1 1 1 0 0 1 0 1 1 0 1 0 1 1 1 1 0 0 0 1 0 1 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n759, new_n760, new_n761, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n775, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n869, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1013, new_n1014;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  NAND2_X1  g001(.A1(G225gat), .A2(G233gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  OR2_X1    g003(.A1(G113gat), .A2(G120gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT1), .ZN(new_n206));
  NAND2_X1  g005(.A1(G113gat), .A2(G120gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G127gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G134gat), .ZN(new_n210));
  INV_X1    g009(.A(G134gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G127gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT69), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n210), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n209), .A2(KEYINPUT69), .A3(G134gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n208), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G127gat), .B(G134gat), .ZN(new_n217));
  XNOR2_X1  g016(.A(KEYINPUT70), .B(KEYINPUT1), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n217), .A2(new_n218), .A3(new_n205), .A4(new_n207), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n216), .A2(new_n219), .ZN(new_n220));
  AND2_X1   g019(.A1(G155gat), .A2(G162gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(G155gat), .A2(G162gat), .ZN(new_n222));
  OAI21_X1  g021(.A(KEYINPUT77), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  AND2_X1   g022(.A1(G141gat), .A2(G148gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(G141gat), .A2(G148gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G155gat), .ZN(new_n227));
  INV_X1    g026(.A(G162gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT77), .ZN(new_n230));
  AOI21_X1  g029(.A(KEYINPUT2), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  OAI211_X1 g030(.A(new_n223), .B(new_n226), .C1(new_n231), .C2(new_n221), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT2), .ZN(new_n233));
  NOR3_X1   g032(.A1(new_n224), .A2(new_n225), .A3(KEYINPUT76), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT76), .ZN(new_n235));
  INV_X1    g034(.A(G141gat), .ZN(new_n236));
  INV_X1    g035(.A(G148gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(G141gat), .A2(G148gat), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n235), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n233), .B1(new_n234), .B2(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(G155gat), .B(G162gat), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n220), .B1(new_n232), .B2(new_n244), .ZN(new_n245));
  OAI21_X1  g044(.A(KEYINPUT76), .B1(new_n224), .B2(new_n225), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n238), .A2(new_n235), .A3(new_n239), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT2), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n232), .B1(new_n248), .B2(new_n242), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n216), .A2(new_n219), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n204), .B1(new_n245), .B2(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(KEYINPUT78), .B(KEYINPUT4), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n254), .B1(new_n249), .B2(new_n250), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n220), .A2(new_n244), .A3(KEYINPUT4), .A4(new_n232), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n255), .A2(new_n256), .A3(new_n203), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n246), .A2(new_n247), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n242), .B1(new_n258), .B2(new_n233), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n223), .A2(new_n226), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n230), .B1(G155gat), .B2(G162gat), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n221), .B1(new_n261), .B2(new_n233), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(KEYINPUT3), .B1(new_n259), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT3), .ZN(new_n265));
  OAI211_X1 g064(.A(new_n232), .B(new_n265), .C1(new_n248), .C2(new_n242), .ZN(new_n266));
  AND3_X1   g065(.A1(new_n264), .A2(new_n266), .A3(new_n250), .ZN(new_n267));
  OAI211_X1 g066(.A(new_n252), .B(KEYINPUT5), .C1(new_n257), .C2(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n264), .A2(new_n266), .A3(new_n250), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n270), .B1(new_n249), .B2(new_n250), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n220), .A2(new_n244), .A3(new_n232), .A4(new_n253), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n204), .A2(KEYINPUT5), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n269), .A2(new_n271), .A3(new_n272), .A4(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n268), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(G57gat), .B(G85gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n276), .B(KEYINPUT80), .ZN(new_n277));
  XNOR2_X1  g076(.A(G1gat), .B(G29gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n275), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT6), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n268), .A2(new_n281), .A3(new_n274), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n275), .A2(KEYINPUT6), .A3(new_n282), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(G226gat), .A2(G233gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n289), .B(KEYINPUT73), .ZN(new_n290));
  NOR2_X1   g089(.A1(G169gat), .A2(G176gat), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT26), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(G169gat), .A2(G176gat), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n295), .A2(KEYINPUT26), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n293), .B1(new_n296), .B2(new_n291), .ZN(new_n297));
  NAND2_X1  g096(.A1(G183gat), .A2(G190gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(G183gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT27), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT27), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(G183gat), .ZN(new_n303));
  INV_X1    g102(.A(G190gat), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n301), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT68), .ZN(new_n306));
  XNOR2_X1  g105(.A(KEYINPUT27), .B(G183gat), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT68), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n307), .A2(new_n308), .A3(new_n304), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  OR2_X1    g109(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n306), .A2(new_n309), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n299), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n295), .B1(KEYINPUT23), .B2(new_n291), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT23), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n317), .B1(G169gat), .B2(G176gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n300), .A2(new_n304), .ZN(new_n319));
  NAND3_X1  g118(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT65), .ZN(new_n322));
  OAI211_X1 g121(.A(new_n319), .B(new_n320), .C1(new_n321), .C2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n321), .A2(new_n322), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n316), .B(new_n318), .C1(new_n323), .C2(new_n325), .ZN(new_n326));
  XOR2_X1   g125(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n327));
  INV_X1    g126(.A(new_n321), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n328), .A2(new_n319), .A3(new_n320), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n291), .A2(KEYINPUT23), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT66), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n330), .A2(new_n331), .A3(new_n294), .ZN(new_n332));
  AND2_X1   g131(.A1(new_n329), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n318), .A2(KEYINPUT25), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n330), .A2(new_n294), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n334), .B1(new_n335), .B2(KEYINPUT66), .ZN(new_n336));
  AOI22_X1  g135(.A1(new_n326), .A2(new_n327), .B1(new_n333), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n290), .B1(new_n315), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(G211gat), .A2(G218gat), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT22), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(G204gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(G197gat), .ZN(new_n343));
  INV_X1    g142(.A(G197gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(G204gat), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n341), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  XOR2_X1   g145(.A(G211gat), .B(G218gat), .Z(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(G211gat), .B(G218gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(G197gat), .B(G204gat), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n349), .A2(new_n350), .A3(new_n341), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(KEYINPUT72), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT72), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n348), .A2(new_n351), .A3(new_n354), .ZN(new_n355));
  AND2_X1   g154(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  AND2_X1   g155(.A1(new_n297), .A2(new_n298), .ZN(new_n357));
  AND3_X1   g156(.A1(new_n306), .A2(new_n309), .A3(new_n313), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n313), .B1(new_n306), .B2(new_n309), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n335), .A2(KEYINPUT66), .ZN(new_n361));
  INV_X1    g160(.A(new_n334), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n361), .A2(new_n362), .A3(new_n329), .A4(new_n332), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n330), .A2(new_n294), .A3(new_n318), .ZN(new_n364));
  INV_X1    g163(.A(new_n323), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n364), .B1(new_n365), .B2(new_n324), .ZN(new_n366));
  INV_X1    g165(.A(new_n327), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n363), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT29), .B1(new_n360), .B2(new_n368), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n338), .B(new_n356), .C1(new_n369), .C2(new_n290), .ZN(new_n370));
  XNOR2_X1  g169(.A(G8gat), .B(G36gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(G64gat), .B(G92gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n371), .B(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n290), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n375), .B1(new_n360), .B2(new_n368), .ZN(new_n376));
  XNOR2_X1  g175(.A(KEYINPUT74), .B(KEYINPUT29), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n377), .B1(new_n315), .B2(new_n337), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n376), .B1(new_n378), .B2(new_n375), .ZN(new_n379));
  OAI211_X1 g178(.A(new_n370), .B(new_n374), .C1(new_n379), .C2(new_n356), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT75), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT30), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n353), .A2(new_n355), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n360), .A2(new_n368), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n290), .B1(new_n385), .B2(new_n377), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n384), .B1(new_n386), .B2(new_n376), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n387), .A2(KEYINPUT75), .A3(new_n370), .A4(new_n374), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n382), .A2(new_n383), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n374), .B1(new_n387), .B2(new_n370), .ZN(new_n390));
  INV_X1    g189(.A(new_n380), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n390), .B1(new_n391), .B2(KEYINPUT30), .ZN(new_n392));
  AND4_X1   g191(.A1(new_n202), .A2(new_n288), .A3(new_n389), .A4(new_n392), .ZN(new_n393));
  XOR2_X1   g192(.A(KEYINPUT31), .B(G50gat), .Z(new_n394));
  AOI21_X1  g193(.A(KEYINPUT29), .B1(new_n348), .B2(new_n351), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT83), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n265), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  AOI211_X1 g196(.A(KEYINPUT83), .B(KEYINPUT29), .C1(new_n348), .C2(new_n351), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n249), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n266), .A2(new_n377), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(new_n384), .ZN(new_n401));
  NAND2_X1  g200(.A1(G228gat), .A2(G233gat), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n399), .A2(new_n401), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(KEYINPUT84), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT84), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n399), .A2(new_n401), .A3(new_n406), .A4(new_n403), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n238), .A2(new_n239), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n409), .B1(KEYINPUT77), .B2(new_n242), .ZN(new_n410));
  INV_X1    g209(.A(new_n262), .ZN(new_n411));
  AOI22_X1  g210(.A1(new_n241), .A2(new_n243), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n352), .A2(new_n377), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n412), .B1(new_n265), .B2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT82), .ZN(new_n416));
  AND3_X1   g215(.A1(new_n400), .A2(new_n416), .A3(new_n384), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n416), .B1(new_n400), .B2(new_n384), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n415), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n402), .B(KEYINPUT81), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(G22gat), .ZN(new_n422));
  AND3_X1   g221(.A1(new_n408), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n422), .B1(new_n408), .B2(new_n421), .ZN(new_n424));
  XNOR2_X1  g223(.A(G78gat), .B(G106gat), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NOR3_X1   g225(.A1(new_n423), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT29), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n346), .A2(new_n347), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n349), .B1(new_n341), .B2(new_n350), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n428), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(KEYINPUT83), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n395), .A2(new_n396), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n432), .A2(new_n265), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n402), .B1(new_n434), .B2(new_n249), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n406), .B1(new_n435), .B2(new_n401), .ZN(new_n436));
  INV_X1    g235(.A(new_n407), .ZN(new_n437));
  INV_X1    g236(.A(new_n377), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n438), .B1(new_n412), .B2(new_n265), .ZN(new_n439));
  OAI21_X1  g238(.A(KEYINPUT82), .B1(new_n439), .B2(new_n356), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n400), .A2(new_n416), .A3(new_n384), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n414), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n420), .ZN(new_n443));
  OAI22_X1  g242(.A1(new_n436), .A2(new_n437), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(G22gat), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n408), .A2(new_n421), .A3(new_n422), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n425), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n394), .B1(new_n427), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n426), .B1(new_n423), .B2(new_n424), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n445), .A2(new_n446), .A3(new_n425), .ZN(new_n450));
  INV_X1    g249(.A(new_n394), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(G227gat), .ZN(new_n453));
  INV_X1    g252(.A(G233gat), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n385), .A2(new_n220), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n360), .A2(new_n250), .A3(new_n368), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n455), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n458), .B(KEYINPUT34), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n456), .A2(new_n455), .A3(new_n457), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT33), .ZN(new_n461));
  XOR2_X1   g260(.A(G15gat), .B(G43gat), .Z(new_n462));
  XNOR2_X1  g261(.A(G71gat), .B(G99gat), .ZN(new_n463));
  XNOR2_X1  g262(.A(new_n462), .B(new_n463), .ZN(new_n464));
  XNOR2_X1  g263(.A(new_n464), .B(KEYINPUT71), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n460), .B(KEYINPUT32), .C1(new_n461), .C2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n460), .A2(KEYINPUT32), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n460), .A2(new_n461), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n467), .A2(new_n468), .A3(new_n464), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n459), .A2(new_n466), .A3(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n459), .B1(new_n466), .B2(new_n469), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n393), .A2(new_n448), .A3(new_n452), .A4(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT87), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AND3_X1   g275(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n451), .B1(new_n449), .B2(new_n450), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n479), .A2(KEYINPUT87), .A3(new_n473), .A4(new_n393), .ZN(new_n480));
  AND3_X1   g279(.A1(new_n288), .A2(new_n389), .A3(new_n392), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n448), .A2(new_n481), .A3(new_n452), .A4(new_n473), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT35), .ZN(new_n483));
  AOI22_X1  g282(.A1(new_n476), .A2(new_n480), .B1(new_n483), .B2(KEYINPUT88), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT88), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n482), .A2(new_n485), .A3(KEYINPUT35), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT37), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n370), .B(new_n487), .C1(new_n379), .C2(new_n356), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(new_n373), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT38), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n338), .B(new_n384), .C1(new_n369), .C2(new_n290), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT37), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n378), .A2(new_n375), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n384), .B1(new_n493), .B2(new_n338), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n490), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n489), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n382), .A2(new_n388), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AND2_X1   g297(.A1(new_n286), .A2(new_n287), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n487), .B1(new_n387), .B2(new_n370), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT38), .B1(new_n489), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n498), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n389), .A2(new_n392), .ZN(new_n503));
  INV_X1    g302(.A(new_n283), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n271), .A2(new_n272), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n204), .B1(new_n267), .B2(new_n505), .ZN(new_n506));
  OR2_X1    g305(.A1(new_n245), .A2(new_n251), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n506), .B(KEYINPUT39), .C1(new_n204), .C2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT39), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n509), .B(new_n204), .C1(new_n267), .C2(new_n505), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT85), .ZN(new_n511));
  AND3_X1   g310(.A1(new_n510), .A2(new_n511), .A3(new_n281), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n511), .B1(new_n510), .B2(new_n281), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n508), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT40), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n504), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OAI211_X1 g315(.A(KEYINPUT40), .B(new_n508), .C1(new_n512), .C2(new_n513), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n503), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n448), .A2(new_n502), .A3(new_n518), .A4(new_n452), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n519), .A2(KEYINPUT86), .ZN(new_n520));
  OAI22_X1  g319(.A1(new_n477), .A2(new_n478), .B1(new_n499), .B2(new_n503), .ZN(new_n521));
  NOR3_X1   g320(.A1(new_n471), .A2(new_n472), .A3(KEYINPUT36), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT36), .ZN(new_n523));
  INV_X1    g322(.A(new_n459), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n469), .A2(new_n466), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n523), .B1(new_n526), .B2(new_n470), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n522), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n521), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n520), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n519), .A2(KEYINPUT86), .ZN(new_n531));
  AOI22_X1  g330(.A1(new_n484), .A2(new_n486), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  AND2_X1   g331(.A1(G232gat), .A2(G233gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT41), .ZN(new_n534));
  XNOR2_X1  g333(.A(G99gat), .B(G106gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(KEYINPUT95), .ZN(new_n536));
  NAND2_X1  g335(.A1(G85gat), .A2(G92gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(KEYINPUT7), .ZN(new_n538));
  INV_X1    g337(.A(G99gat), .ZN(new_n539));
  INV_X1    g338(.A(G106gat), .ZN(new_n540));
  OAI21_X1  g339(.A(KEYINPUT8), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n538), .B(new_n541), .C1(G85gat), .C2(G92gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n536), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT96), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n536), .A2(new_n542), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n536), .A2(new_n542), .A3(KEYINPUT96), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NOR2_X1   g347(.A1(G29gat), .A2(G36gat), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT14), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(G29gat), .A2(G36gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(G43gat), .B(G50gat), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n553), .A2(KEYINPUT15), .A3(new_n554), .ZN(new_n555));
  OR2_X1    g354(.A1(new_n554), .A2(KEYINPUT15), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n554), .A2(KEYINPUT15), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n552), .B(KEYINPUT90), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n556), .A2(new_n551), .A3(new_n557), .A4(new_n558), .ZN(new_n559));
  AND2_X1   g358(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n534), .B1(new_n548), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(KEYINPUT17), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT91), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n555), .A2(new_n559), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT17), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  AOI211_X1 g365(.A(KEYINPUT91), .B(KEYINPUT17), .C1(new_n555), .C2(new_n559), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n562), .B(new_n548), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  OR2_X1    g367(.A1(new_n568), .A2(KEYINPUT97), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(KEYINPUT97), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n561), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G190gat), .B(G218gat), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT98), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n571), .A2(KEYINPUT98), .A3(new_n573), .ZN(new_n577));
  OR2_X1    g376(.A1(new_n571), .A2(new_n573), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n533), .A2(KEYINPUT41), .ZN(new_n580));
  XNOR2_X1  g379(.A(G134gat), .B(G162gat), .ZN(new_n581));
  XOR2_X1   g380(.A(new_n580), .B(new_n581), .Z(new_n582));
  NAND2_X1  g381(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n582), .B1(new_n571), .B2(new_n573), .ZN(new_n584));
  AOI21_X1  g383(.A(KEYINPUT99), .B1(new_n578), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n578), .A2(KEYINPUT99), .A3(new_n584), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n583), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT16), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n589), .A2(G1gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(G15gat), .B(G22gat), .ZN(new_n591));
  MUX2_X1   g390(.A(G1gat), .B(new_n590), .S(new_n591), .Z(new_n592));
  INV_X1    g391(.A(G8gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  AND2_X1   g393(.A1(G71gat), .A2(G78gat), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n595), .A2(KEYINPUT9), .ZN(new_n596));
  XNOR2_X1  g395(.A(G57gat), .B(G64gat), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(G71gat), .A2(G78gat), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(KEYINPUT94), .A2(KEYINPUT9), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  OAI211_X1 g402(.A(new_n601), .B(new_n600), .C1(new_n596), .C2(new_n597), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n594), .B1(KEYINPUT21), .B2(new_n606), .ZN(new_n607));
  XOR2_X1   g406(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n608));
  INV_X1    g407(.A(KEYINPUT21), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  AND2_X1   g409(.A1(G231gat), .A2(G233gat), .ZN(new_n611));
  OR2_X1    g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(new_n611), .ZN(new_n613));
  XNOR2_X1  g412(.A(G127gat), .B(G155gat), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n614), .B1(new_n612), .B2(new_n613), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n608), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NOR3_X1   g418(.A1(new_n616), .A2(new_n617), .A3(new_n608), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n607), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n620), .ZN(new_n622));
  INV_X1    g421(.A(new_n607), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n622), .A2(new_n623), .A3(new_n618), .ZN(new_n624));
  XNOR2_X1  g423(.A(G183gat), .B(G211gat), .ZN(new_n625));
  AND3_X1   g424(.A1(new_n621), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n625), .B1(new_n621), .B2(new_n624), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n588), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n592), .B(G8gat), .ZN(new_n630));
  OAI211_X1 g429(.A(new_n630), .B(new_n562), .C1(new_n566), .C2(new_n567), .ZN(new_n631));
  NAND2_X1  g430(.A1(G229gat), .A2(G233gat), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n594), .A2(new_n564), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n631), .A2(KEYINPUT18), .A3(new_n632), .A4(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT93), .ZN(new_n635));
  OR2_X1    g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT92), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n630), .A2(new_n560), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n633), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n632), .B(KEYINPUT13), .Z(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n638), .A2(new_n639), .A3(new_n643), .ZN(new_n644));
  AND2_X1   g443(.A1(new_n631), .A2(new_n633), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(new_n632), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT18), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n638), .A2(new_n643), .A3(new_n648), .ZN(new_n649));
  XOR2_X1   g448(.A(G113gat), .B(G141gat), .Z(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT11), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT89), .ZN(new_n652));
  XNOR2_X1  g451(.A(G169gat), .B(G197gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT12), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n644), .A2(new_n649), .A3(new_n656), .ZN(new_n657));
  AOI22_X1  g456(.A1(new_n636), .A2(new_n637), .B1(new_n641), .B2(new_n642), .ZN(new_n658));
  OAI211_X1 g457(.A(new_n658), .B(new_n648), .C1(new_n639), .C2(new_n655), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g459(.A(G120gat), .B(G148gat), .Z(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT100), .ZN(new_n662));
  XOR2_X1   g461(.A(G176gat), .B(G204gat), .Z(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n605), .B1(new_n536), .B2(new_n542), .ZN(new_n665));
  AOI22_X1  g464(.A1(new_n548), .A2(new_n605), .B1(new_n665), .B2(new_n546), .ZN(new_n666));
  NAND2_X1  g465(.A1(G230gat), .A2(G233gat), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n548), .A2(new_n605), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT10), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n665), .A2(new_n546), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  OR3_X1    g471(.A1(new_n548), .A2(new_n670), .A3(new_n605), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AOI211_X1 g473(.A(new_n664), .B(new_n668), .C1(new_n674), .C2(new_n667), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT101), .ZN(new_n677));
  NOR3_X1   g476(.A1(new_n548), .A2(new_n670), .A3(new_n605), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n678), .B1(new_n670), .B2(new_n666), .ZN(new_n679));
  INV_X1    g478(.A(new_n667), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n677), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n674), .A2(KEYINPUT101), .A3(new_n667), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n668), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n664), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n676), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n629), .A2(new_n660), .A3(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n532), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(new_n499), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g489(.A1(new_n688), .A2(new_n503), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(G8gat), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT42), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n589), .A2(new_n593), .ZN(new_n694));
  NAND2_X1  g493(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n688), .A2(new_n503), .A3(new_n694), .A4(new_n695), .ZN(new_n696));
  AND3_X1   g495(.A1(new_n696), .A2(KEYINPUT102), .A3(new_n693), .ZN(new_n697));
  AOI21_X1  g496(.A(KEYINPUT102), .B1(new_n696), .B2(new_n693), .ZN(new_n698));
  OAI221_X1 g497(.A(new_n692), .B1(new_n693), .B2(new_n696), .C1(new_n697), .C2(new_n698), .ZN(G1325gat));
  INV_X1    g498(.A(G15gat), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n688), .A2(new_n700), .A3(new_n473), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n532), .A2(new_n528), .A3(new_n687), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n701), .B1(new_n702), .B2(new_n700), .ZN(G1326gat));
  INV_X1    g502(.A(new_n479), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g504(.A(KEYINPUT43), .B(G22gat), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n705), .B(new_n706), .ZN(G1327gat));
  NAND2_X1  g506(.A1(new_n480), .A2(new_n476), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n483), .A2(KEYINPUT88), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n708), .A2(new_n486), .A3(new_n709), .ZN(new_n710));
  OR2_X1    g509(.A1(new_n519), .A2(KEYINPUT86), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n711), .A2(new_n531), .A3(new_n521), .A4(new_n528), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n657), .A2(new_n659), .ZN(new_n714));
  INV_X1    g513(.A(new_n628), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n714), .A2(new_n715), .A3(new_n685), .ZN(new_n716));
  AND3_X1   g515(.A1(new_n713), .A2(new_n588), .A3(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(G29gat), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n717), .A2(new_n718), .A3(new_n499), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT45), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n721));
  INV_X1    g520(.A(new_n588), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n721), .B1(new_n532), .B2(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n713), .A2(KEYINPUT44), .A3(new_n588), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n725), .A2(new_n716), .ZN(new_n726));
  AND2_X1   g525(.A1(new_n726), .A2(new_n499), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n720), .B1(new_n727), .B2(new_n718), .ZN(G1328gat));
  INV_X1    g527(.A(G36gat), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n717), .A2(new_n729), .A3(new_n503), .ZN(new_n730));
  XOR2_X1   g529(.A(new_n730), .B(KEYINPUT46), .Z(new_n731));
  AND2_X1   g530(.A1(new_n726), .A2(new_n503), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n731), .B1(new_n732), .B2(new_n729), .ZN(G1329gat));
  INV_X1    g532(.A(G43gat), .ZN(new_n734));
  INV_X1    g533(.A(new_n528), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n723), .A2(new_n735), .A3(new_n724), .A4(new_n716), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT104), .ZN(new_n737));
  OR2_X1    g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(new_n737), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n734), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n473), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n741), .A2(G43gat), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n717), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(KEYINPUT47), .ZN(new_n744));
  AOI22_X1  g543(.A1(new_n736), .A2(G43gat), .B1(new_n717), .B2(new_n742), .ZN(new_n745));
  XNOR2_X1  g544(.A(KEYINPUT103), .B(KEYINPUT47), .ZN(new_n746));
  OAI22_X1  g545(.A1(new_n740), .A2(new_n744), .B1(new_n745), .B2(new_n746), .ZN(G1330gat));
  NAND4_X1  g546(.A1(new_n723), .A2(new_n704), .A3(new_n724), .A4(new_n716), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(G50gat), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n479), .A2(G50gat), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n717), .A2(new_n750), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n749), .B(new_n751), .C1(KEYINPUT105), .C2(KEYINPUT48), .ZN(new_n752));
  NAND2_X1  g551(.A1(KEYINPUT105), .A2(KEYINPUT48), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n752), .B(new_n753), .ZN(G1331gat));
  NOR4_X1   g553(.A1(new_n588), .A2(new_n628), .A3(new_n660), .A4(new_n686), .ZN(new_n755));
  AND2_X1   g554(.A1(new_n713), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n499), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g557(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n759));
  AND3_X1   g558(.A1(new_n756), .A2(new_n503), .A3(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n760), .B(new_n761), .ZN(G1333gat));
  INV_X1    g561(.A(G71gat), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n763), .B1(new_n756), .B2(new_n735), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT107), .ZN(new_n765));
  AND4_X1   g564(.A1(new_n763), .A2(new_n713), .A3(new_n473), .A4(new_n755), .ZN(new_n766));
  OR3_X1    g565(.A1(new_n764), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n765), .B1(new_n764), .B2(new_n766), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  XOR2_X1   g568(.A(KEYINPUT106), .B(KEYINPUT50), .Z(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(new_n770), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n767), .A2(new_n768), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n773), .ZN(G1334gat));
  NAND2_X1  g573(.A1(new_n756), .A2(new_n704), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(G78gat), .ZN(G1335gat));
  NAND3_X1  g575(.A1(new_n714), .A2(KEYINPUT108), .A3(new_n628), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT108), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n778), .B1(new_n715), .B2(new_n660), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n780), .A2(new_n686), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n725), .A2(new_n499), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(G85gat), .ZN(new_n783));
  INV_X1    g582(.A(new_n780), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n713), .A2(new_n588), .A3(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT51), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n288), .A2(G85gat), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n787), .A2(new_n685), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n783), .A2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT109), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n783), .A2(KEYINPUT109), .A3(new_n789), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(G1336gat));
  INV_X1    g593(.A(G92gat), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n685), .A2(new_n795), .A3(new_n503), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT110), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n787), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT52), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n723), .A2(new_n503), .A3(new_n724), .A4(new_n781), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(G92gat), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n799), .A2(new_n800), .A3(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT112), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n799), .A2(KEYINPUT112), .A3(new_n800), .A4(new_n802), .ZN(new_n806));
  AOI211_X1 g605(.A(new_n722), .B(new_n780), .C1(new_n710), .C2(new_n712), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT111), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n786), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n785), .A2(KEYINPUT111), .A3(KEYINPUT51), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n809), .A2(new_n798), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n802), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(KEYINPUT52), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n805), .A2(new_n806), .A3(new_n813), .ZN(G1337gat));
  NAND4_X1  g613(.A1(new_n787), .A2(new_n539), .A3(new_n473), .A4(new_n685), .ZN(new_n815));
  AND3_X1   g614(.A1(new_n725), .A2(new_n735), .A3(new_n781), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n815), .B1(new_n816), .B2(new_n539), .ZN(G1338gat));
  NOR3_X1   g616(.A1(new_n479), .A2(G106gat), .A3(new_n686), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n809), .A2(new_n810), .A3(new_n818), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n723), .A2(new_n704), .A3(new_n724), .A4(new_n781), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(G106gat), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(KEYINPUT53), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT113), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT114), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n820), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n820), .A2(new_n826), .ZN(new_n828));
  OAI21_X1  g627(.A(G106gat), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(KEYINPUT53), .B1(new_n787), .B2(new_n818), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n822), .A2(KEYINPUT113), .A3(KEYINPUT53), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n825), .A2(new_n831), .A3(new_n832), .ZN(G1339gat));
  NOR4_X1   g632(.A1(new_n588), .A2(new_n660), .A3(new_n628), .A4(new_n685), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n638), .A2(new_n643), .A3(new_n655), .A4(new_n648), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n645), .A2(new_n632), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n641), .A2(new_n642), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n654), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT115), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n839), .A2(new_n840), .A3(new_n685), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n685), .A2(new_n835), .A3(new_n838), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(KEYINPUT115), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n844), .B1(new_n674), .B2(new_n667), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n679), .A2(new_n680), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n684), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n681), .A2(new_n844), .A3(new_n682), .ZN(new_n848));
  AOI21_X1  g647(.A(KEYINPUT55), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n849), .A2(new_n675), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n847), .A2(new_n848), .A3(KEYINPUT55), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  OAI211_X1 g651(.A(new_n841), .B(new_n843), .C1(new_n714), .C2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n722), .ZN(new_n854));
  INV_X1    g653(.A(new_n851), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n855), .A2(new_n849), .A3(new_n675), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n588), .A2(new_n856), .A3(new_n839), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n834), .B1(new_n858), .B2(new_n628), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n499), .A2(new_n389), .A3(new_n392), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n704), .A2(new_n741), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(new_n660), .ZN(new_n865));
  XNOR2_X1  g664(.A(new_n865), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g665(.A1(new_n864), .A2(new_n685), .ZN(new_n867));
  XNOR2_X1  g666(.A(new_n867), .B(G120gat), .ZN(G1341gat));
  NOR2_X1   g667(.A1(new_n863), .A2(new_n628), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n869), .B(new_n209), .ZN(G1342gat));
  NOR3_X1   g669(.A1(new_n722), .A2(new_n704), .A3(new_n741), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n861), .A2(new_n211), .A3(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n872), .A2(KEYINPUT56), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n873), .B(KEYINPUT116), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n872), .A2(KEYINPUT56), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n861), .A2(new_n871), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(G134gat), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n874), .A2(new_n875), .A3(new_n877), .ZN(G1343gat));
  NOR2_X1   g677(.A1(new_n735), .A2(new_n860), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT57), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n479), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n856), .A2(new_n660), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(new_n842), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(new_n722), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n715), .B1(new_n884), .B2(new_n857), .ZN(new_n885));
  OAI211_X1 g684(.A(KEYINPUT117), .B(new_n881), .C1(new_n885), .C2(new_n834), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT117), .ZN(new_n887));
  AOI22_X1  g686(.A1(new_n856), .A2(new_n660), .B1(new_n685), .B2(new_n839), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n857), .B1(new_n888), .B2(new_n588), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n834), .B1(new_n889), .B2(new_n628), .ZN(new_n890));
  INV_X1    g689(.A(new_n881), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n887), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n886), .A2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(new_n834), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n835), .A2(new_n838), .ZN(new_n895));
  AND3_X1   g694(.A1(new_n578), .A2(KEYINPUT99), .A3(new_n584), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n896), .A2(new_n585), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n895), .B1(new_n897), .B2(new_n583), .ZN(new_n898));
  AOI22_X1  g697(.A1(new_n853), .A2(new_n722), .B1(new_n856), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n894), .B1(new_n899), .B2(new_n715), .ZN(new_n900));
  AOI21_X1  g699(.A(KEYINPUT57), .B1(new_n900), .B2(new_n704), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n660), .B(new_n879), .C1(new_n893), .C2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(G141gat), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n735), .A2(new_n479), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n861), .A2(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n906), .A2(new_n236), .A3(new_n660), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n903), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(KEYINPUT58), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT58), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n903), .A2(new_n907), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n909), .A2(new_n911), .ZN(G1344gat));
  NOR4_X1   g711(.A1(new_n686), .A2(G148gat), .A3(new_n288), .A4(new_n503), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n900), .A2(new_n904), .A3(new_n913), .ZN(new_n914));
  OAI211_X1 g713(.A(new_n685), .B(new_n879), .C1(new_n893), .C2(new_n901), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT118), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n237), .A2(KEYINPUT59), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n880), .B1(new_n900), .B2(new_n704), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n704), .A2(new_n880), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n890), .A2(new_n920), .ZN(new_n921));
  XOR2_X1   g720(.A(new_n879), .B(KEYINPUT119), .Z(new_n922));
  NOR4_X1   g721(.A1(new_n919), .A2(new_n921), .A3(new_n686), .A4(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(KEYINPUT59), .B1(new_n923), .B2(new_n237), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n918), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n916), .B1(new_n915), .B2(new_n917), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n914), .B1(new_n925), .B2(new_n926), .ZN(G1345gat));
  OAI211_X1 g726(.A(new_n715), .B(new_n879), .C1(new_n893), .C2(new_n901), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(G155gat), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n906), .A2(new_n227), .A3(new_n715), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT120), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n929), .A2(new_n930), .A3(KEYINPUT120), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(G1346gat));
  OAI211_X1 g734(.A(new_n588), .B(new_n879), .C1(new_n893), .C2(new_n901), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(G162gat), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n906), .A2(new_n228), .A3(new_n588), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT121), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n937), .A2(new_n938), .A3(KEYINPUT121), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(G1347gat));
  NAND2_X1  g742(.A1(new_n503), .A2(new_n288), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n859), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(new_n862), .ZN(new_n946));
  INV_X1    g745(.A(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(G169gat), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n947), .A2(new_n948), .A3(new_n660), .ZN(new_n949));
  OAI21_X1  g748(.A(G169gat), .B1(new_n946), .B2(new_n714), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(KEYINPUT122), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT122), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n949), .A2(new_n953), .A3(new_n950), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n952), .A2(new_n954), .ZN(G1348gat));
  NAND2_X1  g754(.A1(new_n947), .A2(new_n685), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n956), .B(G176gat), .ZN(G1349gat));
  OAI21_X1  g756(.A(G183gat), .B1(new_n946), .B2(new_n628), .ZN(new_n958));
  NAND4_X1  g757(.A1(new_n945), .A2(new_n307), .A3(new_n862), .A4(new_n715), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT60), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n961), .A2(KEYINPUT123), .ZN(new_n962));
  XNOR2_X1  g761(.A(new_n960), .B(new_n962), .ZN(G1350gat));
  INV_X1    g762(.A(KEYINPUT61), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n946), .A2(new_n722), .ZN(new_n965));
  INV_X1    g764(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n964), .B1(new_n966), .B2(G190gat), .ZN(new_n967));
  NOR3_X1   g766(.A1(new_n965), .A2(KEYINPUT61), .A3(new_n304), .ZN(new_n968));
  OAI22_X1  g767(.A1(new_n967), .A2(new_n968), .B1(G190gat), .B2(new_n966), .ZN(G1351gat));
  NOR2_X1   g768(.A1(new_n735), .A2(new_n944), .ZN(new_n970));
  INV_X1    g769(.A(new_n970), .ZN(new_n971));
  OR2_X1    g770(.A1(new_n890), .A2(new_n920), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n842), .B(new_n840), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n588), .B1(new_n973), .B2(new_n882), .ZN(new_n974));
  INV_X1    g773(.A(new_n857), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n628), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n479), .B1(new_n976), .B2(new_n894), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n972), .B1(new_n977), .B2(new_n880), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT124), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n971), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  OAI211_X1 g779(.A(new_n972), .B(KEYINPUT124), .C1(new_n977), .C2(new_n880), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NOR3_X1   g781(.A1(new_n982), .A2(new_n344), .A3(new_n714), .ZN(new_n983));
  INV_X1    g782(.A(new_n944), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n900), .A2(new_n904), .A3(new_n984), .ZN(new_n985));
  INV_X1    g784(.A(new_n985), .ZN(new_n986));
  AOI21_X1  g785(.A(G197gat), .B1(new_n986), .B2(new_n660), .ZN(new_n987));
  NOR2_X1   g786(.A1(new_n983), .A2(new_n987), .ZN(G1352gat));
  OAI21_X1  g787(.A(new_n979), .B1(new_n919), .B2(new_n921), .ZN(new_n989));
  NAND4_X1  g788(.A1(new_n989), .A2(new_n981), .A3(new_n685), .A4(new_n970), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n990), .A2(KEYINPUT126), .ZN(new_n991));
  INV_X1    g790(.A(KEYINPUT126), .ZN(new_n992));
  NAND4_X1  g791(.A1(new_n980), .A2(new_n992), .A3(new_n685), .A4(new_n981), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n991), .A2(new_n993), .A3(G204gat), .ZN(new_n994));
  NOR3_X1   g793(.A1(new_n985), .A2(G204gat), .A3(new_n686), .ZN(new_n995));
  INV_X1    g794(.A(KEYINPUT62), .ZN(new_n996));
  OAI21_X1  g795(.A(KEYINPUT125), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g796(.A(KEYINPUT125), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n685), .A2(new_n342), .ZN(new_n999));
  OAI211_X1 g798(.A(new_n998), .B(KEYINPUT62), .C1(new_n985), .C2(new_n999), .ZN(new_n1000));
  AOI22_X1  g799(.A1(new_n997), .A2(new_n1000), .B1(new_n996), .B2(new_n995), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n994), .A2(new_n1001), .ZN(G1353gat));
  INV_X1    g801(.A(G211gat), .ZN(new_n1003));
  INV_X1    g802(.A(new_n978), .ZN(new_n1004));
  NOR2_X1   g803(.A1(new_n971), .A2(new_n628), .ZN(new_n1005));
  AOI21_X1  g804(.A(new_n1003), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g805(.A(KEYINPUT63), .ZN(new_n1007));
  OR2_X1    g806(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1009));
  NOR3_X1   g808(.A1(new_n985), .A2(G211gat), .A3(new_n628), .ZN(new_n1010));
  XNOR2_X1  g809(.A(new_n1010), .B(KEYINPUT127), .ZN(new_n1011));
  NAND3_X1  g810(.A1(new_n1008), .A2(new_n1009), .A3(new_n1011), .ZN(G1354gat));
  OAI21_X1  g811(.A(G218gat), .B1(new_n982), .B2(new_n722), .ZN(new_n1013));
  OR2_X1    g812(.A1(new_n722), .A2(G218gat), .ZN(new_n1014));
  OAI21_X1  g813(.A(new_n1013), .B1(new_n985), .B2(new_n1014), .ZN(G1355gat));
endmodule


