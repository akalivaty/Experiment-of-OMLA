//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 1 1 0 0 1 0 0 1 0 1 0 1 0 0 0 1 1 0 1 0 1 1 0 0 0 0 1 0 0 1 1 0 0 1 0 0 1 1 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n751,
    new_n752, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n854, new_n855, new_n856,
    new_n857, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963;
  INV_X1    g000(.A(KEYINPUT85), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT5), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT76), .B(G148gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G141gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT77), .ZN(new_n206));
  INV_X1    g005(.A(G141gat), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n206), .B1(new_n207), .B2(G148gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n205), .A2(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(G155gat), .B(G162gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n204), .A2(new_n206), .A3(G141gat), .ZN(new_n211));
  INV_X1    g010(.A(G162gat), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT2), .B1(new_n212), .B2(KEYINPUT78), .ZN(new_n213));
  NAND4_X1  g012(.A1(new_n209), .A2(new_n210), .A3(new_n211), .A4(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT3), .ZN(new_n215));
  XNOR2_X1  g014(.A(G141gat), .B(G148gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n216), .A2(KEYINPUT2), .ZN(new_n217));
  OR2_X1    g016(.A1(new_n217), .A2(new_n210), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n214), .A2(new_n215), .A3(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n215), .B1(new_n214), .B2(new_n218), .ZN(new_n221));
  XNOR2_X1  g020(.A(G127gat), .B(G134gat), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n222), .B(KEYINPUT68), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT1), .ZN(new_n224));
  INV_X1    g023(.A(G113gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n225), .A2(G120gat), .ZN(new_n226));
  INV_X1    g025(.A(G120gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n227), .A2(G113gat), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n224), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  OR3_X1    g028(.A1(new_n225), .A2(KEYINPUT69), .A3(G120gat), .ZN(new_n230));
  OAI21_X1  g029(.A(KEYINPUT69), .B1(new_n225), .B2(G120gat), .ZN(new_n231));
  XNOR2_X1  g030(.A(KEYINPUT70), .B(G113gat), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n230), .B(new_n231), .C1(new_n232), .C2(new_n227), .ZN(new_n233));
  AND2_X1   g032(.A1(new_n222), .A2(new_n224), .ZN(new_n234));
  AOI22_X1  g033(.A1(new_n223), .A2(new_n229), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NOR3_X1   g034(.A1(new_n220), .A2(new_n221), .A3(new_n235), .ZN(new_n236));
  AND2_X1   g035(.A1(new_n222), .A2(KEYINPUT68), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n222), .A2(KEYINPUT68), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n229), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n233), .A2(new_n234), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n214), .A2(new_n239), .A3(new_n218), .A4(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT4), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  XOR2_X1   g042(.A(KEYINPUT79), .B(KEYINPUT4), .Z(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n235), .A2(new_n218), .A3(new_n214), .A4(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n203), .B1(new_n236), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n221), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n239), .A2(new_n240), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n249), .A2(new_n250), .A3(new_n219), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n214), .A2(new_n218), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n253), .A2(KEYINPUT4), .A3(new_n235), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n241), .A2(new_n244), .ZN(new_n255));
  NAND2_X1  g054(.A1(G225gat), .A2(G233gat), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n257), .A2(new_n203), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n251), .A2(new_n254), .A3(new_n255), .A4(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n252), .A2(new_n250), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT80), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n260), .A2(new_n261), .A3(new_n241), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n252), .A2(KEYINPUT80), .A3(new_n250), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n203), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n248), .B(new_n259), .C1(new_n256), .C2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G1gat), .B(G29gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n266), .B(KEYINPUT0), .ZN(new_n267));
  XNOR2_X1  g066(.A(G57gat), .B(G85gat), .ZN(new_n268));
  XOR2_X1   g067(.A(new_n267), .B(new_n268), .Z(new_n269));
  OAI21_X1  g068(.A(new_n202), .B1(new_n265), .B2(new_n269), .ZN(new_n270));
  XOR2_X1   g069(.A(KEYINPUT81), .B(KEYINPUT6), .Z(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n272), .B1(new_n265), .B2(new_n269), .ZN(new_n273));
  AND2_X1   g072(.A1(new_n248), .A2(new_n259), .ZN(new_n274));
  OR2_X1    g073(.A1(new_n264), .A2(new_n256), .ZN(new_n275));
  INV_X1    g074(.A(new_n269), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n274), .A2(new_n275), .A3(KEYINPUT85), .A4(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n270), .A2(new_n273), .A3(new_n277), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n274), .A2(new_n275), .A3(new_n276), .A4(new_n272), .ZN(new_n279));
  AND2_X1   g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT86), .ZN(new_n281));
  NAND3_X1  g080(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n282), .B1(G183gat), .B2(G190gat), .ZN(new_n283));
  AOI21_X1  g082(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n284));
  OAI21_X1  g083(.A(KEYINPUT64), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n284), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT64), .ZN(new_n287));
  INV_X1    g086(.A(G183gat), .ZN(new_n288));
  INV_X1    g087(.A(G190gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n286), .A2(new_n287), .A3(new_n290), .A4(new_n282), .ZN(new_n291));
  INV_X1    g090(.A(G169gat), .ZN(new_n292));
  INV_X1    g091(.A(G176gat), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n292), .A2(new_n293), .A3(KEYINPUT23), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT23), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n295), .B1(G169gat), .B2(G176gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(G169gat), .A2(G176gat), .ZN(new_n297));
  AND3_X1   g096(.A1(new_n294), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n285), .A2(new_n291), .A3(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT65), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT25), .ZN(new_n301));
  AND3_X1   g100(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n300), .B1(new_n299), .B2(new_n301), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n294), .A2(new_n296), .A3(KEYINPUT25), .A4(new_n297), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n283), .B1(KEYINPUT66), .B2(new_n286), .ZN(new_n305));
  OR2_X1    g104(.A1(new_n286), .A2(KEYINPUT66), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NOR3_X1   g106(.A1(new_n302), .A2(new_n303), .A3(new_n307), .ZN(new_n308));
  NOR2_X1   g107(.A1(G169gat), .A2(G176gat), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n309), .A2(KEYINPUT26), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(new_n297), .ZN(new_n311));
  AOI22_X1  g110(.A1(new_n309), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(KEYINPUT27), .B(G183gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(new_n289), .ZN(new_n314));
  XNOR2_X1  g113(.A(KEYINPUT67), .B(KEYINPUT28), .ZN(new_n315));
  OAI211_X1 g114(.A(new_n311), .B(new_n312), .C1(new_n314), .C2(new_n315), .ZN(new_n316));
  AND2_X1   g115(.A1(new_n314), .A2(new_n315), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(KEYINPUT74), .B1(new_n308), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(G226gat), .A2(G233gat), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n299), .A2(new_n301), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(KEYINPUT65), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n324));
  INV_X1    g123(.A(new_n307), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT74), .ZN(new_n327));
  INV_X1    g126(.A(new_n318), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n319), .A2(new_n321), .A3(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(G197gat), .B(G204gat), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT22), .ZN(new_n332));
  INV_X1    g131(.A(G211gat), .ZN(new_n333));
  INV_X1    g132(.A(G218gat), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n332), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  XOR2_X1   g135(.A(G211gat), .B(G218gat), .Z(new_n337));
  XOR2_X1   g136(.A(new_n336), .B(new_n337), .Z(new_n338));
  INV_X1    g137(.A(KEYINPUT73), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n336), .A2(KEYINPUT73), .A3(new_n337), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT29), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n344), .B(new_n320), .C1(new_n308), .C2(new_n318), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n330), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n319), .A2(new_n329), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n321), .B1(new_n347), .B2(new_n344), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n321), .B1(new_n308), .B2(new_n318), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(new_n342), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n346), .B(KEYINPUT37), .C1(new_n348), .C2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n330), .A2(new_n345), .A3(new_n342), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT37), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n349), .A2(new_n343), .ZN(new_n354));
  OAI211_X1 g153(.A(new_n352), .B(new_n353), .C1(new_n348), .C2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT38), .ZN(new_n356));
  XNOR2_X1  g155(.A(G8gat), .B(G36gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n357), .B(KEYINPUT75), .ZN(new_n358));
  XNOR2_X1  g157(.A(G64gat), .B(G92gat), .ZN(new_n359));
  XOR2_X1   g158(.A(new_n358), .B(new_n359), .Z(new_n360));
  NAND4_X1  g159(.A1(new_n351), .A2(new_n355), .A3(new_n356), .A4(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n360), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n352), .B(new_n362), .C1(new_n348), .C2(new_n354), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n280), .A2(new_n281), .A3(new_n361), .A4(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n278), .A2(new_n279), .A3(new_n363), .ZN(new_n365));
  AND4_X1   g164(.A1(new_n356), .A2(new_n355), .A3(new_n351), .A4(new_n360), .ZN(new_n366));
  OAI21_X1  g165(.A(KEYINPUT86), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n355), .A2(new_n360), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n307), .B1(new_n322), .B2(KEYINPUT65), .ZN(new_n369));
  AOI211_X1 g168(.A(KEYINPUT74), .B(new_n318), .C1(new_n369), .C2(new_n324), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n327), .B1(new_n326), .B2(new_n328), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n344), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n354), .B1(new_n372), .B2(new_n320), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n353), .B1(new_n374), .B2(new_n352), .ZN(new_n375));
  OAI21_X1  g174(.A(KEYINPUT38), .B1(new_n368), .B2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n364), .A2(new_n367), .A3(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n340), .A2(new_n344), .A3(new_n341), .ZN(new_n378));
  AOI21_X1  g177(.A(KEYINPUT3), .B1(new_n378), .B2(KEYINPUT82), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT82), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n340), .A2(new_n380), .A3(new_n344), .A4(new_n341), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n253), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n219), .A2(new_n344), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n342), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  OAI211_X1 g184(.A(G228gat), .B(G233gat), .C1(new_n382), .C2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(G228gat), .A2(G233gat), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n215), .B1(new_n338), .B2(KEYINPUT29), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(new_n252), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n384), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n386), .A2(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(KEYINPUT31), .B(G50gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(G78gat), .B(G106gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n394), .B(G22gat), .ZN(new_n395));
  INV_X1    g194(.A(new_n392), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n379), .A2(new_n381), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n385), .B1(new_n397), .B2(new_n252), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n390), .B(new_n396), .C1(new_n398), .C2(new_n387), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n393), .A2(new_n395), .A3(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n395), .ZN(new_n401));
  INV_X1    g200(.A(new_n399), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n396), .B1(new_n386), .B2(new_n390), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n401), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  AND2_X1   g203(.A1(new_n400), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT30), .ZN(new_n406));
  AND2_X1   g205(.A1(new_n363), .A2(new_n406), .ZN(new_n407));
  AND3_X1   g206(.A1(new_n330), .A2(new_n345), .A3(new_n342), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n360), .B1(new_n408), .B2(new_n373), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n360), .A2(new_n406), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n352), .B(new_n410), .C1(new_n348), .C2(new_n354), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  OAI21_X1  g211(.A(KEYINPUT83), .B1(new_n407), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n363), .A2(new_n406), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT83), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n414), .A2(new_n415), .A3(new_n411), .A4(new_n409), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n257), .B1(new_n236), .B2(new_n247), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n262), .A2(new_n263), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT84), .B1(new_n418), .B2(new_n256), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT84), .ZN(new_n420));
  AOI211_X1 g219(.A(new_n420), .B(new_n257), .C1(new_n262), .C2(new_n263), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n417), .B(KEYINPUT39), .C1(new_n419), .C2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n417), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT39), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n276), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n422), .A2(new_n425), .A3(KEYINPUT40), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n426), .A2(new_n270), .A3(new_n277), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT40), .B1(new_n422), .B2(new_n425), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n413), .A2(new_n416), .A3(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n377), .A2(new_n405), .A3(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT36), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n235), .B1(new_n308), .B2(new_n318), .ZN(new_n433));
  AND2_X1   g232(.A1(G227gat), .A2(G233gat), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n326), .A2(new_n250), .A3(new_n328), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT32), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT33), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  XNOR2_X1  g238(.A(G15gat), .B(G43gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(G71gat), .B(G99gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n440), .B(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n437), .A2(new_n439), .A3(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT34), .ZN(new_n445));
  OR2_X1    g244(.A1(new_n442), .A2(KEYINPUT71), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n442), .A2(KEYINPUT71), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n446), .A2(KEYINPUT33), .A3(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n436), .A2(KEYINPUT32), .A3(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n444), .A2(new_n445), .A3(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n445), .B1(new_n444), .B2(new_n449), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n434), .B1(new_n433), .B2(new_n435), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n453), .A2(KEYINPUT72), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  NOR3_X1   g254(.A1(new_n451), .A2(new_n452), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n444), .A2(new_n449), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT34), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n454), .B1(new_n458), .B2(new_n450), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n432), .B1(new_n456), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n400), .A2(new_n404), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n274), .A2(new_n276), .A3(new_n275), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n273), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(new_n279), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n464), .A2(new_n414), .A3(new_n411), .A4(new_n409), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n455), .B1(new_n451), .B2(new_n452), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n458), .A2(new_n454), .A3(new_n450), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n467), .A2(new_n468), .A3(KEYINPUT36), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n460), .A2(new_n466), .A3(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n431), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n464), .ZN(new_n473));
  NOR3_X1   g272(.A1(new_n473), .A2(new_n407), .A3(new_n412), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n467), .A2(new_n468), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n474), .A2(new_n405), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT35), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n461), .B1(new_n468), .B2(new_n467), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n278), .A2(new_n279), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT35), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n481), .B1(new_n413), .B2(new_n416), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n478), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n477), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n472), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(G134gat), .B(G162gat), .ZN(new_n486));
  XOR2_X1   g285(.A(KEYINPUT87), .B(G29gat), .Z(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(G36gat), .ZN(new_n488));
  NOR2_X1   g287(.A1(G29gat), .A2(G36gat), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT14), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n489), .B(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n488), .A2(KEYINPUT88), .A3(new_n491), .ZN(new_n492));
  AND2_X1   g291(.A1(G43gat), .A2(G50gat), .ZN(new_n493));
  NOR2_X1   g292(.A1(G43gat), .A2(G50gat), .ZN(new_n494));
  OAI21_X1  g293(.A(KEYINPUT15), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  XOR2_X1   g294(.A(new_n492), .B(new_n495), .Z(new_n496));
  INV_X1    g295(.A(KEYINPUT15), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n493), .B1(KEYINPUT89), .B2(new_n497), .ZN(new_n498));
  OR2_X1    g297(.A1(new_n497), .A2(KEYINPUT89), .ZN(new_n499));
  AND2_X1   g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  XOR2_X1   g299(.A(KEYINPUT90), .B(G50gat), .Z(new_n501));
  INV_X1    g300(.A(G43gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n500), .A2(new_n488), .A3(new_n491), .A4(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n496), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT17), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n505), .B(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT95), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT7), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(KEYINPUT95), .A2(KEYINPUT7), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n510), .A2(G85gat), .A3(G92gat), .A4(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(G85gat), .ZN(new_n513));
  INV_X1    g312(.A(G92gat), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n508), .B(new_n509), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(G99gat), .A2(G106gat), .ZN(new_n516));
  AOI22_X1  g315(.A1(KEYINPUT8), .A2(new_n516), .B1(new_n513), .B2(new_n514), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n512), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  OR2_X1    g317(.A1(G99gat), .A2(G106gat), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n518), .A2(new_n516), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n516), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n512), .A2(new_n521), .A3(new_n515), .A4(new_n517), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n507), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT96), .ZN(new_n526));
  AND2_X1   g325(.A1(new_n496), .A2(new_n504), .ZN(new_n527));
  AND2_X1   g326(.A1(G232gat), .A2(G233gat), .ZN(new_n528));
  AOI22_X1  g327(.A1(new_n527), .A2(new_n523), .B1(KEYINPUT41), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n525), .A2(new_n526), .A3(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n526), .B1(new_n525), .B2(new_n529), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n486), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n532), .ZN(new_n534));
  INV_X1    g333(.A(new_n486), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n534), .A2(new_n530), .A3(new_n535), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n528), .A2(KEYINPUT41), .ZN(new_n537));
  XNOR2_X1  g336(.A(G190gat), .B(G218gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n537), .B(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n533), .A2(new_n536), .A3(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n539), .B1(new_n533), .B2(new_n536), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(G15gat), .B(G22gat), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n544), .A2(G1gat), .ZN(new_n545));
  INV_X1    g344(.A(G1gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT16), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n545), .B1(new_n544), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(KEYINPUT91), .ZN(new_n549));
  INV_X1    g348(.A(G8gat), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT91), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n550), .B1(new_n545), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT92), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n548), .A2(new_n550), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT21), .ZN(new_n559));
  XNOR2_X1  g358(.A(G57gat), .B(G64gat), .ZN(new_n560));
  AOI21_X1  g359(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n561));
  OR2_X1    g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  XOR2_X1   g361(.A(G71gat), .B(G78gat), .Z(new_n563));
  OR2_X1    g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n563), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n558), .B1(new_n559), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n559), .ZN(new_n568));
  NAND2_X1  g367(.A1(G231gat), .A2(G233gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(G127gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n567), .B(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(G155gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(G183gat), .B(G211gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n572), .B(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n543), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G120gat), .B(G148gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(G176gat), .B(G204gat), .ZN(new_n581));
  XOR2_X1   g380(.A(new_n580), .B(new_n581), .Z(new_n582));
  XNOR2_X1  g381(.A(new_n523), .B(new_n566), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT10), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(KEYINPUT97), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n523), .A2(KEYINPUT10), .A3(new_n565), .A4(new_n564), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT97), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n583), .A2(new_n588), .A3(new_n584), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n586), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(G230gat), .A2(G233gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT98), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n590), .A2(KEYINPUT98), .A3(new_n591), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OR2_X1    g395(.A1(new_n583), .A2(new_n591), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n582), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  AND3_X1   g397(.A1(new_n592), .A2(new_n597), .A3(new_n582), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n579), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(G229gat), .A2(G233gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(KEYINPUT93), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n557), .A2(new_n527), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n505), .B(KEYINPUT17), .ZN(new_n607));
  OAI211_X1 g406(.A(new_n605), .B(new_n606), .C1(new_n607), .C2(new_n557), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT18), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n507), .A2(new_n558), .ZN(new_n611));
  NAND4_X1  g410(.A1(new_n611), .A2(KEYINPUT18), .A3(new_n605), .A4(new_n606), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n604), .B(KEYINPUT13), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n555), .A2(new_n505), .A3(new_n556), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n614), .B1(new_n606), .B2(new_n615), .ZN(new_n616));
  AND2_X1   g415(.A1(new_n616), .A2(KEYINPUT94), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n616), .A2(KEYINPUT94), .ZN(new_n618));
  OAI211_X1 g417(.A(new_n610), .B(new_n612), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(G113gat), .B(G141gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(G197gat), .ZN(new_n621));
  XOR2_X1   g420(.A(KEYINPUT11), .B(G169gat), .Z(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XOR2_X1   g422(.A(new_n623), .B(KEYINPUT12), .Z(new_n624));
  NAND2_X1  g423(.A1(new_n619), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n616), .B(KEYINPUT94), .ZN(new_n626));
  INV_X1    g425(.A(new_n624), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n626), .A2(new_n627), .A3(new_n612), .A4(new_n610), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n485), .A2(new_n602), .A3(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT99), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n629), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n633), .B1(new_n472), .B2(new_n484), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n634), .A2(KEYINPUT99), .A3(new_n602), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(new_n473), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g437(.A1(new_n413), .A2(new_n416), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n639), .B1(new_n632), .B2(new_n635), .ZN(new_n640));
  XOR2_X1   g439(.A(KEYINPUT16), .B(G8gat), .Z(new_n641));
  NAND3_X1  g440(.A1(new_n640), .A2(KEYINPUT42), .A3(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n639), .ZN(new_n643));
  INV_X1    g442(.A(new_n635), .ZN(new_n644));
  AOI21_X1  g443(.A(KEYINPUT99), .B1(new_n634), .B2(new_n602), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n643), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(KEYINPUT101), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT101), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n640), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n647), .A2(G8gat), .A3(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n641), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n651), .B1(new_n647), .B2(new_n649), .ZN(new_n652));
  XNOR2_X1  g451(.A(KEYINPUT100), .B(KEYINPUT42), .ZN(new_n653));
  OAI211_X1 g452(.A(new_n642), .B(new_n650), .C1(new_n652), .C2(new_n653), .ZN(G1325gat));
  INV_X1    g453(.A(G15gat), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n636), .A2(new_n655), .A3(new_n475), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n460), .A2(new_n469), .ZN(new_n657));
  OR2_X1    g456(.A1(new_n657), .A2(KEYINPUT102), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(KEYINPUT102), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n660), .B1(new_n632), .B2(new_n635), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n656), .B1(new_n661), .B2(new_n655), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT103), .ZN(G1326gat));
  NAND2_X1  g462(.A1(new_n636), .A2(new_n461), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(KEYINPUT104), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT104), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n636), .A2(new_n666), .A3(new_n461), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(KEYINPUT43), .B(G22gat), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n665), .A2(new_n667), .A3(new_n669), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(G1327gat));
  AND2_X1   g472(.A1(new_n430), .A2(new_n405), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n470), .B1(new_n377), .B2(new_n674), .ZN(new_n675));
  AOI22_X1  g474(.A1(new_n476), .A2(KEYINPUT35), .B1(new_n478), .B2(new_n482), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n543), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n678), .A2(new_n577), .A3(new_n600), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n677), .A2(new_n633), .A3(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n487), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n680), .A2(new_n473), .A3(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT45), .ZN(new_n683));
  OR2_X1    g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n685), .B1(new_n677), .B2(new_n543), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n485), .A2(KEYINPUT44), .A3(new_n678), .ZN(new_n687));
  AND3_X1   g486(.A1(new_n625), .A2(KEYINPUT105), .A3(new_n628), .ZN(new_n688));
  AOI21_X1  g487(.A(KEYINPUT105), .B1(new_n625), .B2(new_n628), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n690), .A2(new_n578), .A3(new_n601), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n686), .A2(new_n687), .A3(new_n473), .A4(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(new_n487), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n682), .A2(new_n683), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n684), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(KEYINPUT106), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT106), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n684), .A2(new_n697), .A3(new_n693), .A4(new_n694), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(new_n698), .ZN(G1328gat));
  INV_X1    g498(.A(KEYINPUT107), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n639), .A2(G36gat), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n680), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT46), .ZN(new_n703));
  INV_X1    g502(.A(new_n679), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n634), .A2(new_n704), .A3(new_n701), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(KEYINPUT107), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n702), .A2(new_n703), .A3(new_n706), .ZN(new_n707));
  XOR2_X1   g506(.A(new_n707), .B(KEYINPUT108), .Z(new_n708));
  AOI21_X1  g507(.A(new_n703), .B1(new_n702), .B2(new_n706), .ZN(new_n709));
  AND2_X1   g508(.A1(new_n686), .A2(new_n687), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n710), .A2(new_n643), .A3(new_n691), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n709), .B1(G36gat), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n708), .A2(new_n712), .ZN(G1329gat));
  NAND3_X1  g512(.A1(new_n680), .A2(new_n502), .A3(new_n475), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n686), .A2(new_n687), .A3(new_n657), .A4(new_n691), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(KEYINPUT109), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(G43gat), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n715), .A2(KEYINPUT109), .ZN(new_n718));
  OAI211_X1 g517(.A(KEYINPUT47), .B(new_n714), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n660), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n686), .A2(new_n720), .A3(new_n687), .A4(new_n691), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(G43gat), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n722), .A2(new_n714), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n719), .B1(KEYINPUT47), .B2(new_n723), .ZN(G1330gat));
  NAND4_X1  g523(.A1(new_n686), .A2(new_n687), .A3(new_n461), .A4(new_n691), .ZN(new_n725));
  INV_X1    g524(.A(new_n501), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n680), .A2(new_n461), .A3(new_n501), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(KEYINPUT48), .B1(new_n728), .B2(KEYINPUT110), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n729), .B(new_n730), .ZN(G1331gat));
  NAND4_X1  g530(.A1(new_n690), .A2(new_n578), .A3(new_n543), .A4(new_n601), .ZN(new_n732));
  OR3_X1    g531(.A1(new_n677), .A2(KEYINPUT111), .A3(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(KEYINPUT111), .B1(new_n677), .B2(new_n732), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n735), .A2(new_n464), .ZN(new_n736));
  XOR2_X1   g535(.A(KEYINPUT112), .B(G57gat), .Z(new_n737));
  XNOR2_X1  g536(.A(new_n736), .B(new_n737), .ZN(G1332gat));
  OAI22_X1  g537(.A1(new_n735), .A2(new_n639), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n739));
  XNOR2_X1  g538(.A(KEYINPUT49), .B(G64gat), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n733), .A2(new_n643), .A3(new_n734), .A4(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n739), .A2(new_n741), .ZN(G1333gat));
  OAI21_X1  g541(.A(G71gat), .B1(new_n735), .B2(new_n660), .ZN(new_n743));
  INV_X1    g542(.A(G71gat), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n475), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n743), .B1(new_n735), .B2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT50), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  OAI211_X1 g547(.A(new_n743), .B(KEYINPUT50), .C1(new_n735), .C2(new_n745), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(G1334gat));
  NOR2_X1   g549(.A1(new_n735), .A2(new_n405), .ZN(new_n751));
  XNOR2_X1  g550(.A(KEYINPUT113), .B(G78gat), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n751), .B(new_n752), .ZN(G1335gat));
  INV_X1    g552(.A(KEYINPUT105), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n629), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n625), .A2(KEYINPUT105), .A3(new_n628), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n757), .A2(new_n578), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n759), .A2(new_n600), .ZN(new_n760));
  AND3_X1   g559(.A1(new_n710), .A2(new_n473), .A3(new_n760), .ZN(new_n761));
  OAI211_X1 g560(.A(new_n678), .B(new_n758), .C1(new_n675), .C2(new_n676), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(KEYINPUT51), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n601), .A2(new_n513), .A3(new_n473), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(KEYINPUT114), .ZN(new_n765));
  OAI22_X1  g564(.A1(new_n761), .A2(new_n513), .B1(new_n763), .B2(new_n765), .ZN(G1336gat));
  NAND4_X1  g565(.A1(new_n686), .A2(new_n687), .A3(new_n643), .A4(new_n760), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(G92gat), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT52), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n601), .A2(new_n643), .A3(new_n514), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(KEYINPUT115), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n768), .B(new_n769), .C1(new_n763), .C2(new_n771), .ZN(new_n772));
  XOR2_X1   g571(.A(KEYINPUT116), .B(KEYINPUT51), .Z(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n762), .A2(KEYINPUT117), .A3(new_n774), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n485), .A2(KEYINPUT51), .A3(new_n678), .A4(new_n758), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(KEYINPUT117), .B1(new_n762), .B2(new_n774), .ZN(new_n778));
  OR2_X1    g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(new_n771), .ZN(new_n780));
  AOI22_X1  g579(.A1(new_n779), .A2(new_n780), .B1(G92gat), .B2(new_n767), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n772), .B1(new_n781), .B2(new_n769), .ZN(G1337gat));
  NAND4_X1  g581(.A1(new_n686), .A2(new_n720), .A3(new_n687), .A4(new_n760), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(G99gat), .ZN(new_n784));
  INV_X1    g583(.A(G99gat), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n601), .A2(new_n785), .A3(new_n475), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(KEYINPUT118), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n784), .B1(new_n763), .B2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT119), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n788), .B(new_n789), .ZN(G1338gat));
  NAND4_X1  g589(.A1(new_n686), .A2(new_n687), .A3(new_n461), .A4(new_n760), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(G106gat), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT53), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n600), .A2(new_n405), .A3(G106gat), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n792), .B(new_n793), .C1(new_n763), .C2(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n794), .B1(new_n777), .B2(new_n778), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n792), .ZN(new_n798));
  AOI21_X1  g597(.A(KEYINPUT120), .B1(new_n798), .B2(KEYINPUT53), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT120), .ZN(new_n800));
  AOI211_X1 g599(.A(new_n800), .B(new_n793), .C1(new_n797), .C2(new_n792), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n796), .B1(new_n799), .B2(new_n801), .ZN(G1339gat));
  NOR3_X1   g601(.A1(new_n579), .A2(new_n757), .A3(new_n601), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT121), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT54), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n594), .A2(new_n806), .A3(new_n595), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n806), .B1(new_n590), .B2(new_n591), .ZN(new_n808));
  INV_X1    g607(.A(new_n591), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n586), .A2(new_n809), .A3(new_n587), .A4(new_n589), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n582), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n807), .A2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT55), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n805), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n599), .B1(new_n812), .B2(new_n813), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n807), .A2(new_n811), .A3(KEYINPUT121), .A4(KEYINPUT55), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n814), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n605), .B1(new_n611), .B2(new_n606), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n818), .A2(KEYINPUT122), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n606), .A2(new_n615), .A3(new_n614), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n820), .B1(new_n818), .B2(KEYINPUT122), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n623), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n628), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n817), .A2(new_n543), .A3(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(new_n823), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n601), .A2(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n826), .B1(new_n690), .B2(new_n817), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n824), .B1(new_n827), .B2(new_n543), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n804), .B1(new_n828), .B2(new_n578), .ZN(new_n829));
  INV_X1    g628(.A(new_n478), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n830), .A2(new_n464), .A3(new_n643), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(KEYINPUT123), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT123), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n829), .A2(new_n834), .A3(new_n831), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n833), .A2(new_n629), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(G113gat), .ZN(new_n837));
  AND3_X1   g636(.A1(new_n814), .A2(new_n815), .A3(new_n816), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n838), .A2(new_n678), .A3(new_n825), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n600), .A2(new_n823), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n840), .B1(new_n757), .B2(new_n838), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n839), .B1(new_n841), .B2(new_n678), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n803), .B1(new_n842), .B2(new_n577), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n843), .A2(new_n464), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n830), .A2(new_n643), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(new_n232), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n846), .A2(new_n847), .A3(new_n757), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n837), .A2(new_n848), .ZN(G1340gat));
  AOI21_X1  g648(.A(G120gat), .B1(new_n846), .B2(new_n601), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n833), .A2(new_n835), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n600), .A2(new_n227), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n850), .B1(new_n851), .B2(new_n852), .ZN(G1341gat));
  NAND3_X1  g652(.A1(new_n833), .A2(new_n578), .A3(new_n835), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(G127gat), .ZN(new_n855));
  INV_X1    g654(.A(G127gat), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n846), .A2(new_n856), .A3(new_n578), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n855), .A2(new_n857), .ZN(G1342gat));
  NAND3_X1  g657(.A1(new_n833), .A2(new_n678), .A3(new_n835), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(G134gat), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n543), .A2(G134gat), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n844), .A2(new_n845), .A3(new_n861), .ZN(new_n862));
  OR2_X1    g661(.A1(new_n862), .A2(KEYINPUT56), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(KEYINPUT56), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n860), .A2(new_n863), .A3(new_n864), .ZN(G1343gat));
  NOR3_X1   g664(.A1(new_n720), .A2(new_n405), .A3(new_n643), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n633), .A2(G141gat), .ZN(new_n867));
  AND3_X1   g666(.A1(new_n844), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n657), .A2(new_n464), .A3(new_n643), .ZN(new_n869));
  AOI21_X1  g668(.A(KEYINPUT57), .B1(new_n829), .B2(new_n461), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT57), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n405), .A2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n629), .A2(new_n814), .A3(new_n815), .A4(new_n816), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n678), .B1(new_n874), .B2(new_n826), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n577), .B1(new_n875), .B2(new_n824), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n873), .B1(new_n876), .B2(new_n804), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n757), .B(new_n869), .C1(new_n870), .C2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n868), .B1(new_n878), .B2(G141gat), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT58), .ZN(new_n880));
  INV_X1    g679(.A(new_n869), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n871), .B1(new_n843), .B2(new_n405), .ZN(new_n882));
  INV_X1    g681(.A(new_n877), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n207), .B1(new_n884), .B2(new_n629), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n844), .A2(new_n866), .ZN(new_n886));
  INV_X1    g685(.A(new_n867), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n880), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI22_X1  g687(.A1(new_n879), .A2(new_n880), .B1(new_n885), .B2(new_n888), .ZN(G1344gat));
  INV_X1    g688(.A(new_n204), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n600), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n844), .A2(new_n866), .A3(new_n891), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n892), .B(KEYINPUT124), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT125), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n601), .B1(new_n869), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n896), .B1(new_n895), .B2(new_n869), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n843), .A2(new_n873), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n602), .A2(new_n633), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n876), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(KEYINPUT57), .B1(new_n900), .B2(new_n461), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n897), .B1(new_n898), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n894), .B1(new_n902), .B2(G148gat), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n890), .A2(new_n894), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n904), .B1(new_n884), .B2(new_n601), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n893), .B1(new_n903), .B2(new_n905), .ZN(G1345gat));
  OAI21_X1  g705(.A(new_n869), .B1(new_n870), .B2(new_n877), .ZN(new_n907));
  OAI21_X1  g706(.A(G155gat), .B1(new_n907), .B2(new_n577), .ZN(new_n908));
  OR2_X1    g707(.A1(new_n577), .A2(G155gat), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n908), .B1(new_n886), .B2(new_n909), .ZN(G1346gat));
  NOR2_X1   g709(.A1(new_n907), .A2(new_n543), .ZN(new_n911));
  XNOR2_X1  g710(.A(KEYINPUT78), .B(G162gat), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n678), .A2(new_n912), .ZN(new_n913));
  OAI22_X1  g712(.A1(new_n911), .A2(new_n912), .B1(new_n886), .B2(new_n913), .ZN(G1347gat));
  NOR2_X1   g713(.A1(new_n639), .A2(new_n473), .ZN(new_n915));
  INV_X1    g714(.A(new_n915), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n916), .A2(new_n830), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n829), .A2(new_n917), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n918), .A2(new_n292), .A3(new_n633), .ZN(new_n919));
  INV_X1    g718(.A(new_n918), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(new_n757), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n919), .B1(new_n292), .B2(new_n921), .ZN(G1348gat));
  NOR2_X1   g721(.A1(new_n918), .A2(new_n600), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n923), .B(new_n293), .ZN(G1349gat));
  OR3_X1    g723(.A1(new_n918), .A2(new_n313), .A3(new_n577), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT60), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n288), .B1(new_n918), .B2(new_n577), .ZN(new_n927));
  AND3_X1   g726(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n926), .B1(new_n925), .B2(new_n927), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n928), .A2(new_n929), .ZN(G1350gat));
  OAI22_X1  g729(.A1(new_n918), .A2(new_n543), .B1(KEYINPUT61), .B2(G190gat), .ZN(new_n931));
  NAND2_X1  g730(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n931), .B(new_n932), .ZN(G1351gat));
  NAND2_X1  g732(.A1(new_n660), .A2(new_n915), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n843), .A2(new_n405), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(G197gat), .B1(new_n935), .B2(new_n757), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n900), .A2(new_n461), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(new_n871), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n829), .A2(new_n872), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n934), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n629), .A2(G197gat), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n936), .B1(new_n940), .B2(new_n941), .ZN(G1352gat));
  INV_X1    g741(.A(G204gat), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n935), .A2(new_n943), .A3(new_n601), .ZN(new_n944));
  OR2_X1    g743(.A1(new_n944), .A2(KEYINPUT62), .ZN(new_n945));
  INV_X1    g744(.A(new_n934), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n946), .B1(new_n898), .B2(new_n901), .ZN(new_n947));
  OAI21_X1  g746(.A(G204gat), .B1(new_n947), .B2(new_n600), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n944), .A2(KEYINPUT62), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n945), .A2(new_n948), .A3(new_n949), .ZN(G1353gat));
  NAND3_X1  g749(.A1(new_n935), .A2(new_n333), .A3(new_n578), .ZN(new_n951));
  OAI211_X1 g750(.A(new_n578), .B(new_n946), .C1(new_n898), .C2(new_n901), .ZN(new_n952));
  AND3_X1   g751(.A1(new_n952), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n953));
  AOI21_X1  g752(.A(KEYINPUT63), .B1(new_n952), .B2(G211gat), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n951), .B1(new_n953), .B2(new_n954), .ZN(G1354gat));
  OR2_X1    g754(.A1(new_n940), .A2(KEYINPUT127), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n678), .A2(G218gat), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n957), .B1(new_n940), .B2(KEYINPUT127), .ZN(new_n958));
  NAND4_X1  g757(.A1(new_n829), .A2(new_n461), .A3(new_n678), .A4(new_n946), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(new_n334), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT126), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n959), .A2(KEYINPUT126), .A3(new_n334), .ZN(new_n963));
  AOI22_X1  g762(.A1(new_n956), .A2(new_n958), .B1(new_n962), .B2(new_n963), .ZN(G1355gat));
endmodule


