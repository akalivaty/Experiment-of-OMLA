

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584;

  XNOR2_X1 U321 ( .A(n348), .B(KEYINPUT111), .ZN(n349) );
  XNOR2_X1 U322 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n404) );
  XNOR2_X1 U323 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U324 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U325 ( .A(KEYINPUT9), .B(KEYINPUT80), .Z(n289) );
  NOR2_X1 U326 ( .A1(n575), .A2(n398), .ZN(n399) );
  XNOR2_X1 U327 ( .A(n350), .B(n349), .ZN(n393) );
  XNOR2_X1 U328 ( .A(KEYINPUT122), .B(KEYINPUT54), .ZN(n419) );
  OR2_X1 U329 ( .A1(n301), .A2(n302), .ZN(n304) );
  INV_X1 U330 ( .A(KEYINPUT78), .ZN(n308) );
  NOR2_X1 U331 ( .A1(n475), .A2(n568), .ZN(n440) );
  XNOR2_X1 U332 ( .A(KEYINPUT105), .B(KEYINPUT36), .ZN(n396) );
  XNOR2_X1 U333 ( .A(n558), .B(n396), .ZN(n582) );
  XOR2_X1 U334 ( .A(n457), .B(KEYINPUT124), .Z(n565) );
  XOR2_X1 U335 ( .A(n475), .B(KEYINPUT28), .Z(n534) );
  XNOR2_X1 U336 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U337 ( .A(n464), .B(n463), .ZN(G1351GAT) );
  XNOR2_X1 U338 ( .A(G106GAT), .B(G78GAT), .ZN(n290) );
  XNOR2_X1 U339 ( .A(n290), .B(G148GAT), .ZN(n320) );
  XOR2_X1 U340 ( .A(G64GAT), .B(G92GAT), .Z(n292) );
  XNOR2_X1 U341 ( .A(G176GAT), .B(G204GAT), .ZN(n291) );
  XNOR2_X1 U342 ( .A(n292), .B(n291), .ZN(n409) );
  XNOR2_X1 U343 ( .A(n320), .B(n409), .ZN(n313) );
  XOR2_X1 U344 ( .A(KEYINPUT74), .B(KEYINPUT73), .Z(n298) );
  XOR2_X1 U345 ( .A(G120GAT), .B(G71GAT), .Z(n442) );
  INV_X1 U346 ( .A(KEYINPUT13), .ZN(n293) );
  NAND2_X1 U347 ( .A1(G57GAT), .A2(n293), .ZN(n296) );
  INV_X1 U348 ( .A(G57GAT), .ZN(n294) );
  NAND2_X1 U349 ( .A1(n294), .A2(KEYINPUT13), .ZN(n295) );
  NAND2_X1 U350 ( .A1(n296), .A2(n295), .ZN(n382) );
  XNOR2_X1 U351 ( .A(n442), .B(n382), .ZN(n297) );
  XNOR2_X1 U352 ( .A(n298), .B(n297), .ZN(n301) );
  XOR2_X1 U353 ( .A(KEYINPUT77), .B(KEYINPUT31), .Z(n300) );
  XNOR2_X1 U354 ( .A(KEYINPUT32), .B(KEYINPUT76), .ZN(n299) );
  XNOR2_X1 U355 ( .A(n300), .B(n299), .ZN(n302) );
  NAND2_X1 U356 ( .A1(n302), .A2(n301), .ZN(n303) );
  NAND2_X1 U357 ( .A1(n304), .A2(n303), .ZN(n306) );
  AND2_X1 U358 ( .A1(G230GAT), .A2(G233GAT), .ZN(n305) );
  XNOR2_X1 U359 ( .A(n306), .B(n305), .ZN(n311) );
  XNOR2_X1 U360 ( .A(G99GAT), .B(G85GAT), .ZN(n307) );
  XNOR2_X1 U361 ( .A(n307), .B(KEYINPUT75), .ZN(n365) );
  XNOR2_X1 U362 ( .A(n365), .B(KEYINPUT33), .ZN(n309) );
  XNOR2_X1 U363 ( .A(n313), .B(n312), .ZN(n575) );
  XNOR2_X1 U364 ( .A(KEYINPUT41), .B(n575), .ZN(n550) );
  XOR2_X1 U365 ( .A(n550), .B(KEYINPUT108), .Z(n538) );
  XOR2_X1 U366 ( .A(KEYINPUT95), .B(G218GAT), .Z(n315) );
  XNOR2_X1 U367 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n314) );
  XNOR2_X1 U368 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U369 ( .A(G197GAT), .B(n316), .Z(n415) );
  XOR2_X1 U370 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n318) );
  XNOR2_X1 U371 ( .A(KEYINPUT94), .B(G204GAT), .ZN(n317) );
  XNOR2_X1 U372 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U373 ( .A(n415), .B(n319), .ZN(n330) );
  XOR2_X1 U374 ( .A(KEYINPUT22), .B(n320), .Z(n322) );
  NAND2_X1 U375 ( .A1(G228GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U376 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U377 ( .A(n323), .B(KEYINPUT93), .Z(n328) );
  XNOR2_X1 U378 ( .A(G50GAT), .B(G22GAT), .ZN(n324) );
  XNOR2_X1 U379 ( .A(n324), .B(G141GAT), .ZN(n345) );
  XOR2_X1 U380 ( .A(G155GAT), .B(KEYINPUT3), .Z(n326) );
  XNOR2_X1 U381 ( .A(G162GAT), .B(KEYINPUT2), .ZN(n325) );
  XNOR2_X1 U382 ( .A(n326), .B(n325), .ZN(n425) );
  XNOR2_X1 U383 ( .A(n345), .B(n425), .ZN(n327) );
  XNOR2_X1 U384 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U385 ( .A(n330), .B(n329), .ZN(n475) );
  XOR2_X1 U386 ( .A(KEYINPUT67), .B(KEYINPUT29), .Z(n332) );
  XNOR2_X1 U387 ( .A(KEYINPUT66), .B(KEYINPUT68), .ZN(n331) );
  XNOR2_X1 U388 ( .A(n332), .B(n331), .ZN(n336) );
  XOR2_X1 U389 ( .A(KEYINPUT71), .B(G197GAT), .Z(n334) );
  XOR2_X1 U390 ( .A(G113GAT), .B(G1GAT), .Z(n422) );
  XOR2_X1 U391 ( .A(G15GAT), .B(KEYINPUT70), .Z(n383) );
  XNOR2_X1 U392 ( .A(n422), .B(n383), .ZN(n333) );
  XNOR2_X1 U393 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U394 ( .A(n336), .B(n335), .Z(n338) );
  NAND2_X1 U395 ( .A1(G229GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U396 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U397 ( .A(n339), .B(KEYINPUT69), .Z(n343) );
  XOR2_X1 U398 ( .A(G29GAT), .B(G43GAT), .Z(n341) );
  XNOR2_X1 U399 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n340) );
  XNOR2_X1 U400 ( .A(n341), .B(n340), .ZN(n366) );
  XNOR2_X1 U401 ( .A(n366), .B(KEYINPUT30), .ZN(n342) );
  XNOR2_X1 U402 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U403 ( .A(n345), .B(n344), .ZN(n347) );
  XOR2_X1 U404 ( .A(G169GAT), .B(G36GAT), .Z(n346) );
  XOR2_X1 U405 ( .A(G8GAT), .B(n346), .Z(n406) );
  XNOR2_X1 U406 ( .A(n347), .B(n406), .ZN(n395) );
  NOR2_X1 U407 ( .A1(n395), .A2(n550), .ZN(n350) );
  XNOR2_X1 U408 ( .A(KEYINPUT46), .B(KEYINPUT112), .ZN(n348) );
  XOR2_X1 U409 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n352) );
  XNOR2_X1 U410 ( .A(G218GAT), .B(G92GAT), .ZN(n351) );
  XNOR2_X1 U411 ( .A(n352), .B(n351), .ZN(n355) );
  XNOR2_X1 U412 ( .A(G162GAT), .B(G106GAT), .ZN(n353) );
  XNOR2_X1 U413 ( .A(n289), .B(n353), .ZN(n354) );
  XOR2_X1 U414 ( .A(n355), .B(n354), .Z(n360) );
  XOR2_X1 U415 ( .A(KEYINPUT81), .B(KEYINPUT82), .Z(n357) );
  NAND2_X1 U416 ( .A1(G232GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U417 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U418 ( .A(KEYINPUT65), .B(n358), .ZN(n359) );
  XNOR2_X1 U419 ( .A(n360), .B(n359), .ZN(n364) );
  XOR2_X1 U420 ( .A(G134GAT), .B(G190GAT), .Z(n362) );
  XNOR2_X1 U421 ( .A(G50GAT), .B(G36GAT), .ZN(n361) );
  XNOR2_X1 U422 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U423 ( .A(n364), .B(n363), .ZN(n368) );
  XOR2_X1 U424 ( .A(n366), .B(n365), .Z(n367) );
  XNOR2_X1 U425 ( .A(n368), .B(n367), .ZN(n558) );
  XOR2_X1 U426 ( .A(KEYINPUT85), .B(KEYINPUT15), .Z(n370) );
  XNOR2_X1 U427 ( .A(KEYINPUT12), .B(KEYINPUT83), .ZN(n369) );
  XNOR2_X1 U428 ( .A(n370), .B(n369), .ZN(n391) );
  XOR2_X1 U429 ( .A(G71GAT), .B(G127GAT), .Z(n372) );
  XNOR2_X1 U430 ( .A(G1GAT), .B(G183GAT), .ZN(n371) );
  XNOR2_X1 U431 ( .A(n372), .B(n371), .ZN(n376) );
  XOR2_X1 U432 ( .A(KEYINPUT14), .B(KEYINPUT86), .Z(n374) );
  XNOR2_X1 U433 ( .A(G8GAT), .B(G64GAT), .ZN(n373) );
  XNOR2_X1 U434 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U435 ( .A(n376), .B(n375), .Z(n381) );
  XOR2_X1 U436 ( .A(KEYINPUT87), .B(KEYINPUT88), .Z(n378) );
  NAND2_X1 U437 ( .A1(G231GAT), .A2(G233GAT), .ZN(n377) );
  XNOR2_X1 U438 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U439 ( .A(KEYINPUT84), .B(n379), .ZN(n380) );
  XNOR2_X1 U440 ( .A(n381), .B(n380), .ZN(n387) );
  XOR2_X1 U441 ( .A(n382), .B(G78GAT), .Z(n385) );
  XNOR2_X1 U442 ( .A(n383), .B(G155GAT), .ZN(n384) );
  XNOR2_X1 U443 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U444 ( .A(n387), .B(n386), .Z(n389) );
  XNOR2_X1 U445 ( .A(G22GAT), .B(G211GAT), .ZN(n388) );
  XNOR2_X1 U446 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U447 ( .A(n391), .B(n390), .ZN(n556) );
  INV_X1 U448 ( .A(n556), .ZN(n578) );
  NOR2_X1 U449 ( .A1(n558), .A2(n578), .ZN(n392) );
  AND2_X1 U450 ( .A1(n393), .A2(n392), .ZN(n394) );
  XOR2_X1 U451 ( .A(n394), .B(KEYINPUT47), .Z(n403) );
  INV_X1 U452 ( .A(n395), .ZN(n571) );
  XNOR2_X1 U453 ( .A(KEYINPUT72), .B(n571), .ZN(n563) );
  NOR2_X1 U454 ( .A1(n582), .A2(n556), .ZN(n397) );
  XOR2_X1 U455 ( .A(KEYINPUT45), .B(n397), .Z(n398) );
  XNOR2_X1 U456 ( .A(n399), .B(KEYINPUT113), .ZN(n400) );
  NOR2_X1 U457 ( .A1(n563), .A2(n400), .ZN(n401) );
  XNOR2_X1 U458 ( .A(KEYINPUT114), .B(n401), .ZN(n402) );
  NOR2_X1 U459 ( .A1(n403), .A2(n402), .ZN(n405) );
  XNOR2_X1 U460 ( .A(n405), .B(n404), .ZN(n529) );
  XOR2_X1 U461 ( .A(KEYINPUT97), .B(n406), .Z(n408) );
  NAND2_X1 U462 ( .A1(G226GAT), .A2(G233GAT), .ZN(n407) );
  XNOR2_X1 U463 ( .A(n408), .B(n407), .ZN(n410) );
  XOR2_X1 U464 ( .A(n410), .B(n409), .Z(n417) );
  XNOR2_X1 U465 ( .A(KEYINPUT17), .B(KEYINPUT19), .ZN(n411) );
  XNOR2_X1 U466 ( .A(n411), .B(KEYINPUT18), .ZN(n412) );
  XOR2_X1 U467 ( .A(n412), .B(KEYINPUT90), .Z(n414) );
  XNOR2_X1 U468 ( .A(G183GAT), .B(G190GAT), .ZN(n413) );
  XNOR2_X1 U469 ( .A(n414), .B(n413), .ZN(n455) );
  XNOR2_X1 U470 ( .A(n455), .B(n415), .ZN(n416) );
  XOR2_X1 U471 ( .A(n417), .B(n416), .Z(n523) );
  XOR2_X1 U472 ( .A(n523), .B(KEYINPUT121), .Z(n418) );
  NOR2_X1 U473 ( .A1(n529), .A2(n418), .ZN(n420) );
  XNOR2_X1 U474 ( .A(n420), .B(n419), .ZN(n438) );
  XNOR2_X1 U475 ( .A(G134GAT), .B(G127GAT), .ZN(n421) );
  XNOR2_X1 U476 ( .A(n421), .B(KEYINPUT0), .ZN(n441) );
  XOR2_X1 U477 ( .A(G85GAT), .B(n441), .Z(n424) );
  XNOR2_X1 U478 ( .A(G29GAT), .B(n422), .ZN(n423) );
  XNOR2_X1 U479 ( .A(n424), .B(n423), .ZN(n429) );
  XOR2_X1 U480 ( .A(n425), .B(KEYINPUT4), .Z(n427) );
  NAND2_X1 U481 ( .A1(G225GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U482 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U483 ( .A(n429), .B(n428), .Z(n437) );
  XOR2_X1 U484 ( .A(KEYINPUT1), .B(G148GAT), .Z(n431) );
  XNOR2_X1 U485 ( .A(G141GAT), .B(G120GAT), .ZN(n430) );
  XNOR2_X1 U486 ( .A(n431), .B(n430), .ZN(n435) );
  XOR2_X1 U487 ( .A(KEYINPUT96), .B(G57GAT), .Z(n433) );
  XNOR2_X1 U488 ( .A(KEYINPUT6), .B(KEYINPUT5), .ZN(n432) );
  XNOR2_X1 U489 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U490 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U491 ( .A(n437), .B(n436), .ZN(n530) );
  NAND2_X1 U492 ( .A1(n438), .A2(n530), .ZN(n568) );
  XNOR2_X1 U493 ( .A(KEYINPUT55), .B(KEYINPUT123), .ZN(n439) );
  XNOR2_X1 U494 ( .A(n440), .B(n439), .ZN(n456) );
  XOR2_X1 U495 ( .A(n442), .B(n441), .Z(n444) );
  XNOR2_X1 U496 ( .A(G43GAT), .B(G99GAT), .ZN(n443) );
  XNOR2_X1 U497 ( .A(n444), .B(n443), .ZN(n448) );
  XOR2_X1 U498 ( .A(G15GAT), .B(G176GAT), .Z(n446) );
  NAND2_X1 U499 ( .A1(G227GAT), .A2(G233GAT), .ZN(n445) );
  XNOR2_X1 U500 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U501 ( .A(n448), .B(n447), .Z(n453) );
  XOR2_X1 U502 ( .A(KEYINPUT92), .B(KEYINPUT20), .Z(n450) );
  XNOR2_X1 U503 ( .A(G169GAT), .B(KEYINPUT91), .ZN(n449) );
  XNOR2_X1 U504 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U505 ( .A(G113GAT), .B(n451), .ZN(n452) );
  XNOR2_X1 U506 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U507 ( .A(n455), .B(n454), .ZN(n476) );
  NAND2_X1 U508 ( .A1(n456), .A2(n476), .ZN(n457) );
  NAND2_X1 U509 ( .A1(n538), .A2(n565), .ZN(n460) );
  XOR2_X1 U510 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n458) );
  XNOR2_X1 U511 ( .A(n458), .B(G176GAT), .ZN(n459) );
  XNOR2_X1 U512 ( .A(n460), .B(n459), .ZN(G1349GAT) );
  NAND2_X1 U513 ( .A1(n558), .A2(n565), .ZN(n464) );
  XOR2_X1 U514 ( .A(KEYINPUT58), .B(KEYINPUT126), .Z(n462) );
  INV_X1 U515 ( .A(G190GAT), .ZN(n461) );
  INV_X1 U516 ( .A(n575), .ZN(n465) );
  NAND2_X1 U517 ( .A1(n465), .A2(n563), .ZN(n466) );
  XNOR2_X1 U518 ( .A(n466), .B(KEYINPUT79), .ZN(n498) );
  XOR2_X1 U519 ( .A(n523), .B(KEYINPUT98), .Z(n467) );
  XNOR2_X1 U520 ( .A(n467), .B(KEYINPUT27), .ZN(n532) );
  INV_X1 U521 ( .A(n476), .ZN(n536) );
  NAND2_X1 U522 ( .A1(n475), .A2(n536), .ZN(n468) );
  XOR2_X1 U523 ( .A(n468), .B(KEYINPUT26), .Z(n570) );
  NAND2_X1 U524 ( .A1(n532), .A2(n570), .ZN(n469) );
  NAND2_X1 U525 ( .A1(n530), .A2(n469), .ZN(n474) );
  NOR2_X1 U526 ( .A1(n536), .A2(n523), .ZN(n470) );
  NOR2_X1 U527 ( .A1(n475), .A2(n470), .ZN(n471) );
  XNOR2_X1 U528 ( .A(KEYINPUT99), .B(n471), .ZN(n472) );
  XNOR2_X1 U529 ( .A(KEYINPUT25), .B(n472), .ZN(n473) );
  NOR2_X1 U530 ( .A1(n474), .A2(n473), .ZN(n480) );
  NAND2_X1 U531 ( .A1(n532), .A2(n534), .ZN(n477) );
  NOR2_X1 U532 ( .A1(n477), .A2(n476), .ZN(n478) );
  NOR2_X1 U533 ( .A1(n530), .A2(n478), .ZN(n479) );
  NOR2_X1 U534 ( .A1(n480), .A2(n479), .ZN(n481) );
  XNOR2_X1 U535 ( .A(KEYINPUT100), .B(n481), .ZN(n496) );
  NOR2_X1 U536 ( .A1(n556), .A2(n558), .ZN(n482) );
  XNOR2_X1 U537 ( .A(n482), .B(KEYINPUT89), .ZN(n483) );
  XOR2_X1 U538 ( .A(KEYINPUT16), .B(n483), .Z(n484) );
  AND2_X1 U539 ( .A1(n496), .A2(n484), .ZN(n510) );
  NAND2_X1 U540 ( .A1(n498), .A2(n510), .ZN(n492) );
  NOR2_X1 U541 ( .A1(n530), .A2(n492), .ZN(n486) );
  XNOR2_X1 U542 ( .A(KEYINPUT34), .B(KEYINPUT101), .ZN(n485) );
  XNOR2_X1 U543 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U544 ( .A(G1GAT), .B(n487), .ZN(G1324GAT) );
  NOR2_X1 U545 ( .A1(n523), .A2(n492), .ZN(n488) );
  XOR2_X1 U546 ( .A(G8GAT), .B(n488), .Z(G1325GAT) );
  NOR2_X1 U547 ( .A1(n536), .A2(n492), .ZN(n490) );
  XNOR2_X1 U548 ( .A(KEYINPUT35), .B(KEYINPUT102), .ZN(n489) );
  XNOR2_X1 U549 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U550 ( .A(G15GAT), .B(n491), .ZN(G1326GAT) );
  NOR2_X1 U551 ( .A1(n534), .A2(n492), .ZN(n494) );
  XNOR2_X1 U552 ( .A(G22GAT), .B(KEYINPUT103), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n494), .B(n493), .ZN(G1327GAT) );
  NOR2_X1 U554 ( .A1(n578), .A2(n582), .ZN(n495) );
  NAND2_X1 U555 ( .A1(n496), .A2(n495), .ZN(n497) );
  XNOR2_X1 U556 ( .A(KEYINPUT37), .B(n497), .ZN(n521) );
  NAND2_X1 U557 ( .A1(n498), .A2(n521), .ZN(n499) );
  XNOR2_X1 U558 ( .A(n499), .B(KEYINPUT38), .ZN(n507) );
  NOR2_X1 U559 ( .A1(n530), .A2(n507), .ZN(n502) );
  XNOR2_X1 U560 ( .A(G29GAT), .B(KEYINPUT104), .ZN(n500) );
  XNOR2_X1 U561 ( .A(n500), .B(KEYINPUT39), .ZN(n501) );
  XNOR2_X1 U562 ( .A(n502), .B(n501), .ZN(G1328GAT) );
  NOR2_X1 U563 ( .A1(n507), .A2(n523), .ZN(n503) );
  XOR2_X1 U564 ( .A(G36GAT), .B(n503), .Z(G1329GAT) );
  XNOR2_X1 U565 ( .A(KEYINPUT106), .B(KEYINPUT40), .ZN(n505) );
  NOR2_X1 U566 ( .A1(n536), .A2(n507), .ZN(n504) );
  XNOR2_X1 U567 ( .A(n505), .B(n504), .ZN(n506) );
  XOR2_X1 U568 ( .A(G43GAT), .B(n506), .Z(G1330GAT) );
  XNOR2_X1 U569 ( .A(G50GAT), .B(KEYINPUT107), .ZN(n509) );
  NOR2_X1 U570 ( .A1(n534), .A2(n507), .ZN(n508) );
  XNOR2_X1 U571 ( .A(n509), .B(n508), .ZN(G1331GAT) );
  AND2_X1 U572 ( .A1(n538), .A2(n395), .ZN(n520) );
  NAND2_X1 U573 ( .A1(n520), .A2(n510), .ZN(n515) );
  NOR2_X1 U574 ( .A1(n530), .A2(n515), .ZN(n511) );
  XOR2_X1 U575 ( .A(G57GAT), .B(n511), .Z(n512) );
  XNOR2_X1 U576 ( .A(KEYINPUT42), .B(n512), .ZN(G1332GAT) );
  NOR2_X1 U577 ( .A1(n523), .A2(n515), .ZN(n513) );
  XOR2_X1 U578 ( .A(G64GAT), .B(n513), .Z(G1333GAT) );
  NOR2_X1 U579 ( .A1(n536), .A2(n515), .ZN(n514) );
  XOR2_X1 U580 ( .A(G71GAT), .B(n514), .Z(G1334GAT) );
  NOR2_X1 U581 ( .A1(n515), .A2(n534), .ZN(n519) );
  XOR2_X1 U582 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n517) );
  XNOR2_X1 U583 ( .A(G78GAT), .B(KEYINPUT110), .ZN(n516) );
  XNOR2_X1 U584 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(G1335GAT) );
  NAND2_X1 U586 ( .A1(n521), .A2(n520), .ZN(n526) );
  NOR2_X1 U587 ( .A1(n530), .A2(n526), .ZN(n522) );
  XOR2_X1 U588 ( .A(G85GAT), .B(n522), .Z(G1336GAT) );
  NOR2_X1 U589 ( .A1(n523), .A2(n526), .ZN(n524) );
  XOR2_X1 U590 ( .A(G92GAT), .B(n524), .Z(G1337GAT) );
  NOR2_X1 U591 ( .A1(n536), .A2(n526), .ZN(n525) );
  XOR2_X1 U592 ( .A(G99GAT), .B(n525), .Z(G1338GAT) );
  NOR2_X1 U593 ( .A1(n534), .A2(n526), .ZN(n527) );
  XOR2_X1 U594 ( .A(KEYINPUT44), .B(n527), .Z(n528) );
  XNOR2_X1 U595 ( .A(G106GAT), .B(n528), .ZN(G1339GAT) );
  NOR2_X1 U596 ( .A1(n530), .A2(n529), .ZN(n531) );
  NAND2_X1 U597 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U598 ( .A(KEYINPUT115), .B(n533), .ZN(n548) );
  NAND2_X1 U599 ( .A1(n548), .A2(n534), .ZN(n535) );
  NOR2_X1 U600 ( .A1(n536), .A2(n535), .ZN(n545) );
  NAND2_X1 U601 ( .A1(n545), .A2(n563), .ZN(n537) );
  XNOR2_X1 U602 ( .A(n537), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n540) );
  NAND2_X1 U604 ( .A1(n545), .A2(n538), .ZN(n539) );
  XNOR2_X1 U605 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U606 ( .A(G120GAT), .B(n541), .ZN(G1341GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n543) );
  NAND2_X1 U608 ( .A1(n545), .A2(n578), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U610 ( .A(G127GAT), .B(n544), .ZN(G1342GAT) );
  XOR2_X1 U611 ( .A(G134GAT), .B(KEYINPUT51), .Z(n547) );
  NAND2_X1 U612 ( .A1(n545), .A2(n558), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(G1343GAT) );
  NAND2_X1 U614 ( .A1(n548), .A2(n570), .ZN(n559) );
  NOR2_X1 U615 ( .A1(n395), .A2(n559), .ZN(n549) );
  XOR2_X1 U616 ( .A(G141GAT), .B(n549), .Z(G1344GAT) );
  NOR2_X1 U617 ( .A1(n550), .A2(n559), .ZN(n555) );
  XOR2_X1 U618 ( .A(KEYINPUT119), .B(KEYINPUT53), .Z(n552) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(KEYINPUT118), .ZN(n551) );
  XNOR2_X1 U620 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U621 ( .A(KEYINPUT52), .B(n553), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(G1345GAT) );
  NOR2_X1 U623 ( .A1(n556), .A2(n559), .ZN(n557) );
  XOR2_X1 U624 ( .A(G155GAT), .B(n557), .Z(G1346GAT) );
  INV_X1 U625 ( .A(n558), .ZN(n560) );
  NOR2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U627 ( .A(G162GAT), .B(n561), .Z(n562) );
  XNOR2_X1 U628 ( .A(KEYINPUT120), .B(n562), .ZN(G1347GAT) );
  NAND2_X1 U629 ( .A1(n565), .A2(n563), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U631 ( .A(G183GAT), .B(KEYINPUT125), .Z(n567) );
  NAND2_X1 U632 ( .A1(n578), .A2(n565), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(G1350GAT) );
  INV_X1 U634 ( .A(n568), .ZN(n569) );
  NAND2_X1 U635 ( .A1(n570), .A2(n569), .ZN(n581) );
  INV_X1 U636 ( .A(n581), .ZN(n579) );
  NAND2_X1 U637 ( .A1(n571), .A2(n579), .ZN(n574) );
  XOR2_X1 U638 ( .A(G197GAT), .B(KEYINPUT60), .Z(n572) );
  XNOR2_X1 U639 ( .A(KEYINPUT59), .B(n572), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  XOR2_X1 U641 ( .A(G204GAT), .B(KEYINPUT61), .Z(n577) );
  NAND2_X1 U642 ( .A1(n579), .A2(n575), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  NAND2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n580), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U647 ( .A(KEYINPUT62), .B(n583), .Z(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

