//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 0 0 0 1 0 1 1 0 1 0 0 0 1 1 0 1 0 1 1 0 0 0 0 0 1 0 1 1 1 0 0 0 0 0 0 0 1 1 1 0 0 0 0 1 1 0 0 0 0 0 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:53 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1287, new_n1288, new_n1289, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1358, new_n1359,
    new_n1360;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(new_n204));
  XOR2_X1   g0004(.A(new_n204), .B(KEYINPUT64), .Z(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  INV_X1    g0013(.A(new_n201), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G50), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n208), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G68), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  INV_X1    g0022(.A(G87), .ZN(new_n223));
  INV_X1    g0023(.A(G250), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n210), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n213), .B(new_n219), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT65), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n235), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  OR2_X1    g0047(.A1(KEYINPUT3), .A2(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G1698), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n250), .A2(G222), .A3(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G77), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n250), .A2(G1698), .ZN(new_n254));
  INV_X1    g0054(.A(G223), .ZN(new_n255));
  OAI221_X1 g0055(.A(new_n252), .B1(new_n253), .B2(new_n250), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G274), .ZN(new_n259));
  AND2_X1   g0059(.A1(G1), .A2(G13), .ZN(new_n260));
  NAND2_X1  g0060(.A1(G33), .A2(G41), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n259), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G41), .ZN(new_n263));
  INV_X1    g0063(.A(G45), .ZN(new_n264));
  AOI21_X1  g0064(.A(G1), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n257), .A2(new_n265), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n267), .B1(G226), .B2(new_n268), .ZN(new_n269));
  AND2_X1   g0069(.A1(new_n258), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G179), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(new_n217), .ZN(new_n276));
  NOR3_X1   g0076(.A1(new_n274), .A2(new_n276), .A3(KEYINPUT68), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(KEYINPUT68), .B1(new_n274), .B2(new_n276), .ZN(new_n279));
  AOI22_X1  g0079(.A1(new_n278), .A2(new_n279), .B1(new_n207), .B2(G20), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G50), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n274), .A2(new_n202), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT67), .ZN(new_n283));
  INV_X1    g0083(.A(G33), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n283), .A2(new_n208), .A3(new_n284), .ZN(new_n285));
  OAI21_X1  g0085(.A(KEYINPUT67), .B1(G20), .B2(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n287), .A2(G150), .B1(G20), .B2(new_n203), .ZN(new_n288));
  XNOR2_X1  g0088(.A(KEYINPUT8), .B(G58), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n208), .A2(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(KEYINPUT66), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT66), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n293), .A2(new_n208), .A3(G33), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n290), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n288), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n276), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n281), .A2(new_n282), .A3(new_n297), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n272), .B(new_n298), .C1(G169), .C2(new_n270), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n268), .A2(G244), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(new_n266), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n250), .A2(G232), .A3(new_n251), .ZN(new_n302));
  INV_X1    g0102(.A(G107), .ZN(new_n303));
  OAI221_X1 g0103(.A(new_n302), .B1(new_n303), .B2(new_n250), .C1(new_n254), .C2(new_n222), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n301), .B1(new_n304), .B2(new_n257), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G190), .ZN(new_n306));
  INV_X1    g0106(.A(G200), .ZN(new_n307));
  INV_X1    g0107(.A(new_n287), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n308), .A2(new_n289), .ZN(new_n309));
  XNOR2_X1  g0109(.A(KEYINPUT15), .B(G87), .ZN(new_n310));
  OAI22_X1  g0110(.A1(new_n310), .A2(new_n291), .B1(new_n208), .B2(new_n253), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n276), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n274), .A2(new_n276), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n253), .B1(new_n207), .B2(G20), .ZN(new_n314));
  AOI22_X1  g0114(.A1(new_n313), .A2(new_n314), .B1(new_n253), .B2(new_n274), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT69), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(KEYINPUT69), .B1(new_n312), .B2(new_n315), .ZN(new_n319));
  OAI221_X1 g0119(.A(new_n306), .B1(new_n307), .B2(new_n305), .C1(new_n318), .C2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n304), .A2(new_n257), .ZN(new_n321));
  INV_X1    g0121(.A(new_n301), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n321), .A2(new_n271), .A3(new_n322), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n323), .B(new_n316), .C1(G169), .C2(new_n305), .ZN(new_n324));
  AND2_X1   g0124(.A1(new_n320), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n298), .A2(KEYINPUT9), .ZN(new_n326));
  AND2_X1   g0126(.A1(new_n297), .A2(new_n282), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT9), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n327), .A2(new_n328), .A3(new_n281), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT10), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n307), .B1(new_n258), .B2(new_n269), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n332), .B1(G190), .B2(new_n270), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n330), .A2(new_n331), .A3(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n331), .B1(new_n330), .B2(new_n333), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n299), .B(new_n325), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  XNOR2_X1  g0137(.A(new_n337), .B(KEYINPUT70), .ZN(new_n338));
  AND2_X1   g0138(.A1(KEYINPUT3), .A2(G33), .ZN(new_n339));
  NOR2_X1   g0139(.A1(KEYINPUT3), .A2(G33), .ZN(new_n340));
  OAI211_X1 g0140(.A(G232), .B(G1698), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  OAI211_X1 g0141(.A(G226), .B(new_n251), .C1(new_n339), .C2(new_n340), .ZN(new_n342));
  NAND2_X1  g0142(.A1(G33), .A2(G97), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n257), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n268), .A2(G238), .B1(new_n265), .B2(new_n262), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT13), .ZN(new_n347));
  AND3_X1   g0147(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n347), .B1(new_n345), .B2(new_n346), .ZN(new_n349));
  OAI21_X1  g0149(.A(G200), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n345), .A2(new_n346), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(KEYINPUT13), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n352), .A2(G190), .A3(new_n353), .ZN(new_n354));
  AND2_X1   g0154(.A1(new_n350), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n287), .A2(G50), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n292), .A2(G77), .A3(new_n294), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n221), .A2(G20), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n356), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT71), .ZN(new_n360));
  AND3_X1   g0160(.A1(new_n359), .A2(new_n360), .A3(new_n276), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n360), .B1(new_n359), .B2(new_n276), .ZN(new_n362));
  OAI21_X1  g0162(.A(KEYINPUT11), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n359), .A2(new_n276), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(KEYINPUT71), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT11), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n359), .A2(new_n360), .A3(new_n276), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n365), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(KEYINPUT12), .B1(new_n273), .B2(G68), .ZN(new_n369));
  OR3_X1    g0169(.A1(new_n273), .A2(KEYINPUT12), .A3(G68), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n221), .B1(new_n207), .B2(G20), .ZN(new_n371));
  AOI22_X1  g0171(.A1(new_n369), .A2(new_n370), .B1(new_n313), .B2(new_n371), .ZN(new_n372));
  AND3_X1   g0172(.A1(new_n363), .A2(new_n368), .A3(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(KEYINPUT72), .B1(new_n355), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n350), .A2(new_n354), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n363), .A2(new_n368), .A3(new_n372), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT72), .ZN(new_n377));
  NOR3_X1   g0177(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n374), .A2(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n290), .A2(new_n273), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n207), .A2(G20), .ZN(new_n382));
  INV_X1    g0182(.A(new_n279), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n382), .B1(new_n383), .B2(new_n277), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n381), .B1(new_n384), .B2(new_n289), .ZN(new_n385));
  INV_X1    g0185(.A(new_n276), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n339), .A2(new_n340), .ZN(new_n387));
  AOI21_X1  g0187(.A(KEYINPUT7), .B1(new_n387), .B2(new_n208), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT7), .ZN(new_n389));
  NOR4_X1   g0189(.A1(new_n339), .A2(new_n340), .A3(new_n389), .A4(G20), .ZN(new_n390));
  OAI21_X1  g0190(.A(G68), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  XNOR2_X1  g0191(.A(G58), .B(G68), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n287), .A2(G159), .B1(new_n392), .B2(G20), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT16), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n386), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n391), .A2(KEYINPUT16), .A3(new_n393), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n385), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  OAI211_X1 g0198(.A(G223), .B(new_n251), .C1(new_n339), .C2(new_n340), .ZN(new_n399));
  OAI211_X1 g0199(.A(G226), .B(G1698), .C1(new_n339), .C2(new_n340), .ZN(new_n400));
  NAND2_X1  g0200(.A1(G33), .A2(G87), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n257), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n260), .A2(new_n261), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n404), .A2(G232), .A3(new_n405), .ZN(new_n406));
  AND2_X1   g0206(.A1(new_n266), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n403), .A2(new_n407), .A3(new_n271), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n266), .A2(new_n406), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n409), .B1(new_n257), .B2(new_n402), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n408), .B1(new_n410), .B2(G169), .ZN(new_n411));
  OAI21_X1  g0211(.A(KEYINPUT18), .B1(new_n398), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n389), .B1(new_n250), .B2(G20), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n387), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n221), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n393), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n395), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n417), .A2(new_n276), .A3(new_n397), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n380), .B1(new_n280), .B2(new_n290), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n411), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT18), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(G190), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n403), .A2(new_n407), .A3(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n424), .B1(new_n410), .B2(G200), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n398), .A2(KEYINPUT17), .A3(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n418), .A2(new_n425), .A3(new_n419), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT17), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n412), .A2(new_n422), .A3(new_n426), .A4(new_n429), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n379), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT73), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n352), .A2(G179), .A3(new_n353), .ZN(new_n433));
  OAI21_X1  g0233(.A(G169), .B1(new_n348), .B2(new_n349), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n433), .B1(new_n434), .B2(KEYINPUT14), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT14), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n352), .A2(new_n353), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n436), .B1(new_n437), .B2(G169), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n432), .B1(new_n435), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n434), .A2(KEYINPUT14), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n437), .A2(new_n436), .A3(G169), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n440), .A2(new_n441), .A3(KEYINPUT73), .A4(new_n433), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(new_n376), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n431), .A2(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n338), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  OAI211_X1 g0247(.A(G264), .B(G1698), .C1(new_n339), .C2(new_n340), .ZN(new_n448));
  OAI211_X1 g0248(.A(G257), .B(new_n251), .C1(new_n339), .C2(new_n340), .ZN(new_n449));
  INV_X1    g0249(.A(G303), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n448), .B(new_n449), .C1(new_n450), .C2(new_n250), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(new_n257), .ZN(new_n452));
  XNOR2_X1  g0252(.A(KEYINPUT5), .B(G41), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n264), .A2(G1), .ZN(new_n454));
  AOI22_X1  g0254(.A1(new_n453), .A2(new_n454), .B1(new_n260), .B2(new_n261), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n207), .A2(G45), .ZN(new_n456));
  NOR2_X1   g0256(.A1(KEYINPUT5), .A2(G41), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(KEYINPUT5), .A2(G41), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n456), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  AOI22_X1  g0260(.A1(new_n455), .A2(G270), .B1(new_n262), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n452), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(G169), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G33), .A2(G283), .ZN(new_n465));
  INV_X1    g0265(.A(G97), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n465), .B(new_n208), .C1(G33), .C2(new_n466), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n467), .B(new_n276), .C1(new_n208), .C2(G116), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT20), .ZN(new_n469));
  XNOR2_X1  g0269(.A(new_n468), .B(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n273), .A2(G116), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n207), .A2(G33), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n273), .A2(new_n472), .A3(new_n217), .A4(new_n275), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n471), .B1(new_n474), .B2(G116), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(KEYINPUT21), .B1(new_n464), .B2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n476), .ZN(new_n478));
  AND2_X1   g0278(.A1(new_n452), .A2(new_n461), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(G190), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n462), .A2(G200), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n478), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT21), .ZN(new_n484));
  INV_X1    g0284(.A(G169), .ZN(new_n485));
  AOI211_X1 g0285(.A(new_n484), .B(new_n485), .C1(new_n452), .C2(new_n461), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n462), .A2(new_n271), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n476), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT80), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OAI211_X1 g0290(.A(KEYINPUT80), .B(new_n476), .C1(new_n486), .C2(new_n487), .ZN(new_n491));
  AOI211_X1 g0291(.A(new_n477), .B(new_n483), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT6), .ZN(new_n493));
  AND2_X1   g0293(.A1(G97), .A2(G107), .ZN(new_n494));
  NOR2_X1   g0294(.A1(G97), .A2(G107), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT74), .ZN(new_n497));
  NAND2_X1  g0297(.A1(KEYINPUT6), .A2(G97), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n497), .B1(new_n498), .B2(G107), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n303), .A2(KEYINPUT74), .A3(KEYINPUT6), .A4(G97), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n496), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(KEYINPUT75), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT75), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n496), .A2(new_n499), .A3(new_n503), .A4(new_n500), .ZN(new_n504));
  AND3_X1   g0304(.A1(new_n502), .A2(G20), .A3(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(G107), .B1(new_n388), .B2(new_n390), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n287), .A2(G77), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n276), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n473), .A2(G97), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT76), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n273), .A2(new_n466), .ZN(new_n512));
  AND3_X1   g0312(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n511), .B1(new_n510), .B2(new_n512), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  OAI211_X1 g0316(.A(G250), .B(G1698), .C1(new_n339), .C2(new_n340), .ZN(new_n517));
  OAI211_X1 g0317(.A(G244), .B(new_n251), .C1(new_n339), .C2(new_n340), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT4), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n465), .B(new_n517), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(G1698), .B1(new_n248), .B2(new_n249), .ZN(new_n521));
  AOI21_X1  g0321(.A(KEYINPUT4), .B1(new_n521), .B2(G244), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n257), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n460), .A2(new_n262), .ZN(new_n524));
  INV_X1    g0324(.A(new_n459), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n454), .B1(new_n525), .B2(new_n457), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n526), .A2(G257), .A3(new_n404), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  AND3_X1   g0329(.A1(new_n523), .A2(new_n529), .A3(new_n423), .ZN(new_n530));
  AOI21_X1  g0330(.A(G200), .B1(new_n523), .B2(new_n529), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n509), .B(new_n516), .C1(new_n530), .C2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n523), .A2(new_n529), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n485), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n523), .A2(new_n529), .A3(new_n271), .ZN(new_n535));
  INV_X1    g0335(.A(new_n507), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n413), .A2(new_n414), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n536), .B1(new_n537), .B2(G107), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n502), .A2(G20), .A3(new_n504), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n386), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n534), .B(new_n535), .C1(new_n540), .C2(new_n515), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT77), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n532), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n542), .B1(new_n532), .B2(new_n541), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT23), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n546), .B1(new_n208), .B2(G107), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n303), .A2(KEYINPUT23), .A3(G20), .ZN(new_n548));
  INV_X1    g0348(.A(G116), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n284), .A2(new_n549), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n547), .A2(new_n548), .B1(new_n550), .B2(new_n208), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n208), .B(G87), .C1(new_n339), .C2(new_n340), .ZN(new_n552));
  XOR2_X1   g0352(.A(KEYINPUT81), .B(KEYINPUT22), .Z(new_n553));
  AND2_X1   g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n552), .A2(new_n553), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n551), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  XOR2_X1   g0356(.A(KEYINPUT82), .B(KEYINPUT24), .Z(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n557), .B(new_n551), .C1(new_n554), .C2(new_n555), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n559), .A2(new_n276), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n474), .A2(G107), .ZN(new_n562));
  OAI211_X1 g0362(.A(KEYINPUT83), .B(KEYINPUT25), .C1(new_n273), .C2(G107), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT83), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT25), .ZN(new_n565));
  AOI21_X1  g0365(.A(G107), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n274), .B(new_n566), .C1(new_n564), .C2(new_n565), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n562), .A2(new_n563), .A3(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT84), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n562), .A2(KEYINPUT84), .A3(new_n563), .A4(new_n567), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n561), .A2(new_n572), .ZN(new_n573));
  OAI211_X1 g0373(.A(G257), .B(G1698), .C1(new_n339), .C2(new_n340), .ZN(new_n574));
  OAI211_X1 g0374(.A(G250), .B(new_n251), .C1(new_n339), .C2(new_n340), .ZN(new_n575));
  NAND2_X1  g0375(.A1(G33), .A2(G294), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT85), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n577), .A2(new_n578), .A3(new_n257), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n455), .A2(G264), .B1(new_n262), .B2(new_n460), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n578), .B1(new_n577), .B2(new_n257), .ZN(new_n582));
  NOR3_X1   g0382(.A1(new_n581), .A2(G190), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n577), .A2(new_n257), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n455), .A2(G264), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n584), .A2(new_n524), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(KEYINPUT86), .B1(new_n586), .B2(new_n307), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n586), .A2(KEYINPUT86), .A3(new_n307), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n573), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n586), .A2(new_n271), .ZN(new_n591));
  INV_X1    g0391(.A(new_n582), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n592), .A2(new_n579), .A3(new_n580), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n591), .B1(G169), .B2(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n386), .B1(new_n556), .B2(new_n558), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n595), .A2(new_n560), .B1(new_n570), .B2(new_n571), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n590), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n222), .A2(new_n251), .ZN(new_n599));
  INV_X1    g0399(.A(G244), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(G1698), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n599), .B(new_n601), .C1(new_n339), .C2(new_n340), .ZN(new_n602));
  INV_X1    g0402(.A(new_n550), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n404), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n404), .A2(G274), .A3(new_n454), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n224), .B1(new_n207), .B2(G45), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n404), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n485), .B1(new_n604), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n262), .A2(new_n454), .B1(new_n404), .B2(new_n606), .ZN(new_n610));
  NOR2_X1   g0410(.A1(G238), .A2(G1698), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n611), .B1(new_n600), .B2(G1698), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n550), .B1(new_n612), .B2(new_n250), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n610), .B(new_n271), .C1(new_n613), .C2(new_n404), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n609), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n208), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n495), .A2(new_n223), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n208), .B(G68), .C1(new_n339), .C2(new_n340), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT19), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n621), .B1(new_n291), .B2(new_n466), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n619), .A2(new_n620), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n276), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n310), .A2(new_n274), .ZN(new_n625));
  INV_X1    g0425(.A(new_n310), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n474), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n624), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT78), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AOI22_X1  g0430(.A1(new_n623), .A2(new_n276), .B1(new_n274), .B2(new_n310), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n631), .A2(KEYINPUT78), .A3(new_n627), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n615), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(G200), .B1(new_n604), .B2(new_n608), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n610), .B(G190), .C1(new_n613), .C2(new_n404), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n474), .A2(G87), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n634), .A2(new_n631), .A3(new_n635), .A4(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(KEYINPUT79), .B1(new_n633), .B2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n615), .ZN(new_n640));
  AND4_X1   g0440(.A1(KEYINPUT78), .A2(new_n624), .A3(new_n625), .A4(new_n627), .ZN(new_n641));
  AOI21_X1  g0441(.A(KEYINPUT78), .B1(new_n631), .B2(new_n627), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT79), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(new_n644), .A3(new_n637), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n639), .A2(new_n645), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n492), .A2(new_n545), .A3(new_n598), .A4(new_n646), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n447), .A2(new_n647), .ZN(G372));
  NOR2_X1   g0448(.A1(new_n298), .A2(KEYINPUT9), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n328), .B1(new_n327), .B2(new_n281), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n333), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(KEYINPUT10), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n334), .ZN(new_n653));
  AND2_X1   g0453(.A1(new_n426), .A2(new_n429), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n316), .B1(new_n305), .B2(G169), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  OAI211_X1 g0457(.A(new_n323), .B(new_n657), .C1(new_n375), .C2(new_n376), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n655), .B1(new_n444), .B2(new_n658), .ZN(new_n659));
  XNOR2_X1  g0459(.A(new_n420), .B(KEYINPUT18), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n653), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n662), .A2(new_n299), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT88), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT87), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n665), .B1(new_n613), .B2(new_n404), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n604), .A2(KEYINPUT87), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n608), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n664), .B1(new_n668), .B2(G169), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n630), .A2(new_n632), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n602), .A2(new_n603), .ZN(new_n671));
  AOI21_X1  g0471(.A(KEYINPUT87), .B1(new_n671), .B2(new_n257), .ZN(new_n672));
  AOI211_X1 g0472(.A(new_n665), .B(new_n404), .C1(new_n602), .C2(new_n603), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n610), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n674), .A2(KEYINPUT88), .A3(new_n485), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n669), .A2(new_n670), .A3(new_n614), .A4(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n631), .A2(new_n636), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n604), .A2(new_n608), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n678), .B1(G190), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n680), .B1(new_n307), .B2(new_n668), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n676), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n532), .A2(new_n541), .ZN(new_n683));
  NOR3_X1   g0483(.A1(new_n682), .A2(new_n590), .A3(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n484), .B1(new_n478), .B2(new_n463), .ZN(new_n685));
  OAI211_X1 g0485(.A(new_n685), .B(new_n488), .C1(new_n594), .C2(new_n596), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n677), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n541), .A2(KEYINPUT89), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n509), .A2(new_n516), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT89), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n689), .A2(new_n690), .A3(new_n535), .A4(new_n534), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n688), .A2(new_n691), .A3(new_n676), .A4(new_n681), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT26), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n540), .A2(new_n515), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n518), .A2(new_n519), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n250), .A2(KEYINPUT4), .A3(G244), .A4(new_n251), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n696), .A2(new_n697), .A3(new_n465), .A4(new_n517), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n528), .B1(new_n698), .B2(new_n257), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n535), .B1(new_n699), .B2(G169), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n695), .A2(new_n700), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n639), .A2(new_n645), .A3(new_n701), .A4(KEYINPUT26), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n694), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n687), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n663), .B1(new_n447), .B2(new_n705), .ZN(G369));
  NAND3_X1  g0506(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n707));
  AND3_X1   g0507(.A1(new_n707), .A2(KEYINPUT90), .A3(KEYINPUT27), .ZN(new_n708));
  AOI21_X1  g0508(.A(KEYINPUT90), .B1(new_n707), .B2(KEYINPUT27), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(G213), .B1(new_n707), .B2(KEYINPUT27), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(G343), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n598), .B1(new_n596), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n597), .A2(new_n715), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n685), .A2(new_n488), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n716), .A2(new_n478), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n490), .A2(new_n491), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n723), .A2(new_n685), .A3(new_n482), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n722), .B1(new_n724), .B2(new_n721), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n719), .A2(G330), .A3(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT91), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n597), .A2(new_n716), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n715), .B1(new_n723), .B2(new_n685), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(new_n598), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n728), .A2(new_n729), .A3(new_n731), .ZN(G399));
  INV_X1    g0532(.A(KEYINPUT92), .ZN(new_n733));
  INV_X1    g0533(.A(new_n211), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n733), .B1(new_n734), .B2(G41), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n211), .A2(KEYINPUT92), .A3(new_n263), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n618), .A2(G116), .ZN(new_n738));
  AND3_X1   g0538(.A1(new_n737), .A2(G1), .A3(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n737), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n739), .B1(new_n216), .B2(new_n740), .ZN(new_n741));
  XOR2_X1   g0541(.A(new_n741), .B(KEYINPUT28), .Z(new_n742));
  AND2_X1   g0542(.A1(new_n584), .A2(new_n585), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n743), .A2(new_n679), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n744), .A2(KEYINPUT30), .A3(new_n487), .A4(new_n699), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT30), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n699), .A2(new_n743), .A3(new_n679), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n479), .A2(G179), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n479), .A2(G179), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n750), .A2(new_n586), .A3(new_n533), .A4(new_n674), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n745), .A2(new_n749), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(new_n715), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT31), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n754), .B1(new_n647), .B2(new_n715), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G330), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n715), .B1(new_n687), .B2(new_n703), .ZN(new_n758));
  OR2_X1    g0558(.A1(new_n758), .A2(KEYINPUT29), .ZN(new_n759));
  INV_X1    g0559(.A(new_n597), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n723), .A2(new_n760), .A3(new_n685), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n684), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n646), .A2(new_n693), .A3(new_n701), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n677), .B1(new_n692), .B2(KEYINPUT26), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n762), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n765), .A2(KEYINPUT29), .A3(new_n716), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n757), .B1(new_n759), .B2(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n742), .B1(new_n767), .B2(G1), .ZN(G364));
  AND2_X1   g0568(.A1(new_n208), .A2(G13), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n207), .B1(new_n769), .B2(G45), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n740), .A2(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n772), .B1(new_n725), .B2(G330), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n773), .B1(G330), .B2(new_n725), .ZN(new_n774));
  INV_X1    g0574(.A(new_n772), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n217), .B1(G20), .B2(new_n485), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n208), .A2(G179), .ZN(new_n778));
  NOR2_X1   g0578(.A1(G190), .A2(G200), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G159), .ZN(new_n782));
  XOR2_X1   g0582(.A(KEYINPUT94), .B(KEYINPUT32), .Z(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n208), .A2(new_n271), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n785), .A2(G190), .A3(G200), .ZN(new_n786));
  NOR3_X1   g0586(.A1(new_n423), .A2(G179), .A3(G200), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n787), .A2(new_n208), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n784), .B1(new_n202), .B2(new_n786), .C1(new_n466), .C2(new_n789), .ZN(new_n790));
  NOR4_X1   g0590(.A1(new_n208), .A2(new_n271), .A3(new_n423), .A4(G200), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(G58), .ZN(new_n793));
  AND2_X1   g0593(.A1(new_n785), .A2(new_n779), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  OAI221_X1 g0595(.A(new_n250), .B1(new_n792), .B2(new_n793), .C1(new_n253), .C2(new_n795), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n785), .A2(new_n423), .A3(G200), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n778), .A2(G190), .A3(G200), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n797), .A2(new_n221), .B1(new_n798), .B2(new_n223), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n778), .A2(new_n423), .A3(G200), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n782), .A2(new_n783), .B1(new_n303), .B2(new_n800), .ZN(new_n801));
  OR4_X1    g0601(.A1(new_n790), .A2(new_n796), .A3(new_n799), .A4(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(G311), .ZN(new_n803));
  INV_X1    g0603(.A(G322), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n803), .A2(new_n795), .B1(new_n792), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n805), .B1(G329), .B2(new_n781), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n387), .B1(new_n798), .B2(new_n450), .ZN(new_n807));
  XOR2_X1   g0607(.A(new_n807), .B(KEYINPUT95), .Z(new_n808));
  INV_X1    g0608(.A(new_n797), .ZN(new_n809));
  XNOR2_X1  g0609(.A(KEYINPUT33), .B(G317), .ZN(new_n810));
  INV_X1    g0610(.A(new_n800), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n809), .A2(new_n810), .B1(new_n811), .B2(G283), .ZN(new_n812));
  INV_X1    g0612(.A(new_n786), .ZN(new_n813));
  AOI22_X1  g0613(.A1(G326), .A2(new_n813), .B1(new_n788), .B2(G294), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n806), .A2(new_n808), .A3(new_n812), .A4(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n777), .B1(new_n802), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(G13), .A2(G33), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n818), .A2(G20), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n819), .A2(new_n776), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n211), .A2(new_n250), .ZN(new_n821));
  XOR2_X1   g0621(.A(new_n821), .B(KEYINPUT93), .Z(new_n822));
  INV_X1    g0622(.A(G355), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n822), .A2(new_n823), .B1(G116), .B2(new_n211), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n734), .A2(new_n250), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(G45), .B2(new_n215), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(G45), .B2(new_n246), .ZN(new_n827));
  OR2_X1    g0627(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n775), .B(new_n816), .C1(new_n820), .C2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n819), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n829), .B1(new_n725), .B2(new_n830), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n774), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(G396));
  OAI22_X1  g0633(.A1(new_n223), .A2(new_n800), .B1(new_n798), .B2(new_n303), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n834), .B1(G283), .B2(new_n809), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n250), .B1(new_n794), .B2(G116), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n781), .A2(G311), .B1(new_n791), .B2(G294), .ZN(new_n837));
  AOI22_X1  g0637(.A1(G303), .A2(new_n813), .B1(new_n788), .B2(G97), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n835), .A2(new_n836), .A3(new_n837), .A4(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(G132), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n250), .B1(new_n780), .B2(new_n840), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n789), .A2(new_n793), .B1(new_n800), .B2(new_n221), .ZN(new_n842));
  INV_X1    g0642(.A(new_n798), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n841), .B(new_n842), .C1(G50), .C2(new_n843), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n844), .B(KEYINPUT97), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT34), .ZN(new_n846));
  INV_X1    g0646(.A(G150), .ZN(new_n847));
  INV_X1    g0647(.A(G137), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n797), .A2(new_n847), .B1(new_n786), .B2(new_n848), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n849), .B(KEYINPUT96), .ZN(new_n850));
  INV_X1    g0650(.A(G143), .ZN(new_n851));
  INV_X1    g0651(.A(G159), .ZN(new_n852));
  OAI221_X1 g0652(.A(new_n850), .B1(new_n851), .B2(new_n792), .C1(new_n852), .C2(new_n795), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n845), .B1(new_n846), .B2(new_n853), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n853), .A2(new_n846), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n839), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT98), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n777), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(new_n857), .B2(new_n856), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n776), .A2(new_n817), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n859), .B(new_n772), .C1(G77), .C2(new_n861), .ZN(new_n862));
  OR2_X1    g0662(.A1(new_n862), .A2(KEYINPUT99), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(KEYINPUT99), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT100), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(new_n324), .B2(new_n716), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n657), .A2(KEYINPUT100), .A3(new_n323), .A4(new_n715), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n715), .A2(new_n316), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n320), .A2(new_n324), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n863), .B(new_n864), .C1(new_n818), .C2(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n758), .A2(new_n871), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n873), .B(KEYINPUT101), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n715), .B1(new_n868), .B2(new_n870), .ZN(new_n875));
  AND4_X1   g0675(.A1(KEYINPUT26), .A2(new_n639), .A3(new_n645), .A4(new_n701), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n876), .B1(new_n693), .B2(new_n692), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n676), .A2(new_n681), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n588), .A2(new_n589), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n596), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n532), .A2(new_n541), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n878), .A2(new_n880), .A3(new_n881), .A4(new_n686), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n676), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n875), .B1(new_n877), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n874), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n775), .B1(new_n886), .B2(new_n757), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n885), .A2(new_n756), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n872), .B1(new_n887), .B2(new_n888), .ZN(G384));
  NAND2_X1  g0689(.A1(new_n502), .A2(new_n504), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT35), .ZN(new_n891));
  OAI211_X1 g0691(.A(G116), .B(new_n218), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n892), .B1(new_n891), .B2(new_n890), .ZN(new_n893));
  XOR2_X1   g0693(.A(KEYINPUT102), .B(KEYINPUT36), .Z(new_n894));
  XNOR2_X1  g0694(.A(new_n893), .B(new_n894), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n216), .B(G77), .C1(new_n793), .C2(new_n221), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n202), .A2(G68), .ZN(new_n897));
  AOI211_X1 g0697(.A(new_n207), .B(G13), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n660), .A2(new_n712), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT37), .ZN(new_n902));
  AND3_X1   g0702(.A1(new_n418), .A2(new_n425), .A3(new_n419), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n903), .A2(new_n420), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n418), .A2(new_n419), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n712), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n902), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n398), .A2(new_n713), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n907), .A2(KEYINPUT104), .B1(new_n430), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n427), .B1(new_n398), .B2(new_n411), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT37), .B1(new_n910), .B2(new_n908), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT104), .ZN(new_n912));
  INV_X1    g0712(.A(new_n420), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n913), .A2(new_n906), .A3(new_n902), .A4(new_n427), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n911), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT38), .B1(new_n909), .B2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n909), .A2(KEYINPUT38), .A3(new_n915), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n373), .A2(new_n716), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n439), .B(new_n442), .C1(new_n374), .C2(new_n378), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n920), .B1(new_n373), .B2(new_n355), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n920), .A2(new_n921), .B1(new_n444), .B2(new_n922), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n324), .A2(new_n715), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n923), .B1(new_n884), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n919), .B1(new_n926), .B2(KEYINPUT103), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT103), .ZN(new_n928));
  AOI211_X1 g0728(.A(new_n928), .B(new_n923), .C1(new_n884), .C2(new_n925), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n901), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT105), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT106), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n911), .A2(new_n933), .A3(new_n914), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n933), .B1(new_n911), .B2(new_n914), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n906), .B1(new_n660), .B2(new_n654), .ZN(new_n937));
  NOR3_X1   g0737(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n918), .B1(new_n938), .B2(KEYINPUT38), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT39), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n444), .A2(new_n715), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n430), .A2(new_n908), .ZN(new_n943));
  OAI211_X1 g0743(.A(KEYINPUT104), .B(KEYINPUT37), .C1(new_n910), .C2(new_n908), .ZN(new_n944));
  AND4_X1   g0744(.A1(KEYINPUT38), .A2(new_n915), .A3(new_n943), .A4(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n916), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(KEYINPUT39), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n941), .A2(new_n942), .A3(new_n947), .ZN(new_n948));
  OAI211_X1 g0748(.A(KEYINPUT105), .B(new_n901), .C1(new_n927), .C2(new_n929), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n932), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n446), .A2(new_n759), .A3(new_n766), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n663), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n950), .B(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n871), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n444), .A2(new_n922), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n920), .B1(new_n379), .B2(new_n443), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n755), .A2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT40), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n911), .A2(new_n914), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(KEYINPUT106), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n961), .A2(new_n943), .A3(new_n934), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT38), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n959), .B1(new_n964), .B2(new_n918), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n755), .B(new_n957), .C1(new_n945), .C2(new_n916), .ZN(new_n966));
  AOI22_X1  g0766(.A1(new_n958), .A2(new_n965), .B1(new_n966), .B2(new_n959), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n446), .A2(new_n755), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n967), .A2(new_n968), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n969), .A2(G330), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n953), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n207), .B2(new_n769), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n953), .A2(new_n971), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n899), .B1(new_n973), .B2(new_n974), .ZN(G367));
  OAI21_X1  g0775(.A(new_n820), .B1(new_n211), .B2(new_n310), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n976), .B1(new_n825), .B2(new_n234), .ZN(new_n977));
  AOI22_X1  g0777(.A1(G294), .A2(new_n809), .B1(new_n811), .B2(G97), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n978), .B1(new_n303), .B2(new_n789), .C1(new_n803), .C2(new_n786), .ZN(new_n979));
  AOI22_X1  g0779(.A1(G283), .A2(new_n794), .B1(new_n781), .B2(G317), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n843), .A2(KEYINPUT46), .A3(G116), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT46), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n798), .B2(new_n549), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n250), .B1(new_n791), .B2(G303), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n980), .A2(new_n981), .A3(new_n983), .A4(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n811), .A2(G77), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n986), .B1(new_n793), .B2(new_n798), .C1(new_n851), .C2(new_n786), .ZN(new_n987));
  AOI22_X1  g0787(.A1(G159), .A2(new_n809), .B1(new_n788), .B2(G68), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n387), .B1(new_n794), .B2(G50), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n781), .A2(G137), .B1(new_n791), .B2(G150), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n988), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n979), .A2(new_n985), .B1(new_n987), .B2(new_n991), .ZN(new_n992));
  XOR2_X1   g0792(.A(KEYINPUT113), .B(KEYINPUT47), .Z(new_n993));
  XNOR2_X1  g0793(.A(new_n992), .B(new_n993), .ZN(new_n994));
  AOI211_X1 g0794(.A(new_n775), .B(new_n977), .C1(new_n994), .C2(new_n776), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n715), .A2(new_n678), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n878), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(new_n676), .B2(new_n996), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n995), .B1(new_n998), .B2(new_n830), .ZN(new_n999));
  NOR3_X1   g0799(.A1(new_n998), .A2(KEYINPUT110), .A3(KEYINPUT43), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n998), .A2(KEYINPUT43), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT109), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n532), .B(new_n541), .C1(new_n695), .C2(new_n716), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n701), .A2(new_n715), .ZN(new_n1006));
  AND2_X1   g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT107), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(KEYINPUT107), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n597), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n715), .B1(new_n1013), .B2(new_n541), .ZN(new_n1014));
  AND2_X1   g0814(.A1(new_n730), .A2(new_n598), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT42), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1015), .A2(new_n1016), .A3(new_n1010), .ZN(new_n1017));
  OAI21_X1  g0817(.A(KEYINPUT42), .B1(new_n731), .B2(new_n1007), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(KEYINPUT108), .B1(new_n1014), .B2(new_n1019), .ZN(new_n1020));
  AND2_X1   g0820(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT108), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n760), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n716), .B1(new_n1023), .B2(new_n701), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1021), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1004), .B1(new_n1020), .B2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n998), .A2(KEYINPUT43), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT110), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1001), .B1(new_n1026), .B2(new_n1029), .ZN(new_n1030));
  NOR3_X1   g0830(.A1(new_n1014), .A2(KEYINPUT108), .A3(new_n1019), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1022), .B1(new_n1021), .B2(new_n1024), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1003), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1033), .A2(new_n1028), .A3(new_n1027), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n728), .B1(new_n1011), .B2(new_n1009), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1030), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n737), .B(KEYINPUT41), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n728), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n731), .A2(new_n729), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT44), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n1040), .A2(KEYINPUT111), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1010), .B1(KEYINPUT111), .B2(new_n1040), .ZN(new_n1043));
  AND3_X1   g0843(.A1(new_n1039), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1042), .B1(new_n1039), .B2(new_n1043), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n731), .A2(new_n729), .A3(new_n1010), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT45), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1047), .B(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1046), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1038), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n730), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1052), .A2(new_n717), .A3(new_n718), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT112), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1015), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  AND2_X1   g0855(.A1(new_n725), .A2(G330), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n731), .A2(KEYINPUT112), .ZN(new_n1057));
  OR3_X1    g0857(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  OAI211_X1 g0858(.A(G330), .B(new_n725), .C1(new_n1055), .C2(new_n1057), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n728), .A2(new_n1046), .A3(new_n1049), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1051), .A2(new_n1060), .A3(new_n767), .A4(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1037), .B1(new_n1062), .B2(new_n767), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1036), .B1(new_n1063), .B2(new_n771), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1035), .B1(new_n1030), .B2(new_n1034), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n999), .B1(new_n1064), .B2(new_n1065), .ZN(G387));
  OAI21_X1  g0866(.A(new_n825), .B1(new_n239), .B2(new_n264), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(new_n738), .B2(new_n822), .ZN(new_n1068));
  OR3_X1    g0868(.A1(new_n289), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1069));
  OAI21_X1  g0869(.A(KEYINPUT50), .B1(new_n289), .B2(G50), .ZN(new_n1070));
  AOI21_X1  g0870(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1069), .A2(new_n738), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n1068), .A2(new_n1072), .B1(new_n303), .B2(new_n734), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n820), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n772), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n221), .A2(new_n795), .B1(new_n792), .B2(new_n202), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n387), .B(new_n1076), .C1(G150), .C2(new_n781), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n809), .A2(new_n290), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n626), .A2(new_n788), .B1(new_n843), .B2(G77), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(G159), .A2(new_n813), .B1(new_n811), .B2(G97), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1077), .A2(new_n1078), .A3(new_n1079), .A4(new_n1080), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(G283), .A2(new_n788), .B1(new_n843), .B2(G294), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(G303), .A2(new_n794), .B1(new_n791), .B2(G317), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n1083), .B1(new_n803), .B2(new_n797), .C1(new_n804), .C2(new_n786), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT48), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1082), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT114), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1086), .B(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1088), .A2(KEYINPUT49), .A3(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n250), .B1(new_n781), .B2(G326), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1090), .B(new_n1091), .C1(new_n549), .C2(new_n800), .ZN(new_n1092));
  AOI21_X1  g0892(.A(KEYINPUT49), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1081), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1075), .B1(new_n1094), .B2(new_n776), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1095), .B1(new_n719), .B2(new_n830), .ZN(new_n1096));
  XOR2_X1   g0896(.A(new_n1096), .B(KEYINPUT115), .Z(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(new_n771), .B2(new_n1060), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1060), .A2(new_n767), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1060), .A2(new_n767), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(new_n740), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1098), .B1(new_n1099), .B2(new_n1101), .ZN(G393));
  NAND2_X1  g0902(.A1(new_n1051), .A2(new_n1061), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n1100), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1104), .A2(new_n740), .A3(new_n1062), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1051), .A2(new_n771), .A3(new_n1061), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n820), .B1(new_n466), .B2(new_n211), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(new_n825), .B2(new_n243), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n813), .A2(G317), .B1(new_n791), .B2(G311), .ZN(new_n1109));
  XOR2_X1   g0909(.A(new_n1109), .B(KEYINPUT52), .Z(new_n1110));
  INV_X1    g0910(.A(G294), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n387), .B1(new_n795), .B2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(G322), .B2(new_n781), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(G116), .A2(new_n788), .B1(new_n811), .B2(G107), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(G303), .A2(new_n809), .B1(new_n843), .B2(G283), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n1110), .A2(new_n1113), .A3(new_n1114), .A4(new_n1115), .ZN(new_n1116));
  OR2_X1    g0916(.A1(new_n1116), .A2(KEYINPUT116), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n792), .A2(new_n852), .B1(new_n786), .B2(new_n847), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(new_n1118), .B(KEYINPUT51), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n250), .B1(new_n851), .B2(new_n780), .C1(new_n795), .C2(new_n289), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n789), .A2(new_n253), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(G87), .B2(new_n811), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(G50), .A2(new_n809), .B1(new_n843), .B2(G68), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1119), .A2(new_n1121), .A3(new_n1123), .A4(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1116), .A2(KEYINPUT116), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1117), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n775), .B(new_n1108), .C1(new_n1127), .C2(new_n776), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(new_n1012), .B2(new_n830), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1105), .A2(new_n1106), .A3(new_n1129), .ZN(G390));
  NAND2_X1  g0930(.A1(new_n955), .A2(new_n956), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n871), .A2(new_n716), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(new_n687), .B2(new_n703), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1131), .B1(new_n1133), .B2(new_n924), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n942), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n941), .A2(new_n947), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n755), .A2(G330), .A3(new_n871), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1138), .A2(new_n923), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n765), .A2(new_n716), .A3(new_n871), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n925), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n1135), .B(new_n939), .C1(new_n1143), .C2(new_n923), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1137), .A2(new_n1140), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n939), .A2(new_n1135), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1146), .B1(new_n1131), .B2(new_n1142), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1139), .B1(new_n1147), .B2(new_n1136), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1145), .A2(new_n1148), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1149), .A2(new_n770), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n941), .A2(new_n947), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n817), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n772), .B1(new_n290), .B2(new_n861), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n813), .A2(G283), .B1(new_n794), .B2(G97), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1154), .B1(new_n303), .B2(new_n797), .ZN(new_n1155));
  XOR2_X1   g0955(.A(new_n1155), .B(KEYINPUT119), .Z(new_n1156));
  OAI221_X1 g0956(.A(new_n387), .B1(new_n780), .B2(new_n1111), .C1(new_n792), .C2(new_n549), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n221), .A2(new_n800), .B1(new_n798), .B2(new_n223), .ZN(new_n1158));
  NOR4_X1   g0958(.A1(new_n1156), .A2(new_n1122), .A3(new_n1157), .A4(new_n1158), .ZN(new_n1159));
  XOR2_X1   g0959(.A(KEYINPUT54), .B(G143), .Z(new_n1160));
  AOI22_X1  g0960(.A1(new_n788), .A2(G159), .B1(new_n794), .B2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n848), .B2(new_n797), .ZN(new_n1162));
  XOR2_X1   g0962(.A(new_n1162), .B(KEYINPUT118), .Z(new_n1163));
  INV_X1    g0963(.A(G125), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n250), .B1(new_n780), .B2(new_n1164), .C1(new_n792), .C2(new_n840), .ZN(new_n1165));
  INV_X1    g0965(.A(G128), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n786), .A2(new_n1166), .B1(new_n800), .B2(new_n202), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n843), .A2(G150), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1168), .B(KEYINPUT53), .ZN(new_n1169));
  NOR4_X1   g0969(.A1(new_n1163), .A2(new_n1165), .A3(new_n1167), .A4(new_n1169), .ZN(new_n1170));
  OR2_X1    g0970(.A1(new_n1159), .A2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1153), .B1(new_n1171), .B2(new_n776), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1150), .B1(new_n1152), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1138), .A2(new_n923), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n1175), .A2(new_n1139), .B1(new_n1133), .B2(new_n924), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1140), .A2(new_n1143), .A3(new_n1174), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n447), .A2(new_n756), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n952), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1178), .A2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n737), .B1(new_n1149), .B2(new_n1181), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1145), .A2(new_n1178), .A3(new_n1148), .A4(new_n1180), .ZN(new_n1183));
  AND3_X1   g0983(.A1(new_n1182), .A2(KEYINPUT117), .A3(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(KEYINPUT117), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1173), .B1(new_n1184), .B2(new_n1185), .ZN(G378));
  AND3_X1   g0986(.A1(new_n941), .A2(new_n947), .A3(new_n942), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n946), .B1(new_n1134), .B2(new_n928), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n926), .A2(KEYINPUT103), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n900), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1187), .B1(new_n1190), .B2(KEYINPUT105), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n298), .A2(new_n712), .ZN(new_n1192));
  AND3_X1   g0992(.A1(new_n653), .A2(new_n299), .A3(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1192), .B1(new_n653), .B2(new_n299), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  OR3_X1    g0996(.A1(new_n1193), .A2(new_n1194), .A3(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1196), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n967), .A2(G330), .A3(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n965), .A2(new_n958), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n966), .A2(new_n959), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1201), .A2(new_n1202), .A3(G330), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1199), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1191), .A2(new_n932), .A3(new_n1200), .A4(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n949), .A2(new_n948), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1208));
  AOI21_X1  g1008(.A(KEYINPUT105), .B1(new_n1208), .B2(new_n901), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1199), .B1(new_n967), .B2(G330), .ZN(new_n1210));
  AND4_X1   g1010(.A1(G330), .A2(new_n1201), .A3(new_n1202), .A4(new_n1199), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n1207), .A2(new_n1209), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n770), .B1(new_n1206), .B2(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n772), .B1(G50), .B2(new_n861), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n800), .A2(new_n793), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n786), .A2(new_n549), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n1215), .B(new_n1216), .C1(G97), .C2(new_n809), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n626), .A2(new_n794), .B1(new_n781), .B2(G283), .ZN(new_n1218));
  AOI211_X1 g1018(.A(G41), .B(new_n250), .C1(new_n791), .C2(G107), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(G68), .A2(new_n788), .B1(new_n843), .B2(G77), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1217), .A2(new_n1218), .A3(new_n1219), .A4(new_n1220), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(new_n1221), .B(KEYINPUT58), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n250), .A2(G41), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n848), .A2(new_n795), .B1(new_n792), .B2(new_n1166), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(G150), .A2(new_n788), .B1(new_n843), .B2(new_n1160), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1226), .B1(new_n1164), .B2(new_n786), .ZN(new_n1227));
  AOI211_X1 g1027(.A(new_n1225), .B(new_n1227), .C1(G132), .C2(new_n809), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n1228), .B(KEYINPUT59), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(KEYINPUT120), .ZN(new_n1230));
  AOI211_X1 g1030(.A(G33), .B(G41), .C1(new_n781), .C2(G124), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1230), .B(new_n1231), .C1(new_n852), .C2(new_n800), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1229), .A2(KEYINPUT120), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n1222), .B1(new_n1223), .B2(new_n1224), .C1(new_n1232), .C2(new_n1233), .ZN(new_n1234));
  OR2_X1    g1034(.A1(new_n1234), .A2(KEYINPUT121), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n777), .B1(new_n1234), .B2(KEYINPUT121), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1214), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1204), .A2(new_n817), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1213), .A2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1205), .A2(new_n1200), .ZN(new_n1242));
  AOI21_X1  g1042(.A(KEYINPUT122), .B1(new_n950), .B2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1206), .A2(new_n1212), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1243), .B1(new_n1244), .B2(KEYINPUT122), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1183), .A2(new_n1180), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(KEYINPUT57), .ZN(new_n1247));
  OAI211_X1 g1047(.A(KEYINPUT123), .B(new_n740), .C1(new_n1245), .C2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1246), .A2(new_n1244), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT57), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1248), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT122), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(new_n1206), .B2(new_n1212), .ZN(new_n1254));
  OAI211_X1 g1054(.A(KEYINPUT57), .B(new_n1246), .C1(new_n1254), .C2(new_n1243), .ZN(new_n1255));
  AOI21_X1  g1055(.A(KEYINPUT123), .B1(new_n1255), .B2(new_n740), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1241), .B1(new_n1252), .B2(new_n1256), .ZN(G375));
  OR2_X1    g1057(.A1(new_n1178), .A2(new_n1180), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1037), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1258), .A2(new_n1259), .A3(new_n1181), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1178), .A2(new_n771), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n781), .A2(G128), .B1(new_n791), .B2(G137), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1262), .B(new_n250), .C1(new_n847), .C2(new_n795), .ZN(new_n1263));
  AOI211_X1 g1063(.A(new_n1215), .B(new_n1263), .C1(G132), .C2(new_n813), .ZN(new_n1264));
  AOI22_X1  g1064(.A1(new_n809), .A2(new_n1160), .B1(new_n788), .B2(G50), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1264), .B(new_n1265), .C1(new_n852), .C2(new_n798), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n780), .A2(new_n450), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n387), .B1(new_n795), .B2(new_n303), .ZN(new_n1268));
  AOI211_X1 g1068(.A(new_n1267), .B(new_n1268), .C1(G283), .C2(new_n791), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n788), .A2(new_n626), .ZN(new_n1270));
  OAI22_X1  g1070(.A1(new_n786), .A2(new_n1111), .B1(new_n798), .B2(new_n466), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1271), .B1(G116), .B2(new_n809), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1269), .A2(new_n986), .A3(new_n1270), .A4(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n777), .B1(new_n1266), .B2(new_n1273), .ZN(new_n1274));
  AOI211_X1 g1074(.A(new_n775), .B(new_n1274), .C1(new_n221), .C2(new_n860), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1275), .B1(new_n1131), .B2(new_n818), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1261), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1260), .A2(new_n1278), .ZN(G381));
  INV_X1    g1079(.A(G375), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1281));
  AND2_X1   g1081(.A1(new_n1173), .A2(new_n1281), .ZN(new_n1282));
  NOR4_X1   g1082(.A1(G393), .A2(G390), .A3(G384), .A4(G396), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1283), .A2(new_n1278), .A3(new_n1260), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1284), .A2(G387), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1280), .A2(new_n1282), .A3(new_n1285), .ZN(G407));
  NAND2_X1  g1086(.A1(new_n714), .A2(G213), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1280), .A2(new_n1282), .A3(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(G407), .A2(new_n1289), .A3(G213), .ZN(G409));
  XNOR2_X1  g1090(.A(G393), .B(G396), .ZN(new_n1291));
  INV_X1    g1091(.A(G390), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(G387), .A2(new_n1292), .ZN(new_n1293));
  OAI211_X1 g1093(.A(G390), .B(new_n999), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1294));
  AND3_X1   g1094(.A1(new_n1291), .A2(new_n1293), .A3(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1293), .A2(KEYINPUT125), .ZN(new_n1296));
  OR2_X1    g1096(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT124), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1297), .A2(new_n1298), .A3(new_n999), .A4(G390), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT125), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(G387), .A2(new_n1300), .A3(new_n1292), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1294), .A2(KEYINPUT124), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1296), .A2(new_n1299), .A3(new_n1301), .A4(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1291), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1295), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT62), .ZN(new_n1307));
  OAI211_X1 g1107(.A(G378), .B(new_n1241), .C1(new_n1252), .C2(new_n1256), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1245), .A2(new_n770), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1239), .B1(new_n1249), .B2(new_n1037), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1282), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1308), .A2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT60), .ZN(new_n1313));
  OR3_X1    g1113(.A1(new_n1178), .A2(new_n1180), .A3(new_n1313), .ZN(new_n1314));
  AND2_X1   g1114(.A1(new_n1314), .A2(new_n740), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1181), .A2(KEYINPUT60), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(new_n1258), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1277), .B1(new_n1315), .B2(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(G384), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1319), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1318), .A2(G384), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  AND4_X1   g1122(.A1(new_n1307), .A2(new_n1312), .A3(new_n1287), .A4(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT61), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1288), .B1(new_n1308), .B2(new_n1311), .ZN(new_n1325));
  OAI211_X1 g1125(.A(G2897), .B(new_n1288), .C1(new_n1320), .C2(new_n1321), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1321), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1288), .A2(G2897), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1327), .A2(new_n1319), .A3(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1326), .A2(new_n1329), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1324), .B1(new_n1325), .B2(new_n1330), .ZN(new_n1331));
  NOR2_X1   g1131(.A1(new_n1323), .A2(new_n1331), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1307), .B1(new_n1325), .B2(new_n1322), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1333), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1306), .B1(new_n1332), .B2(new_n1334), .ZN(new_n1335));
  AND2_X1   g1135(.A1(new_n1299), .A2(new_n1302), .ZN(new_n1336));
  AND3_X1   g1136(.A1(G387), .A2(new_n1300), .A3(new_n1292), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1300), .B1(G387), .B2(new_n1292), .ZN(new_n1338));
  NOR2_X1   g1138(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1291), .B1(new_n1336), .B2(new_n1339), .ZN(new_n1340));
  OAI211_X1 g1140(.A(KEYINPUT126), .B(new_n1324), .C1(new_n1340), .C2(new_n1295), .ZN(new_n1341));
  INV_X1    g1141(.A(KEYINPUT126), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1342), .B1(new_n1305), .B2(KEYINPUT61), .ZN(new_n1343));
  OAI211_X1 g1143(.A(new_n1341), .B(new_n1343), .C1(new_n1325), .C2(new_n1330), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1325), .A2(KEYINPUT63), .A3(new_n1322), .ZN(new_n1345));
  INV_X1    g1145(.A(new_n1345), .ZN(new_n1346));
  AOI21_X1  g1146(.A(KEYINPUT63), .B1(new_n1325), .B2(new_n1322), .ZN(new_n1347));
  NOR3_X1   g1147(.A1(new_n1344), .A2(new_n1346), .A3(new_n1347), .ZN(new_n1348));
  OAI21_X1  g1148(.A(KEYINPUT127), .B1(new_n1335), .B2(new_n1348), .ZN(new_n1349));
  AND2_X1   g1149(.A1(new_n1341), .A2(new_n1343), .ZN(new_n1350));
  INV_X1    g1150(.A(new_n1347), .ZN(new_n1351));
  OR2_X1    g1151(.A1(new_n1325), .A2(new_n1330), .ZN(new_n1352));
  NAND4_X1  g1152(.A1(new_n1350), .A2(new_n1351), .A3(new_n1352), .A4(new_n1345), .ZN(new_n1353));
  INV_X1    g1153(.A(KEYINPUT127), .ZN(new_n1354));
  NOR3_X1   g1154(.A1(new_n1323), .A2(new_n1331), .A3(new_n1333), .ZN(new_n1355));
  OAI211_X1 g1155(.A(new_n1353), .B(new_n1354), .C1(new_n1355), .C2(new_n1306), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1349), .A2(new_n1356), .ZN(G405));
  INV_X1    g1157(.A(new_n1282), .ZN(new_n1358));
  OAI21_X1  g1158(.A(new_n1308), .B1(new_n1280), .B2(new_n1358), .ZN(new_n1359));
  XNOR2_X1  g1159(.A(new_n1359), .B(new_n1322), .ZN(new_n1360));
  XNOR2_X1  g1160(.A(new_n1360), .B(new_n1305), .ZN(G402));
endmodule


