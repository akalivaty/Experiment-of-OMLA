

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592;

  XNOR2_X1 U323 ( .A(n396), .B(n395), .ZN(n402) );
  XNOR2_X1 U324 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U325 ( .A(G15GAT), .B(G22GAT), .ZN(n353) );
  XNOR2_X1 U326 ( .A(n354), .B(G36GAT), .ZN(n355) );
  XNOR2_X1 U327 ( .A(KEYINPUT47), .B(KEYINPUT119), .ZN(n395) );
  XNOR2_X1 U328 ( .A(n356), .B(n355), .ZN(n364) );
  XNOR2_X1 U329 ( .A(n348), .B(n451), .ZN(n349) );
  XNOR2_X1 U330 ( .A(n327), .B(n326), .ZN(n408) );
  XNOR2_X1 U331 ( .A(n350), .B(n349), .ZN(n352) );
  INV_X1 U332 ( .A(n408), .ZN(n328) );
  NOR2_X1 U333 ( .A1(n441), .A2(n527), .ZN(n577) );
  XNOR2_X1 U334 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U335 ( .A(n372), .B(n371), .ZN(n578) );
  NOR2_X1 U336 ( .A1(n543), .A2(n462), .ZN(n572) );
  XOR2_X1 U337 ( .A(KEYINPUT41), .B(n485), .Z(n561) );
  NOR2_X1 U338 ( .A1(n516), .A2(n525), .ZN(n522) );
  XNOR2_X1 U339 ( .A(n416), .B(n415), .ZN(n531) );
  XNOR2_X1 U340 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n463) );
  XNOR2_X1 U341 ( .A(n491), .B(G43GAT), .ZN(n492) );
  XNOR2_X1 U342 ( .A(n464), .B(n463), .ZN(G1351GAT) );
  XNOR2_X1 U343 ( .A(n493), .B(n492), .ZN(G1330GAT) );
  XOR2_X1 U344 ( .A(KEYINPUT75), .B(KEYINPUT11), .Z(n292) );
  XOR2_X1 U345 ( .A(G29GAT), .B(G134GAT), .Z(n427) );
  XNOR2_X1 U346 ( .A(G99GAT), .B(G85GAT), .ZN(n351) );
  XOR2_X1 U347 ( .A(n427), .B(n351), .Z(n291) );
  XNOR2_X1 U348 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U349 ( .A(n293), .B(KEYINPUT76), .Z(n300) );
  XOR2_X1 U350 ( .A(G36GAT), .B(G190GAT), .Z(n412) );
  XOR2_X1 U351 ( .A(G43GAT), .B(G50GAT), .Z(n295) );
  XNOR2_X1 U352 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n294) );
  XNOR2_X1 U353 ( .A(n295), .B(n294), .ZN(n366) );
  XOR2_X1 U354 ( .A(n412), .B(n366), .Z(n297) );
  NAND2_X1 U355 ( .A1(G232GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U356 ( .A(n297), .B(n296), .ZN(n298) );
  XNOR2_X1 U357 ( .A(G218GAT), .B(n298), .ZN(n299) );
  XNOR2_X1 U358 ( .A(n300), .B(n299), .ZN(n308) );
  XOR2_X1 U359 ( .A(KEYINPUT64), .B(KEYINPUT78), .Z(n302) );
  XNOR2_X1 U360 ( .A(KEYINPUT77), .B(KEYINPUT9), .ZN(n301) );
  XNOR2_X1 U361 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U362 ( .A(KEYINPUT10), .B(G92GAT), .Z(n304) );
  XNOR2_X1 U363 ( .A(G162GAT), .B(G106GAT), .ZN(n303) );
  XNOR2_X1 U364 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U365 ( .A(n306), .B(n305), .Z(n307) );
  XNOR2_X1 U366 ( .A(n308), .B(n307), .ZN(n567) );
  XOR2_X1 U367 ( .A(KEYINPUT86), .B(KEYINPUT82), .Z(n310) );
  XNOR2_X1 U368 ( .A(G15GAT), .B(KEYINPUT83), .ZN(n309) );
  XNOR2_X1 U369 ( .A(n310), .B(n309), .ZN(n323) );
  XOR2_X1 U370 ( .A(G99GAT), .B(G134GAT), .Z(n312) );
  XNOR2_X1 U371 ( .A(G43GAT), .B(G190GAT), .ZN(n311) );
  XNOR2_X1 U372 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U373 ( .A(G71GAT), .B(G176GAT), .Z(n314) );
  XNOR2_X1 U374 ( .A(KEYINPUT20), .B(KEYINPUT84), .ZN(n313) );
  XNOR2_X1 U375 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U376 ( .A(n316), .B(n315), .Z(n321) );
  XOR2_X1 U377 ( .A(G113GAT), .B(KEYINPUT0), .Z(n428) );
  XOR2_X1 U378 ( .A(G127GAT), .B(G120GAT), .Z(n318) );
  NAND2_X1 U379 ( .A1(G227GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U380 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U381 ( .A(n428), .B(n319), .ZN(n320) );
  XNOR2_X1 U382 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U383 ( .A(n323), .B(n322), .ZN(n329) );
  XOR2_X1 U384 ( .A(KEYINPUT85), .B(G183GAT), .Z(n325) );
  XNOR2_X1 U385 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n324) );
  XNOR2_X1 U386 ( .A(n325), .B(n324), .ZN(n327) );
  XOR2_X1 U387 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n326) );
  XOR2_X1 U388 ( .A(n329), .B(n328), .Z(n543) );
  INV_X1 U389 ( .A(G92GAT), .ZN(n330) );
  NAND2_X1 U390 ( .A1(G64GAT), .A2(n330), .ZN(n333) );
  INV_X1 U391 ( .A(G64GAT), .ZN(n331) );
  NAND2_X1 U392 ( .A1(n331), .A2(G92GAT), .ZN(n332) );
  NAND2_X1 U393 ( .A1(n333), .A2(n332), .ZN(n335) );
  XNOR2_X1 U394 ( .A(G176GAT), .B(G204GAT), .ZN(n334) );
  XNOR2_X1 U395 ( .A(n335), .B(n334), .ZN(n406) );
  XNOR2_X1 U396 ( .A(G120GAT), .B(G148GAT), .ZN(n336) );
  XNOR2_X1 U397 ( .A(n336), .B(G57GAT), .ZN(n425) );
  XNOR2_X1 U398 ( .A(n406), .B(n425), .ZN(n344) );
  INV_X1 U399 ( .A(n344), .ZN(n342) );
  XOR2_X1 U400 ( .A(KEYINPUT31), .B(KEYINPUT74), .Z(n338) );
  NAND2_X1 U401 ( .A1(G230GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U402 ( .A(n338), .B(n337), .ZN(n340) );
  INV_X1 U403 ( .A(KEYINPUT73), .ZN(n339) );
  XNOR2_X1 U404 ( .A(n340), .B(n339), .ZN(n343) );
  INV_X1 U405 ( .A(n343), .ZN(n341) );
  NAND2_X1 U406 ( .A1(n342), .A2(n341), .ZN(n346) );
  NAND2_X1 U407 ( .A1(n344), .A2(n343), .ZN(n345) );
  NAND2_X1 U408 ( .A1(n346), .A2(n345), .ZN(n347) );
  XNOR2_X1 U409 ( .A(n347), .B(KEYINPUT33), .ZN(n350) );
  XOR2_X1 U410 ( .A(G71GAT), .B(KEYINPUT13), .Z(n387) );
  XOR2_X1 U411 ( .A(n387), .B(KEYINPUT32), .Z(n348) );
  XOR2_X1 U412 ( .A(G106GAT), .B(G78GAT), .Z(n451) );
  XOR2_X1 U413 ( .A(n352), .B(n351), .Z(n485) );
  XNOR2_X1 U414 ( .A(n353), .B(KEYINPUT71), .ZN(n383) );
  XOR2_X1 U415 ( .A(G29GAT), .B(n383), .Z(n356) );
  NAND2_X1 U416 ( .A1(G229GAT), .A2(G233GAT), .ZN(n354) );
  XOR2_X1 U417 ( .A(G197GAT), .B(G141GAT), .Z(n358) );
  XNOR2_X1 U418 ( .A(G169GAT), .B(G113GAT), .ZN(n357) );
  XNOR2_X1 U419 ( .A(n358), .B(n357), .ZN(n362) );
  XOR2_X1 U420 ( .A(KEYINPUT66), .B(KEYINPUT67), .Z(n360) );
  XNOR2_X1 U421 ( .A(G8GAT), .B(KEYINPUT72), .ZN(n359) );
  XNOR2_X1 U422 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U423 ( .A(n362), .B(n361), .Z(n363) );
  XNOR2_X1 U424 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U425 ( .A(n365), .B(KEYINPUT29), .Z(n372) );
  XNOR2_X1 U426 ( .A(n366), .B(KEYINPUT69), .ZN(n370) );
  XOR2_X1 U427 ( .A(KEYINPUT70), .B(G1GAT), .Z(n368) );
  XNOR2_X1 U428 ( .A(KEYINPUT30), .B(KEYINPUT68), .ZN(n367) );
  XNOR2_X1 U429 ( .A(n368), .B(n367), .ZN(n369) );
  INV_X1 U430 ( .A(n578), .ZN(n570) );
  NAND2_X1 U431 ( .A1(n561), .A2(n570), .ZN(n375) );
  XOR2_X1 U432 ( .A(KEYINPUT46), .B(KEYINPUT118), .Z(n373) );
  XOR2_X1 U433 ( .A(KEYINPUT117), .B(n373), .Z(n374) );
  XNOR2_X1 U434 ( .A(n375), .B(n374), .ZN(n376) );
  NOR2_X1 U435 ( .A1(n376), .A2(n567), .ZN(n394) );
  XOR2_X1 U436 ( .A(G57GAT), .B(G64GAT), .Z(n378) );
  XNOR2_X1 U437 ( .A(G211GAT), .B(G78GAT), .ZN(n377) );
  XNOR2_X1 U438 ( .A(n378), .B(n377), .ZN(n382) );
  XOR2_X1 U439 ( .A(KEYINPUT15), .B(KEYINPUT80), .Z(n380) );
  XNOR2_X1 U440 ( .A(KEYINPUT81), .B(KEYINPUT12), .ZN(n379) );
  XNOR2_X1 U441 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U442 ( .A(n382), .B(n381), .ZN(n393) );
  XOR2_X1 U443 ( .A(G8GAT), .B(KEYINPUT79), .Z(n407) );
  XOR2_X1 U444 ( .A(n383), .B(KEYINPUT14), .Z(n385) );
  NAND2_X1 U445 ( .A1(G231GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U446 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U447 ( .A(n407), .B(n386), .ZN(n391) );
  XOR2_X1 U448 ( .A(G1GAT), .B(G127GAT), .Z(n422) );
  XOR2_X1 U449 ( .A(n422), .B(n387), .Z(n389) );
  XNOR2_X1 U450 ( .A(G183GAT), .B(G155GAT), .ZN(n388) );
  XNOR2_X1 U451 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U452 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U453 ( .A(n393), .B(n392), .Z(n573) );
  INV_X1 U454 ( .A(n573), .ZN(n585) );
  NAND2_X1 U455 ( .A1(n394), .A2(n585), .ZN(n396) );
  XNOR2_X1 U456 ( .A(KEYINPUT36), .B(KEYINPUT107), .ZN(n397) );
  XNOR2_X1 U457 ( .A(n397), .B(n567), .ZN(n590) );
  NOR2_X1 U458 ( .A1(n585), .A2(n590), .ZN(n398) );
  XOR2_X1 U459 ( .A(KEYINPUT45), .B(n398), .Z(n399) );
  NOR2_X1 U460 ( .A1(n485), .A2(n399), .ZN(n400) );
  NAND2_X1 U461 ( .A1(n400), .A2(n578), .ZN(n401) );
  NAND2_X1 U462 ( .A1(n402), .A2(n401), .ZN(n403) );
  XNOR2_X1 U463 ( .A(n403), .B(KEYINPUT48), .ZN(n558) );
  XOR2_X1 U464 ( .A(G211GAT), .B(KEYINPUT21), .Z(n405) );
  XNOR2_X1 U465 ( .A(G197GAT), .B(G218GAT), .ZN(n404) );
  XNOR2_X1 U466 ( .A(n405), .B(n404), .ZN(n450) );
  XNOR2_X1 U467 ( .A(n406), .B(n450), .ZN(n416) );
  XOR2_X1 U468 ( .A(n407), .B(KEYINPUT97), .Z(n410) );
  XOR2_X1 U469 ( .A(n408), .B(KEYINPUT98), .Z(n409) );
  XNOR2_X1 U470 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U471 ( .A(n412), .B(n411), .Z(n414) );
  NAND2_X1 U472 ( .A1(G226GAT), .A2(G233GAT), .ZN(n413) );
  XNOR2_X1 U473 ( .A(n414), .B(n413), .ZN(n415) );
  AND2_X1 U474 ( .A1(n558), .A2(n531), .ZN(n418) );
  XNOR2_X1 U475 ( .A(KEYINPUT125), .B(KEYINPUT54), .ZN(n417) );
  XNOR2_X1 U476 ( .A(n418), .B(n417), .ZN(n441) );
  XOR2_X1 U477 ( .A(KEYINPUT92), .B(KEYINPUT5), .Z(n420) );
  XNOR2_X1 U478 ( .A(KEYINPUT94), .B(KEYINPUT4), .ZN(n419) );
  XNOR2_X1 U479 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U480 ( .A(n421), .B(KEYINPUT6), .Z(n424) );
  XNOR2_X1 U481 ( .A(G85GAT), .B(n422), .ZN(n423) );
  XNOR2_X1 U482 ( .A(n424), .B(n423), .ZN(n426) );
  XOR2_X1 U483 ( .A(n426), .B(n425), .Z(n430) );
  XNOR2_X1 U484 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U485 ( .A(n430), .B(n429), .ZN(n434) );
  XOR2_X1 U486 ( .A(KEYINPUT93), .B(KEYINPUT95), .Z(n432) );
  NAND2_X1 U487 ( .A1(G225GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U488 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U489 ( .A(n434), .B(n433), .Z(n440) );
  XOR2_X1 U490 ( .A(KEYINPUT3), .B(G162GAT), .Z(n436) );
  XNOR2_X1 U491 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n435) );
  XNOR2_X1 U492 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U493 ( .A(G141GAT), .B(n437), .Z(n458) );
  INV_X1 U494 ( .A(n458), .ZN(n438) );
  XOR2_X1 U495 ( .A(n438), .B(KEYINPUT1), .Z(n439) );
  XNOR2_X1 U496 ( .A(n440), .B(n439), .ZN(n473) );
  XOR2_X1 U497 ( .A(KEYINPUT96), .B(n473), .Z(n475) );
  INV_X1 U498 ( .A(n475), .ZN(n527) );
  XOR2_X1 U499 ( .A(KEYINPUT91), .B(KEYINPUT24), .Z(n443) );
  XNOR2_X1 U500 ( .A(G50GAT), .B(KEYINPUT23), .ZN(n442) );
  XNOR2_X1 U501 ( .A(n443), .B(n442), .ZN(n447) );
  XOR2_X1 U502 ( .A(G148GAT), .B(G204GAT), .Z(n445) );
  XNOR2_X1 U503 ( .A(G22GAT), .B(KEYINPUT87), .ZN(n444) );
  XNOR2_X1 U504 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U505 ( .A(n447), .B(n446), .Z(n457) );
  XOR2_X1 U506 ( .A(KEYINPUT90), .B(KEYINPUT89), .Z(n449) );
  XNOR2_X1 U507 ( .A(KEYINPUT22), .B(KEYINPUT88), .ZN(n448) );
  XNOR2_X1 U508 ( .A(n449), .B(n448), .ZN(n455) );
  XOR2_X1 U509 ( .A(n451), .B(n450), .Z(n453) );
  NAND2_X1 U510 ( .A1(G228GAT), .A2(G233GAT), .ZN(n452) );
  XNOR2_X1 U511 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U512 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U513 ( .A(n457), .B(n456), .ZN(n459) );
  XOR2_X1 U514 ( .A(n459), .B(n458), .Z(n476) );
  NAND2_X1 U515 ( .A1(n577), .A2(n476), .ZN(n461) );
  INV_X1 U516 ( .A(KEYINPUT55), .ZN(n460) );
  NAND2_X1 U517 ( .A1(n567), .A2(n572), .ZN(n464) );
  INV_X1 U518 ( .A(n543), .ZN(n533) );
  NAND2_X1 U519 ( .A1(n531), .A2(n533), .ZN(n465) );
  NAND2_X1 U520 ( .A1(n465), .A2(n476), .ZN(n466) );
  XNOR2_X1 U521 ( .A(n466), .B(KEYINPUT100), .ZN(n467) );
  XNOR2_X1 U522 ( .A(n467), .B(KEYINPUT25), .ZN(n471) );
  NOR2_X1 U523 ( .A1(n476), .A2(n533), .ZN(n468) );
  XOR2_X1 U524 ( .A(n468), .B(KEYINPUT26), .Z(n575) );
  XNOR2_X1 U525 ( .A(n531), .B(KEYINPUT99), .ZN(n469) );
  XNOR2_X1 U526 ( .A(n469), .B(KEYINPUT27), .ZN(n474) );
  NOR2_X1 U527 ( .A1(n575), .A2(n474), .ZN(n470) );
  NOR2_X1 U528 ( .A1(n471), .A2(n470), .ZN(n472) );
  NOR2_X1 U529 ( .A1(n473), .A2(n472), .ZN(n480) );
  NOR2_X1 U530 ( .A1(n475), .A2(n474), .ZN(n557) );
  XOR2_X1 U531 ( .A(n476), .B(KEYINPUT65), .Z(n477) );
  XOR2_X1 U532 ( .A(KEYINPUT28), .B(n477), .Z(n536) );
  INV_X1 U533 ( .A(n536), .ZN(n478) );
  NAND2_X1 U534 ( .A1(n557), .A2(n478), .ZN(n542) );
  NOR2_X1 U535 ( .A1(n533), .A2(n542), .ZN(n479) );
  NOR2_X1 U536 ( .A1(n480), .A2(n479), .ZN(n481) );
  XNOR2_X1 U537 ( .A(KEYINPUT101), .B(n481), .ZN(n498) );
  INV_X1 U538 ( .A(n590), .ZN(n482) );
  AND2_X1 U539 ( .A1(n498), .A2(n482), .ZN(n483) );
  NAND2_X1 U540 ( .A1(n483), .A2(n585), .ZN(n484) );
  XOR2_X1 U541 ( .A(KEYINPUT37), .B(n484), .Z(n526) );
  INV_X1 U542 ( .A(n485), .ZN(n582) );
  NAND2_X1 U543 ( .A1(n570), .A2(n582), .ZN(n500) );
  NOR2_X1 U544 ( .A1(n526), .A2(n500), .ZN(n487) );
  XNOR2_X1 U545 ( .A(KEYINPUT38), .B(KEYINPUT108), .ZN(n486) );
  XNOR2_X1 U546 ( .A(n487), .B(n486), .ZN(n513) );
  NAND2_X1 U547 ( .A1(n513), .A2(n527), .ZN(n490) );
  XOR2_X1 U548 ( .A(G29GAT), .B(KEYINPUT39), .Z(n488) );
  XNOR2_X1 U549 ( .A(n488), .B(KEYINPUT106), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n490), .B(n489), .ZN(G1328GAT) );
  NAND2_X1 U551 ( .A1(n513), .A2(n533), .ZN(n493) );
  XOR2_X1 U552 ( .A(KEYINPUT40), .B(KEYINPUT109), .Z(n491) );
  NAND2_X1 U553 ( .A1(n572), .A2(n561), .ZN(n496) );
  XOR2_X1 U554 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n494) );
  XNOR2_X1 U555 ( .A(n494), .B(G176GAT), .ZN(n495) );
  XNOR2_X1 U556 ( .A(n496), .B(n495), .ZN(G1349GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT34), .B(KEYINPUT103), .Z(n503) );
  NOR2_X1 U558 ( .A1(n585), .A2(n567), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n497), .B(KEYINPUT16), .ZN(n499) );
  NAND2_X1 U560 ( .A1(n499), .A2(n498), .ZN(n516) );
  NOR2_X1 U561 ( .A1(n500), .A2(n516), .ZN(n501) );
  XNOR2_X1 U562 ( .A(KEYINPUT102), .B(n501), .ZN(n510) );
  NAND2_X1 U563 ( .A1(n510), .A2(n527), .ZN(n502) );
  XNOR2_X1 U564 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U565 ( .A(G1GAT), .B(n504), .ZN(G1324GAT) );
  NAND2_X1 U566 ( .A1(n510), .A2(n531), .ZN(n505) );
  XNOR2_X1 U567 ( .A(n505), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U568 ( .A(KEYINPUT35), .B(KEYINPUT105), .Z(n507) );
  NAND2_X1 U569 ( .A1(n533), .A2(n510), .ZN(n506) );
  XNOR2_X1 U570 ( .A(n507), .B(n506), .ZN(n509) );
  XOR2_X1 U571 ( .A(G15GAT), .B(KEYINPUT104), .Z(n508) );
  XNOR2_X1 U572 ( .A(n509), .B(n508), .ZN(G1326GAT) );
  NAND2_X1 U573 ( .A1(n510), .A2(n536), .ZN(n511) );
  XNOR2_X1 U574 ( .A(n511), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U575 ( .A1(n513), .A2(n531), .ZN(n512) );
  XNOR2_X1 U576 ( .A(n512), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U577 ( .A1(n513), .A2(n536), .ZN(n514) );
  XNOR2_X1 U578 ( .A(n514), .B(KEYINPUT110), .ZN(n515) );
  XNOR2_X1 U579 ( .A(G50GAT), .B(n515), .ZN(G1331GAT) );
  XNOR2_X1 U580 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n518) );
  NAND2_X1 U581 ( .A1(n561), .A2(n578), .ZN(n525) );
  NAND2_X1 U582 ( .A1(n522), .A2(n527), .ZN(n517) );
  XNOR2_X1 U583 ( .A(n518), .B(n517), .ZN(G1332GAT) );
  XOR2_X1 U584 ( .A(G64GAT), .B(KEYINPUT111), .Z(n520) );
  NAND2_X1 U585 ( .A1(n522), .A2(n531), .ZN(n519) );
  XNOR2_X1 U586 ( .A(n520), .B(n519), .ZN(G1333GAT) );
  NAND2_X1 U587 ( .A1(n522), .A2(n533), .ZN(n521) );
  XNOR2_X1 U588 ( .A(n521), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U589 ( .A(G78GAT), .B(KEYINPUT43), .Z(n524) );
  NAND2_X1 U590 ( .A1(n522), .A2(n536), .ZN(n523) );
  XNOR2_X1 U591 ( .A(n524), .B(n523), .ZN(G1335GAT) );
  XOR2_X1 U592 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n529) );
  NOR2_X1 U593 ( .A1(n526), .A2(n525), .ZN(n537) );
  NAND2_X1 U594 ( .A1(n537), .A2(n527), .ZN(n528) );
  XNOR2_X1 U595 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U596 ( .A(G85GAT), .B(n530), .ZN(G1336GAT) );
  NAND2_X1 U597 ( .A1(n537), .A2(n531), .ZN(n532) );
  XNOR2_X1 U598 ( .A(n532), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U599 ( .A1(n537), .A2(n533), .ZN(n534) );
  XNOR2_X1 U600 ( .A(n534), .B(KEYINPUT114), .ZN(n535) );
  XNOR2_X1 U601 ( .A(G99GAT), .B(n535), .ZN(G1338GAT) );
  XNOR2_X1 U602 ( .A(G106GAT), .B(KEYINPUT115), .ZN(n541) );
  XOR2_X1 U603 ( .A(KEYINPUT44), .B(KEYINPUT116), .Z(n539) );
  NAND2_X1 U604 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U605 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n541), .B(n540), .ZN(G1339GAT) );
  NOR2_X1 U607 ( .A1(n543), .A2(n542), .ZN(n544) );
  NAND2_X1 U608 ( .A1(n544), .A2(n558), .ZN(n545) );
  XOR2_X1 U609 ( .A(KEYINPUT120), .B(n545), .Z(n553) );
  NAND2_X1 U610 ( .A1(n553), .A2(n570), .ZN(n546) );
  XNOR2_X1 U611 ( .A(n546), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U612 ( .A(G120GAT), .B(KEYINPUT49), .Z(n548) );
  NAND2_X1 U613 ( .A1(n561), .A2(n553), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(G1341GAT) );
  XNOR2_X1 U615 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n552) );
  XOR2_X1 U616 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n550) );
  NAND2_X1 U617 ( .A1(n553), .A2(n573), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(G1342GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT51), .B(KEYINPUT123), .Z(n555) );
  NAND2_X1 U621 ( .A1(n553), .A2(n567), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U623 ( .A(G134GAT), .B(n556), .Z(G1343GAT) );
  NAND2_X1 U624 ( .A1(n558), .A2(n557), .ZN(n559) );
  NOR2_X1 U625 ( .A1(n575), .A2(n559), .ZN(n566) );
  NAND2_X1 U626 ( .A1(n566), .A2(n570), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n560), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n563) );
  NAND2_X1 U629 ( .A1(n566), .A2(n561), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U631 ( .A(G148GAT), .B(n564), .ZN(G1345GAT) );
  NAND2_X1 U632 ( .A1(n573), .A2(n566), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n565), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U634 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n568), .B(KEYINPUT124), .ZN(n569) );
  XNOR2_X1 U636 ( .A(G162GAT), .B(n569), .ZN(G1347GAT) );
  NAND2_X1 U637 ( .A1(n570), .A2(n572), .ZN(n571) );
  XNOR2_X1 U638 ( .A(G169GAT), .B(n571), .ZN(G1348GAT) );
  NAND2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n574), .B(G183GAT), .ZN(G1350GAT) );
  INV_X1 U641 ( .A(n575), .ZN(n576) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n589) );
  NOR2_X1 U643 ( .A1(n578), .A2(n589), .ZN(n580) );
  XNOR2_X1 U644 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(G197GAT), .B(n581), .ZN(G1352GAT) );
  NOR2_X1 U647 ( .A1(n582), .A2(n589), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1353GAT) );
  NOR2_X1 U650 ( .A1(n585), .A2(n589), .ZN(n586) );
  XOR2_X1 U651 ( .A(G211GAT), .B(n586), .Z(G1354GAT) );
  XOR2_X1 U652 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n588) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n587) );
  XNOR2_X1 U654 ( .A(n588), .B(n587), .ZN(n592) );
  NOR2_X1 U655 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U656 ( .A(n592), .B(n591), .Z(G1355GAT) );
endmodule

