

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591;

  NOR2_X1 U324 ( .A1(n538), .A2(n478), .ZN(n575) );
  NOR2_X1 U325 ( .A1(n467), .A2(n466), .ZN(n469) );
  XNOR2_X1 U326 ( .A(n464), .B(KEYINPUT97), .ZN(n487) );
  NAND2_X1 U327 ( .A1(n411), .A2(n529), .ZN(n412) );
  INV_X1 U328 ( .A(n554), .ZN(n411) );
  XNOR2_X1 U329 ( .A(n448), .B(KEYINPUT125), .ZN(n585) );
  AND2_X1 U330 ( .A1(n475), .A2(n552), .ZN(n448) );
  XNOR2_X1 U331 ( .A(n306), .B(n305), .ZN(n312) );
  XOR2_X1 U332 ( .A(n445), .B(n444), .Z(n531) );
  XOR2_X1 U333 ( .A(n416), .B(G204GAT), .Z(n292) );
  AND2_X1 U334 ( .A1(G230GAT), .A2(G233GAT), .ZN(n293) );
  XOR2_X1 U335 ( .A(G211GAT), .B(KEYINPUT21), .Z(n294) );
  XOR2_X1 U336 ( .A(n355), .B(n414), .Z(n295) );
  XOR2_X1 U337 ( .A(n406), .B(n405), .Z(n296) );
  OR2_X1 U338 ( .A1(n386), .A2(n385), .ZN(n387) );
  XNOR2_X1 U339 ( .A(n438), .B(n293), .ZN(n353) );
  NOR2_X1 U340 ( .A1(n463), .A2(n462), .ZN(n464) );
  XNOR2_X1 U341 ( .A(n353), .B(n424), .ZN(n354) );
  XNOR2_X1 U342 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U343 ( .A(n407), .B(n296), .ZN(n408) );
  XNOR2_X1 U344 ( .A(n361), .B(n360), .ZN(n363) );
  XNOR2_X1 U345 ( .A(n312), .B(n311), .ZN(n561) );
  XNOR2_X1 U346 ( .A(n409), .B(n408), .ZN(n410) );
  INV_X1 U347 ( .A(G218GAT), .ZN(n449) );
  INV_X1 U348 ( .A(G43GAT), .ZN(n471) );
  XNOR2_X1 U349 ( .A(n449), .B(KEYINPUT62), .ZN(n450) );
  XNOR2_X1 U350 ( .A(n479), .B(G183GAT), .ZN(n480) );
  XNOR2_X1 U351 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U352 ( .A(n451), .B(n450), .ZN(G1355GAT) );
  XNOR2_X1 U353 ( .A(n481), .B(n480), .ZN(G1350GAT) );
  XNOR2_X1 U354 ( .A(n474), .B(n473), .ZN(G1330GAT) );
  XOR2_X1 U355 ( .A(G43GAT), .B(G29GAT), .Z(n298) );
  XNOR2_X1 U356 ( .A(KEYINPUT7), .B(G50GAT), .ZN(n297) );
  XNOR2_X1 U357 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U358 ( .A(n299), .B(KEYINPUT68), .Z(n301) );
  XNOR2_X1 U359 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n300) );
  XNOR2_X1 U360 ( .A(n301), .B(n300), .ZN(n337) );
  XOR2_X1 U361 ( .A(KEYINPUT65), .B(KEYINPUT10), .Z(n303) );
  XNOR2_X1 U362 ( .A(KEYINPUT66), .B(KEYINPUT9), .ZN(n302) );
  XNOR2_X1 U363 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U364 ( .A(n337), .B(n304), .ZN(n306) );
  XOR2_X1 U365 ( .A(G190GAT), .B(G134GAT), .Z(n437) );
  XNOR2_X1 U366 ( .A(n437), .B(KEYINPUT77), .ZN(n305) );
  XOR2_X1 U367 ( .A(G92GAT), .B(G85GAT), .Z(n308) );
  XNOR2_X1 U368 ( .A(G99GAT), .B(G106GAT), .ZN(n307) );
  XNOR2_X1 U369 ( .A(n308), .B(n307), .ZN(n355) );
  XOR2_X1 U370 ( .A(G218GAT), .B(G162GAT), .Z(n414) );
  NAND2_X1 U371 ( .A1(G232GAT), .A2(G233GAT), .ZN(n309) );
  XNOR2_X1 U372 ( .A(n295), .B(n309), .ZN(n310) );
  XOR2_X1 U373 ( .A(n310), .B(KEYINPUT11), .Z(n311) );
  XOR2_X1 U374 ( .A(KEYINPUT78), .B(n561), .Z(n483) );
  INV_X1 U375 ( .A(n483), .ZN(n576) );
  XOR2_X1 U376 ( .A(KEYINPUT36), .B(n576), .Z(n467) );
  XOR2_X1 U377 ( .A(G148GAT), .B(G120GAT), .Z(n314) );
  XNOR2_X1 U378 ( .A(G141GAT), .B(G1GAT), .ZN(n313) );
  XNOR2_X1 U379 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U380 ( .A(KEYINPUT4), .B(KEYINPUT90), .Z(n316) );
  XNOR2_X1 U381 ( .A(KEYINPUT1), .B(KEYINPUT6), .ZN(n315) );
  XNOR2_X1 U382 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U383 ( .A(n318), .B(n317), .Z(n323) );
  XOR2_X1 U384 ( .A(KEYINPUT5), .B(KEYINPUT91), .Z(n320) );
  NAND2_X1 U385 ( .A1(G225GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U386 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U387 ( .A(G57GAT), .B(n321), .ZN(n322) );
  XNOR2_X1 U388 ( .A(n323), .B(n322), .ZN(n328) );
  XNOR2_X1 U389 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n324) );
  XNOR2_X1 U390 ( .A(n324), .B(KEYINPUT2), .ZN(n423) );
  XOR2_X1 U391 ( .A(G85GAT), .B(n423), .Z(n326) );
  XNOR2_X1 U392 ( .A(G29GAT), .B(G162GAT), .ZN(n325) );
  XNOR2_X1 U393 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U394 ( .A(n328), .B(n327), .Z(n333) );
  XOR2_X1 U395 ( .A(KEYINPUT83), .B(KEYINPUT0), .Z(n330) );
  XNOR2_X1 U396 ( .A(KEYINPUT84), .B(G127GAT), .ZN(n329) );
  XNOR2_X1 U397 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U398 ( .A(G113GAT), .B(n331), .Z(n429) );
  XNOR2_X1 U399 ( .A(n429), .B(G134GAT), .ZN(n332) );
  XOR2_X1 U400 ( .A(n333), .B(n332), .Z(n490) );
  INV_X1 U401 ( .A(n490), .ZN(n527) );
  XNOR2_X1 U402 ( .A(KEYINPUT112), .B(KEYINPUT46), .ZN(n365) );
  XOR2_X1 U403 ( .A(KEYINPUT67), .B(KEYINPUT71), .Z(n335) );
  XNOR2_X1 U404 ( .A(KEYINPUT29), .B(KEYINPUT30), .ZN(n334) );
  XNOR2_X1 U405 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U406 ( .A(n337), .B(n336), .ZN(n346) );
  XOR2_X1 U407 ( .A(G141GAT), .B(G22GAT), .Z(n415) );
  XOR2_X1 U408 ( .A(KEYINPUT69), .B(KEYINPUT70), .Z(n339) );
  XNOR2_X1 U409 ( .A(G15GAT), .B(G1GAT), .ZN(n338) );
  XNOR2_X1 U410 ( .A(n339), .B(n338), .ZN(n366) );
  XOR2_X1 U411 ( .A(n415), .B(n366), .Z(n341) );
  NAND2_X1 U412 ( .A1(G229GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U413 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U414 ( .A(G169GAT), .B(G8GAT), .Z(n404) );
  XOR2_X1 U415 ( .A(n342), .B(n404), .Z(n344) );
  XNOR2_X1 U416 ( .A(G197GAT), .B(G113GAT), .ZN(n343) );
  XNOR2_X1 U417 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U418 ( .A(n346), .B(n345), .ZN(n579) );
  XOR2_X1 U419 ( .A(G120GAT), .B(G71GAT), .Z(n438) );
  INV_X1 U420 ( .A(G148GAT), .ZN(n347) );
  NAND2_X1 U421 ( .A1(G78GAT), .A2(n347), .ZN(n350) );
  INV_X1 U422 ( .A(G78GAT), .ZN(n348) );
  NAND2_X1 U423 ( .A1(n348), .A2(G148GAT), .ZN(n349) );
  NAND2_X1 U424 ( .A1(n350), .A2(n349), .ZN(n352) );
  XNOR2_X1 U425 ( .A(KEYINPUT75), .B(G204GAT), .ZN(n351) );
  XNOR2_X1 U426 ( .A(n352), .B(n351), .ZN(n424) );
  XNOR2_X1 U427 ( .A(n354), .B(KEYINPUT76), .ZN(n361) );
  XOR2_X1 U428 ( .A(n355), .B(KEYINPUT74), .Z(n359) );
  XOR2_X1 U429 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n357) );
  XNOR2_X1 U430 ( .A(KEYINPUT33), .B(KEYINPUT73), .ZN(n356) );
  XOR2_X1 U431 ( .A(n357), .B(n356), .Z(n358) );
  XOR2_X1 U432 ( .A(G57GAT), .B(KEYINPUT13), .Z(n377) );
  XOR2_X1 U433 ( .A(G176GAT), .B(G64GAT), .Z(n403) );
  XNOR2_X1 U434 ( .A(n377), .B(n403), .ZN(n362) );
  XNOR2_X1 U435 ( .A(n363), .B(n362), .ZN(n584) );
  XNOR2_X1 U436 ( .A(KEYINPUT41), .B(n584), .ZN(n568) );
  AND2_X1 U437 ( .A1(n579), .A2(n568), .ZN(n364) );
  XNOR2_X1 U438 ( .A(n365), .B(n364), .ZN(n386) );
  XOR2_X1 U439 ( .A(n366), .B(KEYINPUT12), .Z(n368) );
  NAND2_X1 U440 ( .A1(G231GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U441 ( .A(n368), .B(n367), .ZN(n384) );
  XOR2_X1 U442 ( .A(KEYINPUT81), .B(G64GAT), .Z(n370) );
  XNOR2_X1 U443 ( .A(G8GAT), .B(G127GAT), .ZN(n369) );
  XNOR2_X1 U444 ( .A(n370), .B(n369), .ZN(n374) );
  XOR2_X1 U445 ( .A(KEYINPUT80), .B(KEYINPUT79), .Z(n372) );
  XNOR2_X1 U446 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n371) );
  XNOR2_X1 U447 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U448 ( .A(n374), .B(n373), .ZN(n382) );
  XOR2_X1 U449 ( .A(G211GAT), .B(G78GAT), .Z(n376) );
  XNOR2_X1 U450 ( .A(G183GAT), .B(G71GAT), .ZN(n375) );
  XNOR2_X1 U451 ( .A(n376), .B(n375), .ZN(n378) );
  XOR2_X1 U452 ( .A(n378), .B(n377), .Z(n380) );
  XNOR2_X1 U453 ( .A(G22GAT), .B(G155GAT), .ZN(n379) );
  XNOR2_X1 U454 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U455 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U456 ( .A(n384), .B(n383), .Z(n588) );
  OR2_X1 U457 ( .A1(n561), .A2(n588), .ZN(n385) );
  XNOR2_X1 U458 ( .A(KEYINPUT113), .B(n387), .ZN(n388) );
  XNOR2_X1 U459 ( .A(n388), .B(KEYINPUT47), .ZN(n394) );
  INV_X1 U460 ( .A(KEYINPUT45), .ZN(n390) );
  INV_X1 U461 ( .A(n588), .ZN(n465) );
  NOR2_X1 U462 ( .A1(n465), .A2(n467), .ZN(n389) );
  XNOR2_X1 U463 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U464 ( .A(n579), .B(KEYINPUT72), .ZN(n565) );
  NOR2_X1 U465 ( .A1(n391), .A2(n565), .ZN(n392) );
  NAND2_X1 U466 ( .A1(n392), .A2(n584), .ZN(n393) );
  NAND2_X1 U467 ( .A1(n394), .A2(n393), .ZN(n396) );
  XOR2_X1 U468 ( .A(KEYINPUT114), .B(KEYINPUT48), .Z(n395) );
  XNOR2_X1 U469 ( .A(n396), .B(n395), .ZN(n554) );
  XNOR2_X1 U470 ( .A(KEYINPUT18), .B(KEYINPUT86), .ZN(n397) );
  XNOR2_X1 U471 ( .A(n397), .B(G183GAT), .ZN(n398) );
  XOR2_X1 U472 ( .A(n398), .B(KEYINPUT87), .Z(n400) );
  XNOR2_X1 U473 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n399) );
  XNOR2_X1 U474 ( .A(n400), .B(n399), .ZN(n430) );
  XNOR2_X1 U475 ( .A(G197GAT), .B(KEYINPUT89), .ZN(n401) );
  XNOR2_X1 U476 ( .A(n294), .B(n401), .ZN(n416) );
  NAND2_X1 U477 ( .A1(G226GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U478 ( .A(n292), .B(n402), .ZN(n409) );
  XNOR2_X1 U479 ( .A(n404), .B(n403), .ZN(n407) );
  XOR2_X1 U480 ( .A(G92GAT), .B(G218GAT), .Z(n406) );
  XNOR2_X1 U481 ( .A(G36GAT), .B(G190GAT), .ZN(n405) );
  XOR2_X1 U482 ( .A(n430), .B(n410), .Z(n529) );
  INV_X1 U483 ( .A(n529), .ZN(n494) );
  XNOR2_X1 U484 ( .A(n412), .B(KEYINPUT54), .ZN(n413) );
  NOR2_X1 U485 ( .A1(n527), .A2(n413), .ZN(n475) );
  XNOR2_X1 U486 ( .A(n415), .B(n414), .ZN(n428) );
  XOR2_X1 U487 ( .A(n416), .B(KEYINPUT22), .Z(n418) );
  NAND2_X1 U488 ( .A1(G228GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U489 ( .A(n418), .B(n417), .ZN(n422) );
  XOR2_X1 U490 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n420) );
  XNOR2_X1 U491 ( .A(G50GAT), .B(G106GAT), .ZN(n419) );
  XNOR2_X1 U492 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U493 ( .A(n422), .B(n421), .Z(n426) );
  XNOR2_X1 U494 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U495 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U496 ( .A(n428), .B(n427), .ZN(n476) );
  XNOR2_X1 U497 ( .A(n430), .B(n429), .ZN(n445) );
  XOR2_X1 U498 ( .A(KEYINPUT85), .B(KEYINPUT20), .Z(n432) );
  XNOR2_X1 U499 ( .A(G43GAT), .B(G99GAT), .ZN(n431) );
  XNOR2_X1 U500 ( .A(n432), .B(n431), .ZN(n436) );
  XOR2_X1 U501 ( .A(G176GAT), .B(KEYINPUT88), .Z(n434) );
  XNOR2_X1 U502 ( .A(G169GAT), .B(KEYINPUT64), .ZN(n433) );
  XNOR2_X1 U503 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U504 ( .A(n436), .B(n435), .Z(n443) );
  XOR2_X1 U505 ( .A(n438), .B(n437), .Z(n440) );
  NAND2_X1 U506 ( .A1(G227GAT), .A2(G233GAT), .ZN(n439) );
  XNOR2_X1 U507 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U508 ( .A(G15GAT), .B(n441), .ZN(n442) );
  XNOR2_X1 U509 ( .A(n443), .B(n442), .ZN(n444) );
  NOR2_X1 U510 ( .A1(n476), .A2(n531), .ZN(n447) );
  XNOR2_X1 U511 ( .A(KEYINPUT26), .B(KEYINPUT94), .ZN(n446) );
  XNOR2_X1 U512 ( .A(n447), .B(n446), .ZN(n552) );
  NOR2_X1 U513 ( .A1(n467), .A2(n585), .ZN(n451) );
  NAND2_X1 U514 ( .A1(n584), .A2(n565), .ZN(n482) );
  XNOR2_X1 U515 ( .A(KEYINPUT27), .B(n529), .ZN(n457) );
  NAND2_X1 U516 ( .A1(n457), .A2(n527), .ZN(n452) );
  XOR2_X1 U517 ( .A(KEYINPUT92), .B(n452), .Z(n551) );
  XOR2_X1 U518 ( .A(n476), .B(KEYINPUT28), .Z(n534) );
  INV_X1 U519 ( .A(n534), .ZN(n500) );
  NAND2_X1 U520 ( .A1(n551), .A2(n500), .ZN(n540) );
  NOR2_X1 U521 ( .A1(n531), .A2(n540), .ZN(n453) );
  XOR2_X1 U522 ( .A(KEYINPUT93), .B(n453), .Z(n463) );
  NAND2_X1 U523 ( .A1(n531), .A2(n529), .ZN(n454) );
  NAND2_X1 U524 ( .A1(n454), .A2(n476), .ZN(n455) );
  XNOR2_X1 U525 ( .A(n455), .B(KEYINPUT25), .ZN(n456) );
  XNOR2_X1 U526 ( .A(KEYINPUT95), .B(n456), .ZN(n459) );
  NAND2_X1 U527 ( .A1(n457), .A2(n552), .ZN(n458) );
  NAND2_X1 U528 ( .A1(n459), .A2(n458), .ZN(n460) );
  NAND2_X1 U529 ( .A1(n490), .A2(n460), .ZN(n461) );
  XOR2_X1 U530 ( .A(KEYINPUT96), .B(n461), .Z(n462) );
  NAND2_X1 U531 ( .A1(n465), .A2(n487), .ZN(n466) );
  XNOR2_X1 U532 ( .A(KEYINPUT37), .B(KEYINPUT102), .ZN(n468) );
  XNOR2_X1 U533 ( .A(n469), .B(n468), .ZN(n525) );
  NOR2_X1 U534 ( .A1(n482), .A2(n525), .ZN(n470) );
  XNOR2_X1 U535 ( .A(n470), .B(KEYINPUT38), .ZN(n507) );
  NAND2_X1 U536 ( .A1(n507), .A2(n531), .ZN(n474) );
  XOR2_X1 U537 ( .A(KEYINPUT40), .B(KEYINPUT104), .Z(n472) );
  INV_X1 U538 ( .A(n531), .ZN(n538) );
  AND2_X1 U539 ( .A1(n476), .A2(n475), .ZN(n477) );
  XNOR2_X1 U540 ( .A(KEYINPUT55), .B(n477), .ZN(n478) );
  NAND2_X1 U541 ( .A1(n575), .A2(n588), .ZN(n481) );
  XOR2_X1 U542 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n479) );
  INV_X1 U543 ( .A(n482), .ZN(n489) );
  XOR2_X1 U544 ( .A(KEYINPUT82), .B(KEYINPUT16), .Z(n485) );
  NAND2_X1 U545 ( .A1(n483), .A2(n588), .ZN(n484) );
  XNOR2_X1 U546 ( .A(n485), .B(n484), .ZN(n486) );
  NAND2_X1 U547 ( .A1(n487), .A2(n486), .ZN(n488) );
  XOR2_X1 U548 ( .A(KEYINPUT98), .B(n488), .Z(n513) );
  NAND2_X1 U549 ( .A1(n489), .A2(n513), .ZN(n499) );
  NOR2_X1 U550 ( .A1(n490), .A2(n499), .ZN(n492) );
  XNOR2_X1 U551 ( .A(KEYINPUT99), .B(KEYINPUT34), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U553 ( .A(G1GAT), .B(n493), .ZN(G1324GAT) );
  NOR2_X1 U554 ( .A1(n494), .A2(n499), .ZN(n495) );
  XOR2_X1 U555 ( .A(KEYINPUT100), .B(n495), .Z(n496) );
  XNOR2_X1 U556 ( .A(G8GAT), .B(n496), .ZN(G1325GAT) );
  NOR2_X1 U557 ( .A1(n538), .A2(n499), .ZN(n498) );
  XNOR2_X1 U558 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n498), .B(n497), .ZN(G1326GAT) );
  NOR2_X1 U560 ( .A1(n500), .A2(n499), .ZN(n502) );
  XNOR2_X1 U561 ( .A(G22GAT), .B(KEYINPUT101), .ZN(n501) );
  XNOR2_X1 U562 ( .A(n502), .B(n501), .ZN(G1327GAT) );
  XOR2_X1 U563 ( .A(G29GAT), .B(KEYINPUT39), .Z(n504) );
  NAND2_X1 U564 ( .A1(n527), .A2(n507), .ZN(n503) );
  XNOR2_X1 U565 ( .A(n504), .B(n503), .ZN(G1328GAT) );
  XOR2_X1 U566 ( .A(G36GAT), .B(KEYINPUT103), .Z(n506) );
  NAND2_X1 U567 ( .A1(n529), .A2(n507), .ZN(n505) );
  XNOR2_X1 U568 ( .A(n506), .B(n505), .ZN(G1329GAT) );
  XOR2_X1 U569 ( .A(G50GAT), .B(KEYINPUT105), .Z(n509) );
  NAND2_X1 U570 ( .A1(n534), .A2(n507), .ZN(n508) );
  XNOR2_X1 U571 ( .A(n509), .B(n508), .ZN(G1331GAT) );
  XOR2_X1 U572 ( .A(KEYINPUT108), .B(KEYINPUT42), .Z(n516) );
  INV_X1 U573 ( .A(n568), .ZN(n510) );
  NOR2_X1 U574 ( .A1(n510), .A2(n579), .ZN(n511) );
  XOR2_X1 U575 ( .A(n511), .B(KEYINPUT106), .Z(n524) );
  INV_X1 U576 ( .A(n524), .ZN(n512) );
  NAND2_X1 U577 ( .A1(n513), .A2(n512), .ZN(n514) );
  XNOR2_X1 U578 ( .A(n514), .B(KEYINPUT107), .ZN(n520) );
  NAND2_X1 U579 ( .A1(n520), .A2(n527), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n516), .B(n515), .ZN(n517) );
  XOR2_X1 U581 ( .A(G57GAT), .B(n517), .Z(G1332GAT) );
  NAND2_X1 U582 ( .A1(n520), .A2(n529), .ZN(n518) );
  XNOR2_X1 U583 ( .A(n518), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U584 ( .A1(n531), .A2(n520), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n519), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n522) );
  NAND2_X1 U587 ( .A1(n520), .A2(n534), .ZN(n521) );
  XNOR2_X1 U588 ( .A(n522), .B(n521), .ZN(n523) );
  XOR2_X1 U589 ( .A(G78GAT), .B(n523), .Z(G1335GAT) );
  NOR2_X1 U590 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U591 ( .A(KEYINPUT110), .B(n526), .ZN(n533) );
  NAND2_X1 U592 ( .A1(n533), .A2(n527), .ZN(n528) );
  XNOR2_X1 U593 ( .A(n528), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U594 ( .A1(n533), .A2(n529), .ZN(n530) );
  XNOR2_X1 U595 ( .A(n530), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U596 ( .A1(n533), .A2(n531), .ZN(n532) );
  XNOR2_X1 U597 ( .A(n532), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT44), .B(KEYINPUT111), .Z(n536) );
  NAND2_X1 U599 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U600 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U601 ( .A(G106GAT), .B(n537), .ZN(G1339GAT) );
  OR2_X1 U602 ( .A1(n538), .A2(n554), .ZN(n539) );
  NOR2_X1 U603 ( .A1(n540), .A2(n539), .ZN(n548) );
  NAND2_X1 U604 ( .A1(n548), .A2(n565), .ZN(n541) );
  XNOR2_X1 U605 ( .A(G113GAT), .B(n541), .ZN(G1340GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT49), .B(KEYINPUT115), .Z(n543) );
  NAND2_X1 U607 ( .A1(n548), .A2(n568), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n543), .B(n542), .ZN(n544) );
  XOR2_X1 U609 ( .A(G120GAT), .B(n544), .Z(G1341GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n546) );
  NAND2_X1 U611 ( .A1(n548), .A2(n588), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U613 ( .A(G127GAT), .B(n547), .Z(G1342GAT) );
  XOR2_X1 U614 ( .A(G134GAT), .B(KEYINPUT51), .Z(n550) );
  NAND2_X1 U615 ( .A1(n548), .A2(n576), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(G1343GAT) );
  NAND2_X1 U617 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X1 U618 ( .A1(n554), .A2(n553), .ZN(n562) );
  NAND2_X1 U619 ( .A1(n562), .A2(n579), .ZN(n555) );
  XNOR2_X1 U620 ( .A(n555), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT117), .B(KEYINPUT52), .Z(n557) );
  NAND2_X1 U622 ( .A1(n562), .A2(n568), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(n559) );
  XOR2_X1 U624 ( .A(G148GAT), .B(KEYINPUT53), .Z(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(G1345GAT) );
  NAND2_X1 U626 ( .A1(n562), .A2(n588), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n560), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(KEYINPUT118), .ZN(n564) );
  XNOR2_X1 U630 ( .A(G162GAT), .B(n564), .ZN(G1347GAT) );
  XOR2_X1 U631 ( .A(G169GAT), .B(KEYINPUT119), .Z(n567) );
  NAND2_X1 U632 ( .A1(n575), .A2(n565), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(G1348GAT) );
  NAND2_X1 U634 ( .A1(n568), .A2(n575), .ZN(n574) );
  XOR2_X1 U635 ( .A(KEYINPUT122), .B(KEYINPUT121), .Z(n570) );
  XNOR2_X1 U636 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n570), .B(n569), .ZN(n572) );
  XOR2_X1 U638 ( .A(G176GAT), .B(KEYINPUT120), .Z(n571) );
  XNOR2_X1 U639 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(G1349GAT) );
  NAND2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n577), .B(KEYINPUT58), .ZN(n578) );
  XNOR2_X1 U643 ( .A(G190GAT), .B(n578), .ZN(G1351GAT) );
  INV_X1 U644 ( .A(n585), .ZN(n589) );
  NAND2_X1 U645 ( .A1(n589), .A2(n579), .ZN(n583) );
  XOR2_X1 U646 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n581) );
  XNOR2_X1 U647 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n580) );
  XNOR2_X1 U648 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n583), .B(n582), .ZN(G1352GAT) );
  XOR2_X1 U650 ( .A(G204GAT), .B(KEYINPUT61), .Z(n587) );
  OR2_X1 U651 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(G1353GAT) );
  XOR2_X1 U653 ( .A(G211GAT), .B(KEYINPUT127), .Z(n591) );
  NAND2_X1 U654 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n591), .B(n590), .ZN(G1354GAT) );
endmodule

