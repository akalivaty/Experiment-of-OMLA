//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 1 0 0 1 1 1 0 1 0 1 0 1 0 0 0 0 0 1 0 0 1 0 1 0 0 1 1 0 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 1 1 1 1 0 1 0 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:11 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n578, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n594, new_n595,
    new_n596, new_n599, new_n600, new_n601, new_n602, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n631, new_n633,
    new_n634, new_n635, new_n636, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1169, new_n1170, new_n1171, new_n1173,
    new_n1174, new_n1175;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT65), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT66), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT67), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G125), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n462), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n463), .A2(G137), .A3(new_n462), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n466), .A2(new_n471), .ZN(G160));
  XOR2_X1   g047(.A(KEYINPUT3), .B(G2104), .Z(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(new_n462), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  XNOR2_X1  g050(.A(new_n475), .B(KEYINPUT69), .ZN(new_n476));
  OR2_X1    g051(.A1(G100), .A2(G2105), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n477), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n478));
  AND2_X1   g053(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n473), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT68), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  INV_X1    g059(.A(new_n469), .ZN(new_n485));
  INV_X1    g060(.A(G102), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(G114), .A2(G2104), .ZN(new_n488));
  INV_X1    g063(.A(G126), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n488), .B1(new_n473), .B2(new_n489), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n487), .B1(new_n490), .B2(G2105), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n463), .A2(G138), .A3(new_n462), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n463), .A2(new_n494), .A3(G138), .A4(new_n462), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n491), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  NAND2_X1  g073(.A1(G75), .A2(G543), .ZN(new_n499));
  INV_X1    g074(.A(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT5), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(G62), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n499), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(G50), .A2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G88), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n508), .B1(new_n504), .B2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(KEYINPUT6), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT6), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n510), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n507), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT70), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n507), .A2(new_n517), .A3(KEYINPUT70), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(G166));
  INV_X1    g097(.A(KEYINPUT74), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT71), .ZN(new_n524));
  AND3_X1   g099(.A1(new_n501), .A2(new_n503), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n524), .B1(new_n501), .B2(new_n503), .ZN(new_n526));
  OAI21_X1  g101(.A(G63), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(G76), .A2(G543), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT7), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n511), .B1(new_n527), .B2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT72), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n513), .A2(G651), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n511), .A2(KEYINPUT6), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n512), .A2(new_n514), .A3(KEYINPUT72), .ZN(new_n537));
  NAND4_X1  g112(.A1(new_n536), .A2(G51), .A3(G543), .A4(new_n537), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n529), .B1(new_n528), .B2(new_n511), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n502), .A2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n500), .A2(KEYINPUT5), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  XNOR2_X1  g117(.A(KEYINPUT73), .B(G89), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n516), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n538), .A2(new_n539), .A3(new_n544), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n523), .B1(new_n532), .B2(new_n545), .ZN(new_n546));
  NAND4_X1  g121(.A1(new_n501), .A2(new_n503), .A3(new_n512), .A4(new_n514), .ZN(new_n547));
  XOR2_X1   g122(.A(KEYINPUT73), .B(G89), .Z(new_n548));
  OAI21_X1  g123(.A(new_n539), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AND3_X1   g124(.A1(new_n512), .A2(new_n514), .A3(KEYINPUT72), .ZN(new_n550));
  AOI21_X1  g125(.A(KEYINPUT72), .B1(new_n512), .B2(new_n514), .ZN(new_n551));
  NOR3_X1   g126(.A1(new_n550), .A2(new_n551), .A3(new_n500), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n549), .B1(new_n552), .B2(G51), .ZN(new_n553));
  INV_X1    g128(.A(G63), .ZN(new_n554));
  OAI21_X1  g129(.A(KEYINPUT71), .B1(new_n540), .B2(new_n541), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n501), .A2(new_n503), .A3(new_n524), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g132(.A(G651), .B1(new_n557), .B2(new_n530), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n553), .A2(new_n558), .A3(KEYINPUT74), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n546), .A2(new_n559), .ZN(G168));
  NAND2_X1  g135(.A1(new_n555), .A2(new_n556), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G64), .ZN(new_n562));
  NAND2_X1  g137(.A1(G77), .A2(G543), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n511), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n536), .A2(G543), .A3(new_n537), .ZN(new_n565));
  INV_X1    g140(.A(G52), .ZN(new_n566));
  INV_X1    g141(.A(G90), .ZN(new_n567));
  OAI22_X1  g142(.A1(new_n565), .A2(new_n566), .B1(new_n567), .B2(new_n547), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n564), .A2(new_n568), .ZN(G171));
  NAND2_X1  g144(.A1(new_n561), .A2(G56), .ZN(new_n570));
  NAND2_X1  g145(.A1(G68), .A2(G543), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n511), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(G43), .ZN(new_n573));
  INV_X1    g148(.A(G81), .ZN(new_n574));
  OAI22_X1  g149(.A1(new_n565), .A2(new_n573), .B1(new_n574), .B2(new_n547), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(G860), .ZN(G153));
  AND3_X1   g152(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(G36), .ZN(G176));
  NAND2_X1  g154(.A1(G1), .A2(G3), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n580), .B(KEYINPUT75), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n581), .B(KEYINPUT8), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  XOR2_X1   g158(.A(new_n583), .B(KEYINPUT76), .Z(G188));
  AOI22_X1  g159(.A1(new_n542), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n585));
  OR2_X1    g160(.A1(new_n585), .A2(new_n511), .ZN(new_n586));
  INV_X1    g161(.A(new_n547), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(G91), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n536), .A2(G53), .A3(G543), .A4(new_n537), .ZN(new_n589));
  AND2_X1   g164(.A1(new_n589), .A2(KEYINPUT9), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n589), .A2(KEYINPUT9), .ZN(new_n591));
  OAI211_X1 g166(.A(new_n586), .B(new_n588), .C1(new_n590), .C2(new_n591), .ZN(G299));
  INV_X1    g167(.A(G171), .ZN(G301));
  AND3_X1   g168(.A1(new_n546), .A2(new_n559), .A3(KEYINPUT77), .ZN(new_n594));
  AOI21_X1  g169(.A(KEYINPUT77), .B1(new_n546), .B2(new_n559), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(G286));
  INV_X1    g172(.A(G166), .ZN(G303));
  NOR2_X1   g173(.A1(new_n525), .A2(new_n526), .ZN(new_n599));
  INV_X1    g174(.A(G74), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n601), .A2(G651), .B1(G87), .B2(new_n587), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n552), .A2(G49), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(G288));
  AOI22_X1  g179(.A1(new_n542), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n605), .A2(new_n511), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n542), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n607), .A2(new_n515), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(G305));
  AND2_X1   g185(.A1(new_n561), .A2(G60), .ZN(new_n611));
  NAND2_X1  g186(.A1(G72), .A2(G543), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(G651), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n552), .A2(G47), .B1(G85), .B2(new_n587), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(new_n615), .ZN(G290));
  NAND2_X1  g191(.A1(G301), .A2(G868), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n542), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n618));
  OR2_X1    g193(.A1(new_n618), .A2(new_n511), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n552), .A2(G54), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n587), .A2(KEYINPUT10), .A3(G92), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT10), .ZN(new_n622));
  INV_X1    g197(.A(G92), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n547), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  AND3_X1   g200(.A1(new_n619), .A2(new_n620), .A3(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n617), .B1(G868), .B2(new_n626), .ZN(G284));
  OAI21_X1  g202(.A(new_n617), .B1(G868), .B2(new_n626), .ZN(G321));
  MUX2_X1   g203(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g204(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g205(.A(G559), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n626), .B1(new_n631), .B2(G860), .ZN(G148));
  NAND2_X1  g207(.A1(new_n626), .A2(new_n631), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(G868), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n634), .A2(KEYINPUT78), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(KEYINPUT78), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n635), .B(new_n636), .C1(G868), .C2(new_n576), .ZN(G323));
  XNOR2_X1  g212(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g213(.A1(new_n463), .A2(new_n469), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT12), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT13), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2100), .ZN(new_n642));
  AOI22_X1  g217(.A1(G123), .A2(new_n474), .B1(new_n480), .B2(G135), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n462), .A2(G111), .ZN(new_n644));
  INV_X1    g219(.A(KEYINPUT79), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n468), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OAI221_X1 g221(.A(new_n646), .B1(new_n645), .B2(new_n644), .C1(G99), .C2(G2105), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n643), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT80), .B(G2096), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n642), .A2(new_n650), .ZN(G156));
  XNOR2_X1  g226(.A(G2451), .B(G2454), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT16), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G1341), .B(G1348), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2427), .B(G2430), .ZN(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT81), .B(G2438), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(KEYINPUT15), .B(G2435), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n662), .A2(KEYINPUT14), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n657), .B(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n664), .A2(G14), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT82), .ZN(G401));
  XNOR2_X1  g241(.A(G2072), .B(G2078), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT17), .Z(new_n668));
  XOR2_X1   g243(.A(G2067), .B(G2678), .Z(new_n669));
  XOR2_X1   g244(.A(G2084), .B(G2090), .Z(new_n670));
  NAND3_X1  g245(.A1(new_n668), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT83), .Z(new_n672));
  NOR2_X1   g247(.A1(new_n668), .A2(new_n669), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n673), .A2(new_n670), .ZN(new_n674));
  INV_X1    g249(.A(new_n669), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n674), .B1(new_n675), .B2(new_n667), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n675), .A2(new_n667), .A3(new_n670), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT18), .Z(new_n678));
  NAND3_X1  g253(.A1(new_n672), .A2(new_n676), .A3(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(G2096), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(G2100), .ZN(G227));
  XNOR2_X1  g256(.A(G1971), .B(G1976), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT84), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n683), .A2(KEYINPUT19), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n683), .A2(KEYINPUT19), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(G1956), .B(G2474), .Z(new_n687));
  XOR2_X1   g262(.A(G1961), .B(G1966), .Z(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n687), .A2(new_n688), .ZN(new_n691));
  OR3_X1    g266(.A1(new_n686), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n689), .B1(new_n684), .B2(new_n685), .ZN(new_n693));
  XOR2_X1   g268(.A(KEYINPUT85), .B(KEYINPUT20), .Z(new_n694));
  AOI22_X1  g269(.A1(new_n693), .A2(new_n694), .B1(new_n686), .B2(new_n691), .ZN(new_n695));
  OAI211_X1 g270(.A(new_n692), .B(new_n695), .C1(new_n693), .C2(new_n694), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT86), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1991), .B(G1996), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n698), .B(new_n699), .Z(new_n700));
  NOR2_X1   g275(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1981), .B(G1986), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n697), .A2(new_n700), .ZN(new_n704));
  AND3_X1   g279(.A1(new_n702), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n703), .B1(new_n702), .B2(new_n704), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n705), .A2(new_n706), .ZN(G229));
  INV_X1    g282(.A(KEYINPUT87), .ZN(new_n708));
  INV_X1    g283(.A(G29), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n709), .A2(G25), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n474), .A2(G119), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT88), .Z(new_n712));
  OR2_X1    g287(.A1(G95), .A2(G2105), .ZN(new_n713));
  OAI211_X1 g288(.A(new_n713), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n480), .A2(G131), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n712), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  AOI211_X1 g291(.A(new_n708), .B(new_n710), .C1(new_n716), .C2(G29), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(new_n708), .B2(new_n710), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT35), .B(G1991), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT89), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n718), .B(new_n720), .ZN(new_n721));
  NOR2_X1   g296(.A1(G16), .A2(G23), .ZN(new_n722));
  INV_X1    g297(.A(G288), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n722), .B1(new_n723), .B2(G16), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT33), .B(G1976), .Z(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G22), .ZN(new_n727));
  OR3_X1    g302(.A1(new_n727), .A2(KEYINPUT91), .A3(G16), .ZN(new_n728));
  OAI21_X1  g303(.A(KEYINPUT91), .B1(new_n727), .B2(G16), .ZN(new_n729));
  INV_X1    g304(.A(G16), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n728), .B(new_n729), .C1(G166), .C2(new_n730), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n731), .A2(G1971), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(G1971), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n730), .A2(G6), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(new_n609), .B2(new_n730), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT32), .B(G1981), .Z(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n732), .A2(new_n733), .A3(new_n737), .ZN(new_n738));
  OR3_X1    g313(.A1(new_n726), .A2(new_n738), .A3(KEYINPUT34), .ZN(new_n739));
  OAI21_X1  g314(.A(KEYINPUT34), .B1(new_n726), .B2(new_n738), .ZN(new_n740));
  NOR2_X1   g315(.A1(G16), .A2(G24), .ZN(new_n741));
  XOR2_X1   g316(.A(G290), .B(KEYINPUT90), .Z(new_n742));
  AOI21_X1  g317(.A(new_n741), .B1(new_n742), .B2(G16), .ZN(new_n743));
  INV_X1    g318(.A(G1986), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND4_X1  g320(.A1(new_n721), .A2(new_n739), .A3(new_n740), .A4(new_n745), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT36), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT23), .ZN(new_n748));
  AND2_X1   g323(.A1(new_n730), .A2(G20), .ZN(new_n749));
  AOI211_X1 g324(.A(new_n748), .B(new_n749), .C1(G299), .C2(G16), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n748), .B2(new_n749), .ZN(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT100), .B(G1956), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n626), .A2(new_n730), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G4), .B2(new_n730), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT92), .B(G1348), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT93), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(G2084), .ZN(new_n759));
  OAI21_X1  g334(.A(G29), .B1(new_n466), .B2(new_n471), .ZN(new_n760));
  OR2_X1    g335(.A1(KEYINPUT24), .A2(G34), .ZN(new_n761));
  NAND2_X1  g336(.A1(KEYINPUT24), .A2(G34), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n761), .A2(new_n709), .A3(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n759), .B1(new_n760), .B2(new_n763), .ZN(new_n764));
  AND3_X1   g339(.A1(new_n760), .A2(new_n759), .A3(new_n763), .ZN(new_n765));
  AOI22_X1  g340(.A1(G129), .A2(new_n474), .B1(new_n480), .B2(G141), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT95), .B(KEYINPUT26), .Z(new_n767));
  NAND3_X1  g342(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n469), .A2(G105), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n766), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n772), .A2(G29), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G29), .B2(G32), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT27), .B(G1996), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT96), .Z(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  AOI211_X1 g352(.A(new_n764), .B(new_n765), .C1(new_n774), .C2(new_n777), .ZN(new_n778));
  NOR2_X1   g353(.A1(G5), .A2(G16), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G171), .B2(G16), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n780), .A2(G1961), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n755), .A2(new_n757), .ZN(new_n782));
  NAND4_X1  g357(.A1(new_n758), .A2(new_n778), .A3(new_n781), .A4(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(new_n774), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n783), .B1(new_n776), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n469), .A2(G103), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT25), .Z(new_n787));
  NAND2_X1  g362(.A1(new_n480), .A2(G139), .ZN(new_n788));
  AOI22_X1  g363(.A1(new_n463), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n789));
  OAI211_X1 g364(.A(new_n787), .B(new_n788), .C1(new_n462), .C2(new_n789), .ZN(new_n790));
  MUX2_X1   g365(.A(G33), .B(new_n790), .S(G29), .Z(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(G2072), .Z(new_n792));
  NAND2_X1  g367(.A1(new_n730), .A2(G19), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n576), .B2(new_n730), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G1341), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n709), .A2(G27), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G164), .B2(new_n709), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G2078), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT94), .B(KEYINPUT28), .Z(new_n799));
  NAND2_X1  g374(.A1(new_n709), .A2(G26), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n480), .A2(G140), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n474), .A2(G128), .ZN(new_n803));
  OR2_X1    g378(.A1(G104), .A2(G2105), .ZN(new_n804));
  OAI211_X1 g379(.A(new_n804), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n802), .A2(new_n803), .A3(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n801), .B1(new_n807), .B2(new_n709), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(G2067), .ZN(new_n809));
  NOR3_X1   g384(.A1(new_n795), .A2(new_n798), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n709), .A2(G35), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(G162), .B2(new_n709), .ZN(new_n812));
  XOR2_X1   g387(.A(KEYINPUT29), .B(G2090), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n785), .A2(new_n792), .A3(new_n810), .A4(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT30), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n709), .B1(new_n816), .B2(G28), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT97), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n816), .A2(G28), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n817), .A2(new_n818), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n819), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(new_n648), .B2(new_n709), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n780), .A2(G1961), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n824), .A2(KEYINPUT98), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(KEYINPUT98), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n823), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(KEYINPUT31), .B(G11), .ZN(new_n828));
  NOR2_X1   g403(.A1(G16), .A2(G21), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(G168), .B2(G16), .ZN(new_n830));
  INV_X1    g405(.A(G1966), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n827), .A2(new_n828), .A3(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT99), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n833), .A2(new_n834), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n815), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n747), .A2(new_n753), .A3(new_n837), .ZN(G150));
  INV_X1    g413(.A(G150), .ZN(G311));
  INV_X1    g414(.A(G67), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n599), .A2(new_n840), .ZN(new_n841));
  AND2_X1   g416(.A1(G80), .A2(G543), .ZN(new_n842));
  OAI21_X1  g417(.A(G651), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n587), .A2(G93), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n536), .A2(G55), .A3(G543), .A4(new_n537), .ZN(new_n845));
  AOI21_X1  g420(.A(KEYINPUT101), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  AND3_X1   g421(.A1(new_n844), .A2(new_n845), .A3(KEYINPUT101), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n843), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(G860), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(KEYINPUT37), .Z(new_n850));
  XNOR2_X1  g425(.A(new_n848), .B(new_n576), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT38), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n626), .A2(G559), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(KEYINPUT39), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n855), .B(KEYINPUT103), .Z(new_n856));
  INV_X1    g431(.A(KEYINPUT102), .ZN(new_n857));
  OR3_X1    g432(.A1(new_n854), .A2(new_n857), .A3(KEYINPUT39), .ZN(new_n858));
  INV_X1    g433(.A(G860), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n857), .B1(new_n854), .B2(KEYINPUT39), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n850), .B1(new_n856), .B2(new_n861), .ZN(G145));
  NAND2_X1  g437(.A1(new_n790), .A2(KEYINPUT104), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n771), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(new_n640), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n648), .B(G160), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(new_n716), .ZN(new_n867));
  OR2_X1    g442(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n865), .A2(new_n867), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(G2104), .B1(new_n462), .B2(G118), .ZN(new_n871));
  INV_X1    g446(.A(G106), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n871), .B1(new_n872), .B2(new_n462), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n474), .A2(G130), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n874), .B(KEYINPUT105), .Z(new_n875));
  AOI211_X1 g450(.A(new_n873), .B(new_n875), .C1(G142), .C2(new_n480), .ZN(new_n876));
  AND2_X1   g451(.A1(new_n876), .A2(new_n483), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n876), .A2(new_n483), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n807), .B(new_n497), .ZN(new_n879));
  OR3_X1    g454(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n879), .B1(new_n877), .B2(new_n878), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n870), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(KEYINPUT106), .B(G37), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n868), .A2(new_n880), .A3(new_n881), .A4(new_n869), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(KEYINPUT40), .ZN(G395));
  OR2_X1    g462(.A1(new_n572), .A2(new_n575), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n848), .B(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(new_n633), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT107), .ZN(new_n891));
  NAND2_X1  g466(.A1(G299), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n550), .A2(new_n551), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT9), .ZN(new_n894));
  NAND4_X1  g469(.A1(new_n893), .A2(new_n894), .A3(G53), .A4(G543), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n589), .A2(KEYINPUT9), .ZN(new_n896));
  AOI22_X1  g471(.A1(new_n895), .A2(new_n896), .B1(G91), .B2(new_n587), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n897), .A2(KEYINPUT107), .A3(new_n586), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n892), .A2(new_n626), .A3(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT41), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n619), .A2(new_n625), .A3(new_n620), .ZN(new_n901));
  NAND3_X1  g476(.A1(G299), .A2(new_n891), .A3(new_n901), .ZN(new_n902));
  AND3_X1   g477(.A1(new_n899), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n900), .B1(new_n899), .B2(new_n902), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OR2_X1    g480(.A1(new_n890), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n899), .A2(KEYINPUT108), .A3(new_n902), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT108), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n626), .B1(G299), .B2(new_n891), .ZN(new_n909));
  AOI21_X1  g484(.A(KEYINPUT107), .B1(new_n897), .B2(new_n586), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n902), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n908), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n890), .A2(new_n907), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n906), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(KEYINPUT42), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n723), .A2(G166), .ZN(new_n917));
  NAND2_X1  g492(.A1(G303), .A2(G288), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n917), .A2(new_n918), .A3(G305), .ZN(new_n919));
  AOI21_X1  g494(.A(G305), .B1(new_n917), .B2(new_n918), .ZN(new_n920));
  OAI21_X1  g495(.A(G290), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n917), .A2(new_n918), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(new_n609), .ZN(new_n923));
  INV_X1    g498(.A(G290), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n917), .A2(new_n918), .A3(G305), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n921), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT42), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n906), .A2(new_n928), .A3(new_n914), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n916), .A2(new_n927), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n927), .B1(new_n916), .B2(new_n929), .ZN(new_n931));
  OAI21_X1  g506(.A(G868), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n848), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n932), .B1(G868), .B2(new_n933), .ZN(G295));
  OAI21_X1  g509(.A(new_n932), .B1(G868), .B2(new_n933), .ZN(G331));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT110), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT77), .ZN(new_n938));
  NOR3_X1   g513(.A1(new_n532), .A2(new_n545), .A3(new_n523), .ZN(new_n939));
  AOI21_X1  g514(.A(KEYINPUT74), .B1(new_n553), .B2(new_n558), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n546), .A2(new_n559), .A3(KEYINPUT77), .ZN(new_n942));
  AOI21_X1  g517(.A(G301), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(G168), .A2(G301), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n889), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(G171), .B1(new_n594), .B2(new_n595), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n947), .A2(new_n851), .A3(new_n944), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n937), .B1(new_n949), .B2(new_n905), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n911), .A2(new_n912), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(KEYINPUT41), .B1(new_n911), .B2(new_n912), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n899), .A2(new_n900), .A3(new_n902), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n955), .A2(KEYINPUT110), .A3(new_n946), .A4(new_n948), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n950), .A2(new_n927), .A3(new_n952), .A4(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n913), .A2(new_n907), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n949), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n921), .A2(new_n926), .ZN(new_n960));
  OAI211_X1 g535(.A(new_n946), .B(new_n948), .C1(KEYINPUT111), .C2(new_n903), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT111), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n953), .B1(new_n962), .B2(new_n954), .ZN(new_n963));
  OAI211_X1 g538(.A(new_n959), .B(new_n960), .C1(new_n961), .C2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n957), .A2(new_n884), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n950), .A2(new_n952), .A3(new_n956), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(new_n960), .ZN(new_n968));
  INV_X1    g543(.A(G37), .ZN(new_n969));
  XNOR2_X1  g544(.A(KEYINPUT109), .B(KEYINPUT43), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n968), .A2(new_n969), .A3(new_n957), .A4(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n936), .B1(new_n966), .B2(new_n972), .ZN(new_n973));
  AND4_X1   g548(.A1(new_n884), .A2(new_n957), .A3(new_n964), .A4(new_n971), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n968), .A2(new_n969), .A3(new_n957), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n974), .B1(new_n970), .B2(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n973), .B1(new_n936), .B2(new_n976), .ZN(G397));
  INV_X1    g552(.A(G40), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n466), .A2(new_n471), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(G1384), .B1(new_n491), .B2(new_n496), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n980), .A2(KEYINPUT50), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT50), .ZN(new_n982));
  AOI211_X1 g557(.A(new_n982), .B(G1384), .C1(new_n491), .C2(new_n496), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n979), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G1956), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n895), .A2(new_n896), .ZN(new_n987));
  AOI21_X1  g562(.A(KEYINPUT57), .B1(new_n987), .B2(KEYINPUT118), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(G299), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT118), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n990), .B1(new_n895), .B2(new_n896), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n897), .B(new_n586), .C1(new_n991), .C2(KEYINPUT57), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n989), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n979), .ZN(new_n994));
  INV_X1    g569(.A(G1384), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n493), .A2(new_n495), .ZN(new_n996));
  AOI22_X1  g571(.A1(new_n463), .A2(G126), .B1(G114), .B2(G2104), .ZN(new_n997));
  OAI22_X1  g572(.A1(new_n997), .A2(new_n462), .B1(new_n486), .B2(new_n485), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n995), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT45), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n994), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g576(.A(KEYINPUT112), .B(G1384), .ZN(new_n1002));
  AOI211_X1 g577(.A(new_n1000), .B(new_n1002), .C1(new_n491), .C2(new_n496), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g579(.A(KEYINPUT56), .B(G2072), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1001), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n986), .A2(new_n993), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n756), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n984), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n497), .A2(new_n979), .A3(new_n995), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(KEYINPUT119), .ZN(new_n1011));
  INV_X1    g586(.A(G2067), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT119), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n980), .A2(new_n1013), .A3(new_n979), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1011), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1009), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1007), .A2(new_n626), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n999), .A2(new_n982), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n980), .A2(KEYINPUT50), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n994), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1006), .B1(new_n1020), .B2(G1956), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n993), .A2(KEYINPUT120), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT120), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1023), .B1(new_n989), .B2(new_n992), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1021), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n1015), .B(KEYINPUT60), .C1(new_n1020), .C2(new_n756), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(KEYINPUT123), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT123), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1009), .A2(new_n1028), .A3(KEYINPUT60), .A4(new_n1015), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1027), .A2(new_n626), .A3(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1026), .A2(KEYINPUT123), .A3(new_n901), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT60), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1016), .A2(new_n1032), .ZN(new_n1033));
  AND3_X1   g608(.A1(new_n1030), .A2(new_n1031), .A3(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1025), .A2(KEYINPUT61), .A3(new_n1007), .ZN(new_n1035));
  XOR2_X1   g610(.A(KEYINPUT122), .B(KEYINPUT61), .Z(new_n1036));
  AND3_X1   g611(.A1(new_n986), .A2(new_n993), .A3(new_n1006), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n993), .B1(new_n986), .B2(new_n1006), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1036), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  AND2_X1   g614(.A1(new_n576), .A2(KEYINPUT121), .ZN(new_n1040));
  XNOR2_X1  g615(.A(KEYINPUT58), .B(G1341), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1041), .B1(new_n1011), .B2(new_n1014), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n979), .B1(new_n980), .B2(KEYINPUT45), .ZN(new_n1043));
  NOR3_X1   g618(.A1(new_n1043), .A2(G1996), .A3(new_n1003), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1040), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(KEYINPUT59), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT59), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1047), .B(new_n1040), .C1(new_n1042), .C2(new_n1044), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1035), .A2(new_n1039), .A3(new_n1049), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1017), .B(new_n1025), .C1(new_n1034), .C2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(G8), .ZN(new_n1052));
  NOR2_X1   g627(.A1(G166), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT55), .ZN(new_n1054));
  XNOR2_X1  g629(.A(new_n1053), .B(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(G1971), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1057));
  INV_X1    g632(.A(G2090), .ZN(new_n1058));
  AOI22_X1  g633(.A1(new_n1056), .A2(new_n1057), .B1(new_n1020), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1055), .B1(new_n1059), .B2(new_n1052), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1043), .A2(new_n1003), .ZN(new_n1061));
  OAI22_X1  g636(.A1(G1971), .A2(new_n1061), .B1(new_n984), .B2(G2090), .ZN(new_n1062));
  XNOR2_X1  g637(.A(new_n1053), .B(KEYINPUT55), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1062), .A2(new_n1063), .A3(G8), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n602), .A2(G1976), .A3(new_n603), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT114), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1052), .B1(new_n980), .B2(new_n979), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n602), .A2(KEYINPUT114), .A3(G1976), .A4(new_n603), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(KEYINPUT52), .ZN(new_n1071));
  OAI21_X1  g646(.A(G1981), .B1(new_n606), .B2(KEYINPUT115), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT49), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT49), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1074), .B(G1981), .C1(new_n606), .C2(KEYINPUT115), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(G305), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1073), .A2(new_n609), .A3(new_n1075), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1077), .A2(new_n1068), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(G1976), .ZN(new_n1080));
  AOI21_X1  g655(.A(KEYINPUT52), .B1(G288), .B2(new_n1080), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1081), .A2(new_n1067), .A3(new_n1068), .A4(new_n1069), .ZN(new_n1082));
  AND3_X1   g657(.A1(new_n1071), .A2(new_n1079), .A3(new_n1082), .ZN(new_n1083));
  AND3_X1   g658(.A1(new_n1060), .A2(new_n1064), .A3(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n999), .A2(new_n1000), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n831), .B1(new_n1085), .B2(new_n1043), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1086), .B1(G2084), .B2(new_n984), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(G8), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n546), .A2(new_n559), .A3(G8), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT124), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT51), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1088), .A2(new_n1089), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1020), .A2(new_n759), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1052), .B1(new_n1095), .B2(new_n1086), .ZN(new_n1096));
  INV_X1    g671(.A(G168), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  OAI211_X1 g673(.A(G8), .B(new_n1092), .C1(new_n1087), .C2(new_n1097), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1094), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT125), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1001), .B1(new_n1000), .B2(new_n999), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1101), .B1(new_n1102), .B2(G2078), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1085), .A2(new_n1043), .ZN(new_n1104));
  INV_X1    g679(.A(G2078), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1104), .A2(KEYINPUT125), .A3(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1103), .A2(KEYINPUT53), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1061), .A2(new_n1105), .ZN(new_n1108));
  XNOR2_X1  g683(.A(KEYINPUT126), .B(KEYINPUT53), .ZN(new_n1109));
  INV_X1    g684(.A(G1961), .ZN(new_n1110));
  AOI22_X1  g685(.A1(new_n1108), .A2(new_n1109), .B1(new_n1110), .B2(new_n984), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1107), .A2(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g687(.A(G171), .B(KEYINPUT54), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1000), .B1(G164), .B2(new_n1002), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n994), .A2(G2078), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1116), .A2(new_n1004), .A3(KEYINPUT53), .A4(new_n1117), .ZN(new_n1118));
  XNOR2_X1  g693(.A(new_n1118), .B(KEYINPUT127), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1119), .A2(new_n1111), .A3(new_n1113), .ZN(new_n1120));
  AND4_X1   g695(.A1(new_n1084), .A2(new_n1100), .A3(new_n1115), .A4(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1051), .A2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1083), .A2(G8), .A3(new_n1063), .A4(new_n1062), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1079), .A2(new_n1080), .A3(new_n723), .ZN(new_n1124));
  NOR2_X1   g699(.A1(G305), .A2(G1981), .ZN(new_n1125));
  XOR2_X1   g700(.A(new_n1125), .B(KEYINPUT116), .Z(new_n1126));
  AND3_X1   g701(.A1(new_n1124), .A2(KEYINPUT117), .A3(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(KEYINPUT117), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1068), .ZN(new_n1129));
  NOR3_X1   g704(.A1(new_n1127), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1084), .A2(KEYINPUT63), .A3(new_n596), .A4(new_n1096), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT63), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1060), .A2(new_n1083), .A3(new_n596), .A4(new_n1064), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1132), .B1(new_n1133), .B2(new_n1088), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1130), .B1(new_n1131), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1100), .A2(KEYINPUT62), .ZN(new_n1136));
  AOI21_X1  g711(.A(G301), .B1(new_n1107), .B2(new_n1111), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT62), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1094), .A2(new_n1138), .A3(new_n1098), .A4(new_n1099), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1136), .A2(new_n1084), .A3(new_n1137), .A4(new_n1139), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1122), .A2(new_n1123), .A3(new_n1135), .A4(new_n1140), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1116), .A2(new_n994), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1142), .A2(new_n744), .A3(new_n924), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1142), .A2(G1986), .A3(G290), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  XOR2_X1   g720(.A(new_n1145), .B(KEYINPUT113), .Z(new_n1146));
  XNOR2_X1  g721(.A(new_n716), .B(new_n719), .ZN(new_n1147));
  OR2_X1    g722(.A1(new_n771), .A2(G1996), .ZN(new_n1148));
  XNOR2_X1  g723(.A(new_n806), .B(new_n1012), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n771), .A2(G1996), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1148), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1142), .B1(new_n1147), .B2(new_n1151), .ZN(new_n1152));
  AND2_X1   g727(.A1(new_n1146), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1141), .A2(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1143), .B(KEYINPUT48), .ZN(new_n1155));
  AND2_X1   g730(.A1(new_n1155), .A2(new_n1152), .ZN(new_n1156));
  NOR3_X1   g731(.A1(new_n1116), .A2(G1996), .A3(new_n994), .ZN(new_n1157));
  OR2_X1    g732(.A1(new_n1157), .A2(KEYINPUT46), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1149), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1142), .B1(new_n771), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1157), .A2(KEYINPUT46), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1158), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  XOR2_X1   g737(.A(new_n1162), .B(KEYINPUT47), .Z(new_n1163));
  OR2_X1    g738(.A1(new_n716), .A2(new_n719), .ZN(new_n1164));
  OAI22_X1  g739(.A1(new_n1164), .A2(new_n1151), .B1(G2067), .B2(new_n806), .ZN(new_n1165));
  AOI211_X1 g740(.A(new_n1156), .B(new_n1163), .C1(new_n1142), .C2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1154), .A2(new_n1166), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g742(.A(G319), .B1(new_n705), .B2(new_n706), .ZN(new_n1169));
  NOR2_X1   g743(.A1(G227), .A2(G401), .ZN(new_n1170));
  NAND2_X1  g744(.A1(new_n886), .A2(new_n1170), .ZN(new_n1171));
  NOR3_X1   g745(.A1(new_n976), .A2(new_n1169), .A3(new_n1171), .ZN(G308));
  INV_X1    g746(.A(new_n1169), .ZN(new_n1173));
  AND2_X1   g747(.A1(new_n886), .A2(new_n1170), .ZN(new_n1174));
  AND2_X1   g748(.A1(new_n975), .A2(new_n970), .ZN(new_n1175));
  OAI211_X1 g749(.A(new_n1173), .B(new_n1174), .C1(new_n1175), .C2(new_n974), .ZN(G225));
endmodule


