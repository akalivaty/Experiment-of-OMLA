//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 0 1 1 1 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 1 1 0 1 0 0 1 0 0 1 0 1 1 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:01 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(G107), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n189), .A2(KEYINPUT75), .A3(G104), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT3), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n189), .A2(G104), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT3), .ZN(new_n194));
  NAND4_X1  g008(.A1(new_n194), .A2(new_n189), .A3(KEYINPUT75), .A4(G104), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n191), .A2(new_n193), .A3(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT4), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(new_n197), .A3(G101), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(KEYINPUT76), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT76), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n196), .A2(new_n200), .A3(new_n197), .A4(G101), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G146), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G143), .ZN(new_n204));
  INV_X1    g018(.A(G143), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G146), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT0), .ZN(new_n208));
  INV_X1    g022(.A(G128), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NOR2_X1   g024(.A1(KEYINPUT0), .A2(G128), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n207), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  OAI211_X1 g026(.A(new_n204), .B(new_n206), .C1(new_n208), .C2(new_n209), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n196), .A2(G101), .ZN(new_n215));
  INV_X1    g029(.A(G101), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n191), .A2(new_n193), .A3(new_n216), .A4(new_n195), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n215), .A2(KEYINPUT4), .A3(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n202), .A2(new_n214), .A3(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G104), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n220), .A2(G107), .ZN(new_n221));
  OAI21_X1  g035(.A(G101), .B1(new_n192), .B2(new_n221), .ZN(new_n222));
  AND2_X1   g036(.A1(new_n217), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT77), .ZN(new_n224));
  OAI211_X1 g038(.A(new_n224), .B(KEYINPUT1), .C1(new_n205), .C2(G146), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G128), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n224), .B1(new_n204), .B2(KEYINPUT1), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n207), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT1), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n204), .A2(new_n206), .A3(new_n229), .A4(G128), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n223), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT10), .ZN(new_n233));
  AND3_X1   g047(.A1(new_n204), .A2(new_n206), .A3(G128), .ZN(new_n234));
  OAI21_X1  g048(.A(KEYINPUT1), .B1(new_n205), .B2(G146), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G128), .ZN(new_n236));
  AOI22_X1  g050(.A1(new_n234), .A2(new_n229), .B1(new_n236), .B2(new_n207), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n237), .A2(new_n233), .ZN(new_n238));
  AOI22_X1  g052(.A1(new_n232), .A2(new_n233), .B1(new_n223), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT11), .ZN(new_n240));
  INV_X1    g054(.A(G134), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n240), .B1(new_n241), .B2(G137), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(G137), .ZN(new_n243));
  INV_X1    g057(.A(G137), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n244), .A2(KEYINPUT11), .A3(G134), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n242), .A2(new_n243), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G131), .ZN(new_n247));
  INV_X1    g061(.A(G131), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n242), .A2(new_n245), .A3(new_n248), .A4(new_n243), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n219), .A2(new_n239), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(KEYINPUT78), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT78), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n219), .A2(new_n239), .A3(new_n254), .A4(new_n251), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g070(.A(G110), .B(G140), .ZN(new_n257));
  XNOR2_X1  g071(.A(new_n257), .B(KEYINPUT74), .ZN(new_n258));
  INV_X1    g072(.A(G953), .ZN(new_n259));
  AND2_X1   g073(.A1(new_n259), .A2(G227), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n258), .B(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n217), .A2(new_n222), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n263), .B1(new_n230), .B2(new_n228), .ZN(new_n264));
  AND2_X1   g078(.A1(new_n263), .A2(new_n237), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n250), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  XOR2_X1   g080(.A(new_n266), .B(KEYINPUT12), .Z(new_n267));
  AND3_X1   g081(.A1(new_n256), .A2(new_n262), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n219), .A2(new_n239), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n250), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n262), .B1(new_n256), .B2(new_n270), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n187), .B(new_n188), .C1(new_n268), .C2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(G469), .A2(G902), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n261), .B1(new_n253), .B2(new_n255), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(new_n270), .ZN(new_n275));
  AND2_X1   g089(.A1(new_n256), .A2(new_n267), .ZN(new_n276));
  OAI211_X1 g090(.A(G469), .B(new_n275), .C1(new_n276), .C2(new_n262), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n272), .A2(new_n273), .A3(new_n277), .ZN(new_n278));
  XOR2_X1   g092(.A(KEYINPUT9), .B(G234), .Z(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(G221), .B1(new_n280), .B2(G902), .ZN(new_n281));
  AND2_X1   g095(.A1(new_n278), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G475), .ZN(new_n283));
  NAND2_X1  g097(.A1(G125), .A2(G140), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  NOR2_X1   g099(.A1(G125), .A2(G140), .ZN(new_n286));
  OAI21_X1  g100(.A(KEYINPUT16), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(G125), .ZN(new_n288));
  NOR3_X1   g102(.A1(new_n288), .A2(KEYINPUT16), .A3(G140), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n287), .A2(new_n290), .A3(G146), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT19), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n292), .B1(new_n285), .B2(new_n286), .ZN(new_n293));
  INV_X1    g107(.A(G140), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n288), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n295), .A2(KEYINPUT19), .A3(new_n284), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n293), .A2(new_n296), .A3(new_n203), .ZN(new_n297));
  NOR2_X1   g111(.A1(G237), .A2(G953), .ZN(new_n298));
  AND3_X1   g112(.A1(new_n298), .A2(G143), .A3(G214), .ZN(new_n299));
  AOI21_X1  g113(.A(G143), .B1(new_n298), .B2(G214), .ZN(new_n300));
  NOR3_X1   g114(.A1(new_n299), .A2(new_n300), .A3(G131), .ZN(new_n301));
  INV_X1    g115(.A(G237), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n302), .A2(new_n259), .A3(G214), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n205), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n298), .A2(G143), .A3(G214), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n248), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n291), .B(new_n297), .C1(new_n301), .C2(new_n306), .ZN(new_n307));
  OAI211_X1 g121(.A(KEYINPUT18), .B(G131), .C1(new_n299), .C2(new_n300), .ZN(new_n308));
  NAND2_X1  g122(.A1(KEYINPUT18), .A2(G131), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n304), .A2(new_n305), .A3(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n203), .B1(new_n285), .B2(new_n286), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n295), .A2(G146), .A3(new_n284), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n308), .A2(new_n310), .A3(new_n313), .ZN(new_n314));
  AND3_X1   g128(.A1(new_n307), .A2(KEYINPUT88), .A3(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(KEYINPUT88), .B1(new_n307), .B2(new_n314), .ZN(new_n316));
  XNOR2_X1  g130(.A(G113), .B(G122), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n317), .B(new_n220), .ZN(new_n318));
  NOR3_X1   g132(.A1(new_n315), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n318), .ZN(new_n320));
  INV_X1    g134(.A(new_n314), .ZN(new_n321));
  OAI21_X1  g135(.A(G131), .B1(new_n299), .B2(new_n300), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT17), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n304), .A2(new_n248), .A3(new_n305), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n306), .A2(KEYINPUT17), .ZN(new_n326));
  AND2_X1   g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT16), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n328), .B1(new_n295), .B2(new_n284), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n203), .B1(new_n329), .B2(new_n289), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n330), .A2(KEYINPUT69), .A3(new_n291), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT69), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n332), .B(new_n203), .C1(new_n329), .C2(new_n289), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  AOI211_X1 g148(.A(new_n320), .B(new_n321), .C1(new_n327), .C2(new_n334), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n283), .B(new_n188), .C1(new_n319), .C2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT20), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n321), .B1(new_n327), .B2(new_n334), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n339), .A2(new_n318), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n188), .B1(new_n340), .B2(new_n335), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G475), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n339), .A2(new_n318), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n307), .A2(new_n314), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT88), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n307), .A2(KEYINPUT88), .A3(new_n314), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n346), .A2(new_n320), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n343), .A2(new_n348), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n349), .A2(KEYINPUT20), .A3(new_n283), .A4(new_n188), .ZN(new_n350));
  AND3_X1   g164(.A1(new_n338), .A2(new_n342), .A3(new_n350), .ZN(new_n351));
  XNOR2_X1  g165(.A(KEYINPUT21), .B(G898), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n352), .B(KEYINPUT91), .ZN(new_n353));
  NAND2_X1  g167(.A1(G234), .A2(G237), .ZN(new_n354));
  AND3_X1   g168(.A1(new_n354), .A2(G902), .A3(G953), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  AND3_X1   g170(.A1(new_n354), .A2(G952), .A3(new_n259), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n279), .A2(G217), .A3(new_n259), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(G116), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(G122), .ZN(new_n363));
  INV_X1    g177(.A(G122), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G116), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT14), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n363), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n362), .A2(KEYINPUT14), .A3(G122), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n367), .A2(G107), .A3(new_n368), .ZN(new_n369));
  XNOR2_X1  g183(.A(G116), .B(G122), .ZN(new_n370));
  AOI21_X1  g184(.A(KEYINPUT89), .B1(new_n370), .B2(new_n189), .ZN(new_n371));
  AND4_X1   g185(.A1(KEYINPUT89), .A2(new_n363), .A3(new_n365), .A4(new_n189), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n369), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n205), .A2(G128), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n209), .A2(G143), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G134), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n374), .A2(new_n375), .A3(new_n241), .ZN(new_n378));
  AND2_X1   g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g193(.A(KEYINPUT90), .B1(new_n373), .B2(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n363), .A2(new_n365), .A3(new_n189), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT89), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n370), .A2(KEYINPUT89), .A3(new_n189), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n377), .A2(new_n378), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT90), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n385), .A2(new_n386), .A3(new_n387), .A4(new_n369), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n380), .A2(new_n388), .ZN(new_n389));
  AND3_X1   g203(.A1(new_n374), .A2(new_n375), .A3(KEYINPUT13), .ZN(new_n390));
  OAI21_X1  g204(.A(G134), .B1(new_n374), .B2(KEYINPUT13), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n378), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n381), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n189), .B1(new_n363), .B2(new_n365), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n361), .B1(new_n389), .B2(new_n397), .ZN(new_n398));
  AOI211_X1 g212(.A(new_n396), .B(new_n360), .C1(new_n380), .C2(new_n388), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n188), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT15), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(G478), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n400), .B(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n351), .A2(new_n359), .A3(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT92), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n351), .A2(KEYINPUT92), .A3(new_n359), .A4(new_n403), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(G214), .B1(G237), .B2(G902), .ZN(new_n409));
  NOR2_X1   g223(.A1(KEYINPUT2), .A2(G113), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(KEYINPUT65), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT65), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n412), .B1(KEYINPUT2), .B2(G113), .ZN(new_n413));
  AOI22_X1  g227(.A1(new_n411), .A2(new_n413), .B1(KEYINPUT2), .B2(G113), .ZN(new_n414));
  INV_X1    g228(.A(G119), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(G116), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n362), .A2(G119), .ZN(new_n417));
  AND2_X1   g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n414), .B(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n202), .A2(new_n419), .A3(new_n218), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n416), .A2(new_n417), .A3(KEYINPUT5), .ZN(new_n421));
  OR3_X1    g235(.A1(new_n362), .A2(KEYINPUT5), .A3(G119), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n421), .A2(new_n422), .A3(G113), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(KEYINPUT79), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n414), .A2(new_n418), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT79), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n421), .A2(new_n422), .A3(new_n426), .A4(G113), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n424), .A2(new_n425), .A3(new_n427), .ZN(new_n428));
  OR2_X1    g242(.A1(new_n428), .A2(new_n263), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n420), .A2(new_n429), .ZN(new_n430));
  XOR2_X1   g244(.A(G110), .B(G122), .Z(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n431), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n420), .A2(new_n429), .A3(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n432), .A2(KEYINPUT6), .A3(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT6), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n430), .A2(new_n436), .A3(new_n431), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n236), .A2(new_n207), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(new_n288), .A3(new_n230), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(KEYINPUT80), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT80), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n438), .A2(new_n441), .A3(new_n288), .A4(new_n230), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n212), .A2(G125), .A3(new_n213), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n259), .A2(G224), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n446), .B(KEYINPUT81), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n445), .B(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n435), .A2(new_n437), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(KEYINPUT82), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT82), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n435), .A2(new_n452), .A3(new_n437), .A4(new_n449), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT83), .ZN(new_n455));
  AND3_X1   g269(.A1(new_n428), .A2(new_n455), .A3(new_n263), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n455), .B1(new_n428), .B2(new_n263), .ZN(new_n457));
  AND3_X1   g271(.A1(new_n223), .A2(new_n425), .A3(new_n423), .ZN(new_n458));
  NOR3_X1   g272(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n431), .B(KEYINPUT8), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n434), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT7), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT85), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n462), .B1(new_n447), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n448), .A2(KEYINPUT85), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n443), .A2(new_n444), .A3(new_n464), .A4(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT84), .ZN(new_n467));
  AND3_X1   g281(.A1(new_n440), .A2(new_n467), .A3(new_n442), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n467), .B1(new_n440), .B2(new_n442), .ZN(new_n469));
  INV_X1    g283(.A(new_n444), .ZN(new_n470));
  NOR3_X1   g284(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n448), .A2(new_n462), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n466), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n188), .B1(new_n461), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT86), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OAI211_X1 g290(.A(KEYINPUT86), .B(new_n188), .C1(new_n461), .C2(new_n473), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(G210), .B1(G237), .B2(G902), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n454), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  AOI22_X1  g294(.A1(new_n453), .A2(new_n451), .B1(new_n476), .B2(new_n477), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n479), .B(KEYINPUT87), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n282), .A2(new_n408), .A3(new_n409), .A4(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n415), .A2(G128), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT23), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n487), .B1(G119), .B2(new_n209), .ZN(new_n488));
  NOR3_X1   g302(.A1(new_n415), .A2(KEYINPUT23), .A3(G128), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n486), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT68), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n491), .B1(new_n209), .B2(G119), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n415), .A2(KEYINPUT68), .A3(G128), .ZN(new_n493));
  AOI22_X1  g307(.A1(new_n492), .A2(new_n493), .B1(G119), .B2(new_n209), .ZN(new_n494));
  XOR2_X1   g308(.A(KEYINPUT24), .B(G110), .Z(new_n495));
  AOI22_X1  g309(.A1(new_n490), .A2(G110), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n331), .A2(new_n496), .A3(new_n333), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(KEYINPUT70), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT70), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n331), .A2(new_n496), .A3(new_n499), .A4(new_n333), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(G110), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n502), .B(new_n486), .C1(new_n488), .C2(new_n489), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT71), .ZN(new_n504));
  OR2_X1    g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n503), .A2(new_n504), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n505), .B(new_n506), .C1(new_n494), .C2(new_n495), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n507), .A2(new_n291), .A3(new_n311), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n501), .A2(KEYINPUT72), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(KEYINPUT72), .B1(new_n501), .B2(new_n508), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n259), .A2(G221), .A3(G234), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n511), .B(KEYINPUT22), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(G137), .ZN(new_n513));
  NOR3_X1   g327(.A1(new_n509), .A2(new_n510), .A3(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n513), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n515), .B1(new_n501), .B2(new_n508), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n188), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(KEYINPUT25), .ZN(new_n518));
  INV_X1    g332(.A(G217), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n519), .B1(G234), .B2(new_n188), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT25), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n521), .B(new_n188), .C1(new_n514), .C2(new_n516), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n518), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(KEYINPUT73), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT73), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n518), .A2(new_n525), .A3(new_n520), .A4(new_n522), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n520), .A2(G902), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n527), .B1(new_n514), .B2(new_n516), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n524), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT30), .ZN(new_n530));
  OR2_X1    g344(.A1(new_n530), .A2(KEYINPUT64), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(KEYINPUT64), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n244), .A2(G134), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n241), .A2(G137), .ZN(new_n534));
  OAI21_X1  g348(.A(G131), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n249), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n237), .A2(new_n536), .ZN(new_n537));
  AOI22_X1  g351(.A1(new_n247), .A2(new_n249), .B1(new_n212), .B2(new_n213), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n531), .B(new_n532), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n250), .A2(new_n214), .ZN(new_n540));
  INV_X1    g354(.A(new_n230), .ZN(new_n541));
  AOI22_X1  g355(.A1(new_n235), .A2(G128), .B1(new_n204), .B2(new_n206), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n249), .B(new_n535), .C1(new_n541), .C2(new_n542), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n540), .A2(KEYINPUT64), .A3(new_n530), .A4(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n539), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n419), .ZN(new_n546));
  XOR2_X1   g360(.A(new_n414), .B(new_n418), .Z(new_n547));
  NAND3_X1  g361(.A1(new_n547), .A2(new_n540), .A3(new_n543), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g363(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n550), .B(G101), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n298), .A2(G210), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n551), .B(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n549), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT29), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n547), .B1(new_n540), .B2(new_n543), .ZN(new_n557));
  NOR3_X1   g371(.A1(new_n419), .A2(new_n537), .A3(new_n538), .ZN(new_n558));
  OAI21_X1  g372(.A(KEYINPUT28), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(KEYINPUT67), .B1(new_n558), .B2(KEYINPUT28), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT67), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT28), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n548), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n559), .A2(new_n560), .A3(new_n553), .A4(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n555), .A2(new_n556), .A3(new_n564), .ZN(new_n565));
  AND2_X1   g379(.A1(new_n560), .A2(new_n563), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n566), .A2(KEYINPUT29), .A3(new_n553), .A4(new_n559), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n565), .A2(new_n567), .A3(new_n188), .ZN(new_n568));
  AND2_X1   g382(.A1(new_n568), .A2(G472), .ZN(new_n569));
  INV_X1    g383(.A(G472), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT31), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n546), .A2(new_n548), .A3(new_n553), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT66), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n558), .B1(new_n545), .B2(new_n419), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n575), .A2(KEYINPUT66), .A3(new_n553), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n571), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n559), .A2(new_n560), .A3(new_n563), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n554), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n575), .A2(new_n571), .A3(new_n553), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n570), .B(new_n188), .C1(new_n577), .C2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(KEYINPUT32), .ZN(new_n583));
  INV_X1    g397(.A(new_n572), .ZN(new_n584));
  AOI22_X1  g398(.A1(new_n584), .A2(new_n571), .B1(new_n578), .B2(new_n554), .ZN(new_n585));
  AOI21_X1  g399(.A(KEYINPUT66), .B1(new_n575), .B2(new_n553), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n547), .B1(new_n539), .B2(new_n544), .ZN(new_n587));
  NOR4_X1   g401(.A1(new_n587), .A2(new_n573), .A3(new_n558), .A4(new_n554), .ZN(new_n588));
  OAI21_X1  g402(.A(KEYINPUT31), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT32), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n590), .A2(new_n591), .A3(new_n570), .A4(new_n188), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n569), .B1(new_n583), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n529), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n485), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(G101), .ZN(G3));
  AND3_X1   g410(.A1(new_n524), .A2(new_n526), .A3(new_n528), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n188), .B1(new_n577), .B2(new_n581), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(G472), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n582), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n597), .A2(new_n282), .A3(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n409), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n454), .A2(new_n478), .ZN(new_n604));
  INV_X1    g418(.A(new_n479), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n603), .B1(new_n606), .B2(new_n480), .ZN(new_n607));
  INV_X1    g421(.A(G478), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n189), .B1(new_n370), .B2(new_n366), .ZN(new_n609));
  AOI22_X1  g423(.A1(new_n368), .A2(new_n609), .B1(new_n383), .B2(new_n384), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n387), .B1(new_n610), .B2(new_n386), .ZN(new_n611));
  INV_X1    g425(.A(new_n388), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n397), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n360), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n389), .A2(new_n397), .A3(new_n361), .ZN(new_n615));
  XOR2_X1   g429(.A(KEYINPUT93), .B(KEYINPUT33), .Z(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n614), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(KEYINPUT93), .A2(KEYINPUT33), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n619), .B1(new_n398), .B2(new_n399), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n608), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  OAI211_X1 g435(.A(new_n608), .B(new_n188), .C1(new_n398), .C2(new_n399), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n608), .A2(new_n188), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n621), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n338), .A2(new_n342), .A3(new_n350), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n607), .A2(new_n359), .A3(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n602), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT34), .B(G104), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(KEYINPUT94), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n630), .B(new_n632), .ZN(G6));
  INV_X1    g447(.A(new_n403), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n351), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  XOR2_X1   g450(.A(new_n359), .B(KEYINPUT95), .Z(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n607), .A2(new_n636), .A3(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n602), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(KEYINPUT35), .B(G107), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G9));
  NOR2_X1   g456(.A1(new_n509), .A2(new_n510), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n515), .A2(KEYINPUT36), .ZN(new_n644));
  XOR2_X1   g458(.A(new_n643), .B(new_n644), .Z(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n527), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n524), .A2(new_n526), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n601), .ZN(new_n648));
  OR2_X1    g462(.A1(new_n484), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(KEYINPUT37), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(new_n502), .ZN(G12));
  NAND2_X1  g465(.A1(new_n278), .A2(new_n281), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n593), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT96), .B(G900), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n357), .B1(new_n355), .B2(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n635), .A2(new_n655), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n653), .A2(new_n607), .A3(new_n647), .A4(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G128), .ZN(G30));
  XNOR2_X1  g472(.A(new_n483), .B(KEYINPUT38), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n554), .B1(new_n557), .B2(new_n558), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n570), .B1(new_n660), .B2(KEYINPUT97), .ZN(new_n661));
  OAI221_X1 g475(.A(new_n661), .B1(KEYINPUT97), .B2(new_n660), .C1(new_n586), .C2(new_n588), .ZN(new_n662));
  NAND2_X1  g476(.A1(G472), .A2(G902), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(KEYINPUT98), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT98), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n662), .A2(new_n666), .A3(new_n663), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n668), .B1(new_n583), .B2(new_n592), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n669), .A2(new_n647), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n351), .A2(new_n403), .ZN(new_n671));
  AND4_X1   g485(.A1(new_n409), .A2(new_n659), .A3(new_n670), .A4(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(new_n655), .B(KEYINPUT39), .Z(new_n673));
  NAND2_X1  g487(.A1(new_n282), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(KEYINPUT99), .ZN(new_n675));
  AND2_X1   g489(.A1(new_n675), .A2(KEYINPUT40), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n675), .A2(KEYINPUT40), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n672), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G143), .ZN(G45));
  NAND2_X1  g493(.A1(new_n618), .A2(new_n620), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n624), .B1(new_n680), .B2(G478), .ZN(new_n681));
  INV_X1    g495(.A(new_n655), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n626), .A2(new_n681), .A3(new_n622), .A4(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT100), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n625), .A2(KEYINPUT100), .A3(new_n626), .A4(new_n682), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n653), .A2(new_n607), .A3(new_n647), .A4(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G146), .ZN(G48));
  INV_X1    g504(.A(new_n569), .ZN(new_n691));
  INV_X1    g505(.A(new_n592), .ZN(new_n692));
  AOI21_X1  g506(.A(G902), .B1(new_n585), .B2(new_n589), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n591), .B1(new_n693), .B2(new_n570), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n691), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n281), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n256), .A2(new_n270), .ZN(new_n697));
  AOI22_X1  g511(.A1(new_n697), .A2(new_n261), .B1(new_n274), .B2(new_n267), .ZN(new_n698));
  OAI21_X1  g512(.A(G469), .B1(new_n698), .B2(G902), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n699), .A2(KEYINPUT101), .A3(new_n272), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT101), .ZN(new_n701));
  OAI211_X1 g515(.A(new_n701), .B(G469), .C1(new_n698), .C2(G902), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n696), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n597), .A2(new_n695), .A3(new_n703), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n704), .A2(new_n629), .ZN(new_n705));
  XOR2_X1   g519(.A(KEYINPUT41), .B(G113), .Z(new_n706));
  XOR2_X1   g520(.A(new_n706), .B(KEYINPUT102), .Z(new_n707));
  XNOR2_X1  g521(.A(new_n705), .B(new_n707), .ZN(G15));
  NOR2_X1   g522(.A1(new_n704), .A2(new_n639), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(new_n362), .ZN(G18));
  NAND4_X1  g524(.A1(new_n703), .A2(new_n647), .A3(new_n607), .A4(new_n695), .ZN(new_n711));
  INV_X1    g525(.A(new_n408), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(new_n415), .ZN(G21));
  NAND3_X1  g528(.A1(new_n599), .A2(KEYINPUT103), .A3(new_n582), .ZN(new_n715));
  OR3_X1    g529(.A1(new_n693), .A2(KEYINPUT103), .A3(new_n570), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n597), .A2(new_n703), .A3(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n607), .A2(new_n638), .A3(new_n671), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(new_n364), .ZN(G24));
  AOI21_X1  g535(.A(new_n687), .B1(new_n716), .B2(new_n715), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n722), .A2(new_n607), .A3(new_n647), .A4(new_n703), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G125), .ZN(G27));
  OAI211_X1 g538(.A(new_n480), .B(new_n409), .C1(new_n482), .C2(new_n481), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n725), .A2(new_n652), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n594), .A2(new_n688), .A3(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT42), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n594), .A2(KEYINPUT42), .A3(new_n688), .A4(new_n726), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G131), .ZN(G33));
  NAND4_X1  g546(.A1(new_n726), .A2(new_n597), .A3(new_n695), .A4(new_n656), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(KEYINPUT104), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT104), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n594), .A2(new_n735), .A3(new_n656), .A4(new_n726), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G134), .ZN(G36));
  OAI21_X1  g552(.A(new_n275), .B1(new_n276), .B2(new_n262), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT45), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  OAI211_X1 g555(.A(KEYINPUT45), .B(new_n275), .C1(new_n276), .C2(new_n262), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n741), .A2(G469), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n273), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT46), .ZN(new_n745));
  OAI21_X1  g559(.A(KEYINPUT105), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n744), .A2(new_n745), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT105), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n743), .A2(new_n748), .A3(KEYINPUT46), .A4(new_n273), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n746), .A2(new_n747), .A3(new_n272), .A4(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n750), .A2(new_n281), .A3(new_n673), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(KEYINPUT106), .ZN(new_n752));
  INV_X1    g566(.A(new_n625), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n753), .A2(new_n626), .ZN(new_n754));
  XOR2_X1   g568(.A(new_n754), .B(KEYINPUT43), .Z(new_n755));
  NOR2_X1   g569(.A1(new_n755), .A2(new_n601), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n647), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT44), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(new_n725), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n756), .A2(KEYINPUT44), .A3(new_n647), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n759), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n752), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G137), .ZN(G39));
  NOR3_X1   g579(.A1(new_n597), .A2(new_n695), .A3(new_n725), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n750), .A2(KEYINPUT47), .A3(new_n281), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(KEYINPUT47), .B1(new_n750), .B2(new_n281), .ZN(new_n769));
  OAI211_X1 g583(.A(new_n688), .B(new_n766), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G140), .ZN(G42));
  NAND2_X1  g585(.A1(new_n272), .A2(KEYINPUT101), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n274), .A2(new_n267), .ZN(new_n773));
  AOI22_X1  g587(.A1(new_n253), .A2(new_n255), .B1(new_n250), .B2(new_n269), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n773), .B1(new_n774), .B2(new_n262), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n187), .B1(new_n775), .B2(new_n188), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n772), .A2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(new_n702), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(KEYINPUT49), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n669), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT107), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n597), .A2(new_n281), .A3(new_n409), .A4(new_n754), .ZN(new_n783));
  AOI211_X1 g597(.A(new_n659), .B(new_n781), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  OAI221_X1 g598(.A(new_n784), .B1(new_n782), .B2(new_n783), .C1(KEYINPUT49), .C2(new_n779), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n755), .A2(new_n358), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n760), .A2(new_n703), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(new_n594), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(KEYINPUT48), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n259), .A2(G952), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n669), .A2(new_n357), .ZN(new_n792));
  NOR3_X1   g606(.A1(new_n792), .A2(new_n787), .A3(new_n529), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n791), .B1(new_n793), .B2(new_n628), .ZN(new_n794));
  INV_X1    g608(.A(new_n718), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n755), .A2(new_n358), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n795), .A2(new_n607), .A3(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n790), .A2(new_n794), .A3(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(KEYINPUT114), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT51), .ZN(new_n800));
  INV_X1    g614(.A(new_n717), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n786), .A2(new_n529), .A3(new_n801), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n281), .B1(new_n777), .B2(new_n778), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n659), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n802), .A2(new_n603), .A3(new_n804), .ZN(new_n805));
  XOR2_X1   g619(.A(new_n805), .B(KEYINPUT50), .Z(new_n806));
  AND2_X1   g620(.A1(new_n802), .A2(new_n760), .ZN(new_n807));
  INV_X1    g621(.A(new_n769), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n808), .A2(KEYINPUT111), .A3(new_n767), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n696), .B1(new_n777), .B2(new_n778), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n768), .A2(new_n769), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n812), .A2(KEYINPUT111), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n807), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n806), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n788), .A2(new_n647), .A3(new_n717), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n793), .A2(new_n351), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n817), .A2(KEYINPUT112), .A3(new_n753), .ZN(new_n818));
  AOI21_X1  g632(.A(KEYINPUT112), .B1(new_n817), .B2(new_n753), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n816), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n800), .B1(new_n815), .B2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT113), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n812), .A2(new_n810), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n800), .B1(new_n824), .B2(new_n807), .ZN(new_n825));
  OAI211_X1 g639(.A(KEYINPUT113), .B(new_n816), .C1(new_n818), .C2(new_n819), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n823), .A2(new_n806), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n821), .A2(new_n827), .ZN(new_n828));
  NOR4_X1   g642(.A1(new_n593), .A2(new_n634), .A3(new_n626), .A4(new_n655), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n647), .B(new_n726), .C1(new_n829), .C2(new_n722), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n731), .A2(new_n737), .A3(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n719), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n803), .A2(new_n529), .A3(new_n593), .ZN(new_n833));
  INV_X1    g647(.A(new_n629), .ZN(new_n834));
  AOI22_X1  g648(.A1(new_n795), .A2(new_n832), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(new_n711), .ZN(new_n836));
  INV_X1    g650(.A(new_n639), .ZN(new_n837));
  AOI22_X1  g651(.A1(new_n836), .A2(new_n408), .B1(new_n833), .B2(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n695), .A2(new_n526), .A3(new_n524), .A4(new_n528), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n484), .B1(new_n839), .B2(new_n648), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n635), .A2(new_n627), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n483), .A2(new_n409), .A3(new_n638), .A4(new_n841), .ZN(new_n842));
  NOR4_X1   g656(.A1(new_n842), .A2(new_n529), .A3(new_n652), .A4(new_n600), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n835), .A2(new_n838), .A3(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n831), .A2(new_n845), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n689), .A2(new_n723), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n606), .A2(new_n480), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n848), .A2(new_n409), .A3(new_n671), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n670), .A2(new_n850), .A3(new_n282), .A4(new_n682), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n847), .A2(KEYINPUT108), .A3(new_n657), .A4(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT108), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n657), .A2(new_n689), .A3(new_n723), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n848), .A2(new_n409), .A3(new_n682), .A4(new_n671), .ZN(new_n855));
  NOR4_X1   g669(.A1(new_n855), .A2(new_n669), .A3(new_n647), .A4(new_n652), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n853), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT52), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n852), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n858), .B1(new_n852), .B2(new_n857), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n846), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(KEYINPUT53), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n852), .A2(new_n857), .A3(new_n858), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n657), .A2(new_n689), .A3(new_n723), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n864), .A2(KEYINPUT52), .A3(new_n851), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT53), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n866), .A2(new_n867), .A3(new_n846), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n862), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n869), .A2(KEYINPUT109), .A3(KEYINPUT54), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n862), .A2(KEYINPUT54), .A3(new_n868), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT109), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n831), .A2(new_n867), .ZN(new_n873));
  INV_X1    g687(.A(new_n844), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n835), .A2(new_n838), .A3(KEYINPUT110), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT110), .ZN(new_n876));
  OAI22_X1  g690(.A1(new_n629), .A2(new_n704), .B1(new_n718), .B2(new_n719), .ZN(new_n877));
  OAI22_X1  g691(.A1(new_n704), .A2(new_n639), .B1(new_n711), .B2(new_n712), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n874), .B1(new_n875), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n866), .A2(new_n873), .A3(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT54), .ZN(new_n882));
  AOI22_X1  g696(.A1(new_n729), .A2(new_n730), .B1(new_n734), .B2(new_n736), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n877), .A2(new_n878), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n883), .A2(new_n884), .A3(new_n844), .A4(new_n830), .ZN(new_n885));
  AOI21_X1  g699(.A(KEYINPUT108), .B1(new_n864), .B2(new_n851), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n854), .A2(new_n856), .A3(new_n853), .ZN(new_n887));
  OAI21_X1  g701(.A(KEYINPUT52), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n885), .B1(new_n888), .B2(new_n863), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n881), .B(new_n882), .C1(new_n889), .C2(KEYINPUT53), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n871), .A2(new_n872), .A3(new_n890), .ZN(new_n891));
  AOI211_X1 g705(.A(new_n799), .B(new_n828), .C1(new_n870), .C2(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(G952), .A2(G953), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT115), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n785), .B1(new_n892), .B2(new_n894), .ZN(G75));
  NOR2_X1   g709(.A1(new_n259), .A2(G952), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n896), .B(KEYINPUT118), .Z(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n861), .A2(new_n867), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n188), .B1(new_n899), .B2(new_n881), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT56), .B1(new_n900), .B2(G210), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n435), .A2(new_n437), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT116), .ZN(new_n903));
  XNOR2_X1  g717(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n449), .B(new_n904), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n903), .B(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n898), .B1(new_n901), .B2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n482), .ZN(new_n908));
  AOI21_X1  g722(.A(KEYINPUT56), .B1(new_n900), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n907), .B1(new_n906), .B2(new_n909), .ZN(G51));
  INV_X1    g724(.A(KEYINPUT119), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n273), .B(KEYINPUT57), .Z(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n888), .A2(new_n863), .ZN(new_n914));
  AOI21_X1  g728(.A(KEYINPUT53), .B1(new_n914), .B2(new_n846), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n866), .A2(new_n873), .A3(new_n880), .ZN(new_n916));
  OAI21_X1  g730(.A(KEYINPUT54), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n913), .B1(new_n917), .B2(new_n890), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n911), .B1(new_n918), .B2(new_n698), .ZN(new_n919));
  INV_X1    g733(.A(new_n890), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n882), .B1(new_n899), .B2(new_n881), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n912), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n922), .A2(KEYINPUT119), .A3(new_n775), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n743), .B(KEYINPUT120), .Z(new_n924));
  NAND2_X1  g738(.A1(new_n900), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n919), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(new_n896), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n926), .A2(new_n927), .ZN(G54));
  NAND3_X1  g742(.A1(new_n900), .A2(KEYINPUT58), .A3(G475), .ZN(new_n929));
  INV_X1    g743(.A(new_n349), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n929), .A2(new_n930), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n931), .A2(new_n932), .A3(new_n896), .ZN(G60));
  XOR2_X1   g747(.A(new_n624), .B(KEYINPUT59), .Z(new_n934));
  NAND3_X1  g748(.A1(new_n870), .A2(new_n891), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n897), .B1(new_n935), .B2(new_n680), .ZN(new_n936));
  INV_X1    g750(.A(new_n680), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n937), .B(new_n934), .C1(new_n920), .C2(new_n921), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n936), .A2(new_n938), .ZN(G63));
  NAND2_X1  g753(.A1(new_n899), .A2(new_n881), .ZN(new_n940));
  XNOR2_X1  g754(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n519), .A2(new_n188), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n941), .B(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n514), .A2(new_n516), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n940), .A2(new_n645), .A3(new_n943), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n946), .A2(new_n898), .A3(new_n947), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(KEYINPUT61), .Z(G66));
  INV_X1    g763(.A(G224), .ZN(new_n950));
  OAI21_X1  g764(.A(G953), .B1(new_n353), .B2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(new_n845), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n951), .B1(new_n952), .B2(G953), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n903), .B1(G898), .B2(new_n259), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n953), .B(new_n954), .ZN(G69));
  AOI21_X1  g769(.A(new_n259), .B1(G227), .B2(G900), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n854), .B(KEYINPUT122), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n762), .B1(new_n839), .B2(new_n849), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n958), .B1(new_n752), .B2(new_n959), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n770), .A2(new_n883), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n960), .A2(new_n259), .A3(new_n961), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n293), .A2(new_n296), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n545), .B(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(G900), .A2(G953), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n962), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n678), .A2(new_n957), .ZN(new_n967));
  XNOR2_X1  g781(.A(KEYINPUT123), .B(KEYINPUT62), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n594), .A2(new_n841), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n970), .A2(new_n674), .A3(new_n725), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n971), .B1(new_n752), .B2(new_n763), .ZN(new_n972));
  NAND2_X1  g786(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n678), .A2(new_n957), .A3(new_n973), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n969), .A2(new_n972), .A3(new_n770), .A4(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n964), .B1(new_n975), .B2(new_n259), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n956), .B1(new_n966), .B2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n976), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n966), .B1(new_n978), .B2(KEYINPUT124), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT125), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT124), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n956), .B1(new_n976), .B2(new_n981), .ZN(new_n982));
  AND3_X1   g796(.A1(new_n979), .A2(new_n980), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n980), .B1(new_n979), .B2(new_n982), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n977), .B1(new_n983), .B2(new_n984), .ZN(G72));
  NOR2_X1   g799(.A1(new_n975), .A2(new_n845), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n663), .B(KEYINPUT63), .ZN(new_n987));
  OAI211_X1 g801(.A(new_n549), .B(new_n553), .C1(new_n986), .C2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(new_n555), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT126), .ZN(new_n990));
  AOI22_X1  g804(.A1(new_n989), .A2(new_n990), .B1(new_n574), .B2(new_n576), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n555), .A2(KEYINPUT126), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n987), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n896), .B1(new_n869), .B2(new_n993), .ZN(new_n994));
  AND3_X1   g808(.A1(new_n960), .A2(new_n952), .A3(new_n961), .ZN(new_n995));
  OAI211_X1 g809(.A(new_n575), .B(new_n554), .C1(new_n995), .C2(new_n987), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n988), .A2(new_n994), .A3(new_n996), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n997), .B(KEYINPUT127), .ZN(G57));
endmodule


