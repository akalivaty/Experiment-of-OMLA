//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 0 0 1 0 1 1 0 0 1 1 0 1 0 0 1 0 1 1 0 1 1 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 1 1 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:47 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n561, new_n562, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n613, new_n614, new_n616, new_n617, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT66), .Z(G173));
  XNOR2_X1  g021(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  AOI22_X1  g037(.A1(new_n462), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n464), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n462), .A2(new_n464), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n465), .A2(new_n470), .ZN(G160));
  AND2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G136), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n474), .A2(new_n464), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n464), .A2(G112), .ZN(new_n479));
  OAI21_X1  g054(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n476), .B(new_n478), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT68), .ZN(G162));
  AND2_X1   g057(.A1(G126), .A2(G2105), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n483), .B1(new_n472), .B2(new_n473), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT69), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OAI211_X1 g061(.A(KEYINPUT69), .B(new_n483), .C1(new_n472), .C2(new_n473), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT70), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n464), .A2(G114), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OR2_X1    g066(.A1(G102), .A2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n492), .A2(new_n494), .A3(KEYINPUT70), .A4(G2104), .ZN(new_n495));
  AOI22_X1  g070(.A1(new_n486), .A2(new_n487), .B1(new_n491), .B2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(G138), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n498), .B1(new_n472), .B2(new_n473), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT4), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  OAI211_X1 g076(.A(new_n498), .B(new_n501), .C1(new_n473), .C2(new_n472), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n496), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  XNOR2_X1  g081(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  OAI21_X1  g083(.A(KEYINPUT72), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n510), .A2(G543), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT72), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT71), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n514), .A2(KEYINPUT5), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n510), .A2(KEYINPUT71), .ZN(new_n516));
  OAI211_X1 g091(.A(new_n513), .B(G543), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  AND3_X1   g092(.A1(new_n509), .A2(new_n512), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G62), .ZN(new_n519));
  NAND2_X1  g094(.A1(G75), .A2(G543), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n506), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AND2_X1   g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  NOR2_X1   g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n509), .A2(new_n512), .A3(new_n517), .A4(new_n524), .ZN(new_n525));
  XOR2_X1   g100(.A(KEYINPUT73), .B(G88), .Z(new_n526));
  INV_X1    g101(.A(G50), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n524), .A2(G543), .ZN(new_n528));
  OAI22_X1  g103(.A1(new_n525), .A2(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n521), .A2(new_n529), .ZN(G166));
  NAND3_X1  g105(.A1(new_n518), .A2(G63), .A3(G651), .ZN(new_n531));
  AND4_X1   g106(.A1(new_n509), .A2(new_n512), .A3(new_n517), .A4(new_n524), .ZN(new_n532));
  XNOR2_X1  g107(.A(KEYINPUT74), .B(G89), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(new_n528), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(KEYINPUT7), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n536), .A2(KEYINPUT7), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n535), .A2(G51), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AND3_X1   g114(.A1(new_n531), .A2(new_n534), .A3(new_n539), .ZN(G168));
  NAND2_X1  g115(.A1(new_n518), .A2(G64), .ZN(new_n541));
  NAND2_X1  g116(.A1(G77), .A2(G543), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n506), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(G90), .ZN(new_n544));
  INV_X1    g119(.A(G52), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n525), .A2(new_n544), .B1(new_n545), .B2(new_n528), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n543), .A2(new_n546), .ZN(G171));
  NAND2_X1  g122(.A1(new_n510), .A2(KEYINPUT71), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n514), .A2(KEYINPUT5), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n508), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n511), .B1(new_n550), .B2(new_n513), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n551), .A2(G56), .A3(new_n509), .ZN(new_n552));
  NAND2_X1  g127(.A1(G68), .A2(G543), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n506), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(G81), .ZN(new_n555));
  INV_X1    g130(.A(G43), .ZN(new_n556));
  OAI22_X1  g131(.A1(new_n525), .A2(new_n555), .B1(new_n556), .B2(new_n528), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  NAND4_X1  g134(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND4_X1  g137(.A1(G319), .A2(G483), .A3(G661), .A4(new_n562), .ZN(G188));
  OAI211_X1 g138(.A(G53), .B(G543), .C1(new_n522), .C2(new_n523), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT9), .ZN(new_n565));
  INV_X1    g140(.A(G91), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n525), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n509), .A2(new_n512), .A3(new_n517), .ZN(new_n569));
  INV_X1    g144(.A(G65), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n567), .B1(G651), .B2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(G299));
  INV_X1    g148(.A(G171), .ZN(G301));
  INV_X1    g149(.A(G168), .ZN(G286));
  INV_X1    g150(.A(G166), .ZN(G303));
  NAND4_X1  g151(.A1(new_n551), .A2(G87), .A3(new_n509), .A4(new_n524), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n535), .A2(G49), .ZN(new_n578));
  AOI21_X1  g153(.A(G74), .B1(new_n551), .B2(new_n509), .ZN(new_n579));
  OAI211_X1 g154(.A(new_n577), .B(new_n578), .C1(new_n579), .C2(new_n506), .ZN(G288));
  INV_X1    g155(.A(G86), .ZN(new_n581));
  INV_X1    g156(.A(G48), .ZN(new_n582));
  OAI22_X1  g157(.A1(new_n525), .A2(new_n581), .B1(new_n582), .B2(new_n528), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n509), .A2(G61), .A3(new_n517), .A4(new_n512), .ZN(new_n584));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n506), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G305));
  NAND2_X1  g163(.A1(G72), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G60), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n569), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n591), .A2(G651), .ZN(new_n592));
  XOR2_X1   g167(.A(KEYINPUT75), .B(G47), .Z(new_n593));
  AOI22_X1  g168(.A1(new_n532), .A2(G85), .B1(new_n535), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n592), .A2(new_n594), .ZN(G290));
  NAND2_X1  g170(.A1(G79), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G66), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n569), .B2(new_n597), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n598), .A2(G651), .B1(G54), .B2(new_n535), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n532), .A2(KEYINPUT10), .A3(G92), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT10), .ZN(new_n601));
  INV_X1    g176(.A(G92), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n525), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n599), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n607), .B1(new_n606), .B2(G171), .ZN(G284));
  OAI21_X1  g183(.A(new_n607), .B1(new_n606), .B2(G171), .ZN(G321));
  NAND2_X1  g184(.A1(G299), .A2(new_n606), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(new_n606), .B2(G168), .ZN(G297));
  OAI21_X1  g186(.A(new_n610), .B1(new_n606), .B2(G168), .ZN(G280));
  AND2_X1   g187(.A1(new_n599), .A2(new_n604), .ZN(new_n613));
  INV_X1    g188(.A(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n614), .B2(G860), .ZN(G148));
  INV_X1    g190(.A(new_n558), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(new_n606), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n605), .A2(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(new_n606), .ZN(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g195(.A1(new_n462), .A2(new_n466), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT12), .Z(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT13), .Z(new_n623));
  INV_X1    g198(.A(G2100), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n623), .A2(new_n624), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n475), .A2(G135), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n477), .A2(G123), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n464), .A2(G111), .ZN(new_n629));
  OAI21_X1  g204(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n627), .B(new_n628), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(G2096), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n625), .A2(new_n626), .A3(new_n633), .ZN(G156));
  XNOR2_X1  g209(.A(G2451), .B(G2454), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT16), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(G2443), .B(G2446), .Z(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT15), .B(G2435), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2438), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2427), .B(G2430), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n643), .A2(KEYINPUT14), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(KEYINPUT76), .ZN(new_n645));
  INV_X1    g220(.A(KEYINPUT76), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n643), .A2(new_n646), .A3(KEYINPUT14), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n641), .A2(new_n642), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n639), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  AOI211_X1 g226(.A(new_n649), .B(new_n638), .C1(new_n645), .C2(new_n647), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n637), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(new_n647), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n646), .B1(new_n643), .B2(KEYINPUT14), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n650), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(new_n638), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n648), .A2(new_n650), .A3(new_n639), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n657), .A2(new_n636), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n653), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1341), .B(G1348), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n662), .A2(KEYINPUT77), .ZN(new_n663));
  INV_X1    g238(.A(KEYINPUT77), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n660), .A2(new_n664), .A3(new_n661), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n660), .A2(new_n661), .ZN(new_n667));
  INV_X1    g242(.A(G14), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(G401));
  INV_X1    g246(.A(KEYINPUT18), .ZN(new_n672));
  XOR2_X1   g247(.A(G2084), .B(G2090), .Z(new_n673));
  XNOR2_X1  g248(.A(G2067), .B(G2678), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(KEYINPUT17), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n673), .A2(new_n674), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n672), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(G2100), .ZN(new_n679));
  XOR2_X1   g254(.A(G2072), .B(G2078), .Z(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(new_n675), .B2(KEYINPUT18), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(new_n632), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n679), .A2(new_n682), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(G227));
  XOR2_X1   g261(.A(G1991), .B(G1996), .Z(new_n687));
  XNOR2_X1  g262(.A(G1971), .B(G1976), .ZN(new_n688));
  INV_X1    g263(.A(KEYINPUT19), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1956), .B(G2474), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1961), .B(G1966), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT20), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n691), .A2(new_n692), .ZN(new_n697));
  INV_X1    g272(.A(new_n693), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n697), .B1(new_n690), .B2(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n688), .B(KEYINPUT19), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(KEYINPUT78), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n699), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  NOR3_X1   g279(.A1(new_n696), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  AND2_X1   g280(.A1(new_n700), .A2(KEYINPUT78), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(new_n699), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n703), .B1(new_n707), .B2(new_n695), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n687), .B1(new_n705), .B2(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(G1981), .B(G1986), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n704), .B1(new_n696), .B2(new_n702), .ZN(new_n711));
  INV_X1    g286(.A(new_n687), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n707), .A2(new_n695), .A3(new_n703), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  AND3_X1   g289(.A1(new_n709), .A2(new_n710), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n710), .B1(new_n709), .B2(new_n714), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(G229));
  XNOR2_X1  g293(.A(KEYINPUT30), .B(G28), .ZN(new_n719));
  INV_X1    g294(.A(G29), .ZN(new_n720));
  OR2_X1    g295(.A1(KEYINPUT31), .A2(G11), .ZN(new_n721));
  NAND2_X1  g296(.A1(KEYINPUT31), .A2(G11), .ZN(new_n722));
  AOI22_X1  g297(.A1(new_n719), .A2(new_n720), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(new_n631), .B2(new_n720), .ZN(new_n724));
  NAND2_X1  g299(.A1(G168), .A2(G16), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT84), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n725), .B(new_n726), .C1(G16), .C2(G21), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(new_n726), .B2(new_n725), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n724), .B1(new_n728), .B2(G1966), .ZN(new_n729));
  INV_X1    g304(.A(G16), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G5), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G171), .B2(new_n730), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G1961), .ZN(new_n733));
  OAI211_X1 g308(.A(new_n729), .B(new_n733), .C1(G1966), .C2(new_n728), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT85), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n720), .A2(G35), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT88), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G162), .B2(new_n720), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT29), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n739), .A2(G2090), .ZN(new_n740));
  NOR2_X1   g315(.A1(G4), .A2(G16), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(new_n613), .B2(G16), .ZN(new_n742));
  AOI22_X1  g317(.A1(new_n740), .A2(KEYINPUT89), .B1(G1348), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(KEYINPUT89), .B2(new_n740), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n720), .A2(G26), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT28), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n475), .A2(G140), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT82), .Z(new_n748));
  OAI21_X1  g323(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n749));
  INV_X1    g324(.A(G116), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n749), .B1(new_n750), .B2(G2105), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(new_n477), .B2(G128), .ZN(new_n752));
  AND2_X1   g327(.A1(new_n748), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n746), .B1(new_n753), .B2(new_n720), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G2067), .ZN(new_n755));
  INV_X1    g330(.A(G160), .ZN(new_n756));
  NAND2_X1  g331(.A1(KEYINPUT24), .A2(G34), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT24), .ZN(new_n758));
  INV_X1    g333(.A(G34), .ZN(new_n759));
  AOI21_X1  g334(.A(G29), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  AOI22_X1  g335(.A1(new_n756), .A2(G29), .B1(new_n757), .B2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(G2084), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT86), .Z(new_n764));
  NAND2_X1  g339(.A1(new_n475), .A2(G141), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n477), .A2(G129), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n466), .A2(G105), .ZN(new_n767));
  NAND3_X1  g342(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT26), .Z(new_n769));
  NAND4_X1  g344(.A1(new_n765), .A2(new_n766), .A3(new_n767), .A4(new_n769), .ZN(new_n770));
  MUX2_X1   g345(.A(G32), .B(new_n770), .S(G29), .Z(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT27), .B(G1996), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT83), .B(KEYINPUT25), .ZN(new_n774));
  AND3_X1   g349(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n774), .A2(new_n775), .ZN(new_n777));
  AOI22_X1  g352(.A1(new_n776), .A2(new_n777), .B1(new_n475), .B2(G139), .ZN(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n780), .A2(new_n464), .ZN(new_n781));
  OAI21_X1  g356(.A(G29), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(G33), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(G29), .B2(new_n783), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n784), .A2(G2072), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n761), .A2(new_n762), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n784), .A2(G2072), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n773), .A2(new_n785), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  NOR3_X1   g363(.A1(new_n755), .A2(new_n764), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n720), .A2(G27), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G164), .B2(new_n720), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT87), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G2078), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n789), .B(new_n793), .C1(G1961), .C2(new_n732), .ZN(new_n794));
  XOR2_X1   g369(.A(KEYINPUT80), .B(G16), .Z(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n796), .A2(G19), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(new_n558), .B2(new_n796), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(G1341), .Z(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G1348), .B2(new_n742), .ZN(new_n800));
  NOR4_X1   g375(.A1(new_n735), .A2(new_n744), .A3(new_n794), .A4(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n796), .A2(G22), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G166), .B2(new_n796), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G1971), .ZN(new_n804));
  NOR2_X1   g379(.A1(G6), .A2(G16), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(new_n587), .B2(G16), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT32), .B(G1981), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n730), .A2(G23), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G288), .B2(G16), .ZN(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT33), .B(G1976), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n808), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n810), .A2(new_n811), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(new_n806), .B2(new_n807), .ZN(new_n814));
  NOR3_X1   g389(.A1(new_n804), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT34), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n815), .A2(new_n816), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n720), .A2(G25), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n477), .A2(G119), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT79), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n823));
  INV_X1    g398(.A(G107), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n823), .B1(new_n824), .B2(G2105), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n825), .B1(new_n475), .B2(G131), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n822), .A2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n819), .B1(new_n828), .B2(new_n720), .ZN(new_n829));
  XOR2_X1   g404(.A(KEYINPUT35), .B(G1991), .Z(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n829), .B(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n796), .A2(G24), .ZN(new_n833));
  INV_X1    g408(.A(G290), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n833), .B1(new_n834), .B2(new_n796), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(G1986), .ZN(new_n836));
  AOI211_X1 g411(.A(new_n832), .B(new_n836), .C1(KEYINPUT81), .C2(KEYINPUT36), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n817), .A2(new_n818), .A3(new_n837), .ZN(new_n838));
  NOR2_X1   g413(.A1(KEYINPUT81), .A2(KEYINPUT36), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n838), .A2(new_n839), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n739), .A2(G2090), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n842), .A2(KEYINPUT90), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(KEYINPUT90), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n795), .A2(G20), .ZN(new_n845));
  XOR2_X1   g420(.A(KEYINPUT91), .B(KEYINPUT23), .Z(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(new_n572), .B2(new_n730), .ZN(new_n848));
  INV_X1    g423(.A(G1956), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n843), .A2(new_n844), .A3(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT92), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n801), .A2(new_n840), .A3(new_n841), .A4(new_n852), .ZN(G150));
  INV_X1    g428(.A(G150), .ZN(G311));
  NAND2_X1  g429(.A1(new_n613), .A2(G559), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT38), .ZN(new_n856));
  NAND2_X1  g431(.A1(G80), .A2(G543), .ZN(new_n857));
  INV_X1    g432(.A(G67), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n857), .B1(new_n569), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(G651), .ZN(new_n860));
  NAND4_X1  g435(.A1(new_n551), .A2(G93), .A3(new_n509), .A4(new_n524), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n535), .A2(G55), .ZN(new_n862));
  AND3_X1   g437(.A1(new_n861), .A2(KEYINPUT93), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(KEYINPUT93), .B1(new_n861), .B2(new_n862), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n860), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(new_n616), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n861), .A2(new_n862), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT93), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n861), .A2(KEYINPUT93), .A3(new_n862), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n871), .A2(new_n558), .A3(new_n860), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n866), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n856), .B(new_n874), .ZN(new_n875));
  OR2_X1    g450(.A1(new_n875), .A2(KEYINPUT39), .ZN(new_n876));
  INV_X1    g451(.A(G860), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n875), .A2(KEYINPUT39), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n865), .A2(G860), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n880), .B(KEYINPUT37), .Z(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(G145));
  XNOR2_X1  g457(.A(new_n631), .B(KEYINPUT94), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(G160), .ZN(new_n884));
  INV_X1    g459(.A(G162), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n884), .B(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n770), .B1(new_n779), .B2(new_n781), .ZN(new_n887));
  AND2_X1   g462(.A1(new_n766), .A2(new_n769), .ZN(new_n888));
  AND2_X1   g463(.A1(new_n765), .A2(new_n767), .ZN(new_n889));
  INV_X1    g464(.A(new_n781), .ZN(new_n890));
  NAND4_X1  g465(.A1(new_n888), .A2(new_n889), .A3(new_n890), .A4(new_n778), .ZN(new_n891));
  AND2_X1   g466(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n491), .A2(new_n495), .ZN(new_n893));
  AOI21_X1  g468(.A(KEYINPUT69), .B1(new_n462), .B2(new_n483), .ZN(new_n894));
  INV_X1    g469(.A(new_n487), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n502), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n501), .B1(new_n462), .B2(new_n498), .ZN(new_n898));
  OAI21_X1  g473(.A(KEYINPUT95), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT95), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n500), .A2(new_n900), .A3(new_n502), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n896), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT96), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n500), .A2(new_n900), .A3(new_n502), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n900), .B1(new_n500), .B2(new_n502), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n496), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(KEYINPUT96), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n904), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n892), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n887), .A2(new_n891), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n911), .A2(new_n908), .A3(new_n904), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n748), .A2(new_n752), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n622), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n828), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n916), .B1(new_n822), .B2(new_n826), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n475), .A2(G142), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT97), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n920), .B(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n923));
  INV_X1    g498(.A(G118), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n923), .B1(new_n924), .B2(G2105), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n477), .A2(G130), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n922), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n917), .A2(new_n919), .A3(new_n929), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n827), .A2(new_n622), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n928), .B1(new_n931), .B2(new_n918), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n910), .A2(new_n753), .A3(new_n912), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n915), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n933), .B1(new_n915), .B2(new_n934), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n886), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(G37), .ZN(new_n938));
  AND2_X1   g513(.A1(new_n930), .A2(new_n932), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT98), .ZN(new_n940));
  INV_X1    g515(.A(new_n934), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n753), .B1(new_n910), .B2(new_n912), .ZN(new_n942));
  OAI211_X1 g517(.A(new_n939), .B(new_n940), .C1(new_n941), .C2(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n915), .A2(new_n933), .A3(new_n934), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n884), .B(G162), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n936), .A2(new_n940), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n937), .B(new_n938), .C1(new_n946), .C2(new_n947), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n948), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g524(.A(KEYINPUT100), .ZN(new_n950));
  XNOR2_X1  g525(.A(G288), .B(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(new_n587), .ZN(new_n952));
  XNOR2_X1  g527(.A(G288), .B(KEYINPUT100), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(G305), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(G303), .A2(new_n834), .ZN(new_n956));
  NAND2_X1  g531(.A1(G166), .A2(G290), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n955), .A2(new_n958), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n952), .A2(new_n954), .A3(new_n956), .A4(new_n957), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  AND2_X1   g537(.A1(KEYINPUT101), .A2(KEYINPUT42), .ZN(new_n963));
  NOR2_X1   g538(.A1(KEYINPUT101), .A2(KEYINPUT42), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n964), .B(KEYINPUT102), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  NOR3_X1   g541(.A1(new_n962), .A2(new_n963), .A3(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n963), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n965), .B1(new_n961), .B2(new_n968), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n613), .A2(new_n572), .ZN(new_n971));
  NAND2_X1  g546(.A1(G299), .A2(new_n605), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(KEYINPUT99), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT99), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n873), .B(new_n618), .ZN(new_n979));
  OR2_X1    g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(KEYINPUT41), .B1(new_n971), .B2(new_n972), .ZN(new_n981));
  AND3_X1   g556(.A1(new_n971), .A2(new_n972), .A3(KEYINPUT41), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n979), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n980), .A2(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n606), .B1(new_n970), .B2(new_n984), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n980), .B(new_n983), .C1(new_n967), .C2(new_n969), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n987), .A2(KEYINPUT103), .ZN(new_n988));
  INV_X1    g563(.A(new_n865), .ZN(new_n989));
  OAI21_X1  g564(.A(KEYINPUT103), .B1(new_n989), .B2(G868), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n990), .B1(new_n985), .B2(new_n986), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n988), .A2(new_n991), .ZN(G295));
  NOR2_X1   g567(.A1(new_n988), .A2(new_n991), .ZN(G331));
  XNOR2_X1  g568(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  AND3_X1   g570(.A1(new_n866), .A2(new_n872), .A3(G301), .ZN(new_n996));
  AOI21_X1  g571(.A(G301), .B1(new_n866), .B2(new_n872), .ZN(new_n997));
  NOR3_X1   g572(.A1(new_n996), .A2(new_n997), .A3(G286), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n873), .A2(G171), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n866), .A2(new_n872), .A3(G301), .ZN(new_n1000));
  AOI21_X1  g575(.A(G168), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n974), .B1(new_n998), .B2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n982), .A2(new_n981), .ZN(new_n1003));
  OAI21_X1  g578(.A(G286), .B1(new_n996), .B2(new_n997), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n999), .A2(G168), .A3(new_n1000), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1002), .A2(new_n962), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(new_n938), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n962), .B1(new_n1002), .B2(new_n1006), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n995), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1006), .ZN(new_n1011));
  AOI22_X1  g586(.A1(new_n1004), .A2(new_n1005), .B1(new_n975), .B2(new_n977), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n961), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1013), .A2(new_n938), .A3(new_n1007), .A4(new_n994), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1010), .A2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1015), .A2(KEYINPUT44), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT44), .ZN(new_n1017));
  OR3_X1    g592(.A1(new_n1008), .A2(new_n1009), .A3(new_n995), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1013), .A2(new_n938), .A3(new_n1007), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT43), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1017), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1016), .A2(new_n1021), .ZN(G397));
  INV_X1    g597(.A(KEYINPUT108), .ZN(new_n1023));
  INV_X1    g598(.A(G1384), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n904), .A2(new_n908), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT45), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G1996), .ZN(new_n1029));
  NAND2_X1  g604(.A1(G160), .A2(G40), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1028), .A2(new_n1029), .A3(new_n1031), .ZN(new_n1032));
  OR3_X1    g607(.A1(new_n1032), .A2(KEYINPUT105), .A3(new_n770), .ZN(new_n1033));
  OAI21_X1  g608(.A(KEYINPUT105), .B1(new_n1032), .B2(new_n770), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1036));
  INV_X1    g611(.A(G2067), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n753), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n914), .A2(G2067), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1036), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT107), .ZN(new_n1042));
  XNOR2_X1  g617(.A(new_n1041), .B(new_n1042), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1028), .A2(G1996), .A3(new_n770), .A4(new_n1031), .ZN(new_n1044));
  XNOR2_X1  g619(.A(new_n1044), .B(KEYINPUT106), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n827), .A2(new_n831), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n828), .A2(new_n830), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1036), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  AND4_X1   g623(.A1(new_n1035), .A2(new_n1043), .A3(new_n1045), .A4(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1036), .ZN(new_n1050));
  INV_X1    g625(.A(G1986), .ZN(new_n1051));
  XNOR2_X1  g626(.A(G290), .B(new_n1051), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1023), .B1(new_n1049), .B2(new_n1054), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1035), .A2(new_n1043), .A3(new_n1045), .A4(new_n1048), .ZN(new_n1056));
  NOR3_X1   g631(.A1(new_n1056), .A2(KEYINPUT108), .A3(new_n1053), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT109), .ZN(new_n1059));
  NOR3_X1   g634(.A1(new_n902), .A2(new_n1059), .A3(G1384), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT109), .B1(new_n907), .B2(new_n1024), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1031), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(G1976), .ZN(new_n1063));
  OAI21_X1  g638(.A(KEYINPUT111), .B1(G288), .B2(new_n1063), .ZN(new_n1064));
  AND2_X1   g639(.A1(new_n577), .A2(new_n578), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT111), .ZN(new_n1066));
  OAI21_X1  g641(.A(G651), .B1(new_n518), .B2(G74), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .A4(G1976), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1064), .A2(new_n1068), .ZN(new_n1069));
  AND3_X1   g644(.A1(new_n1062), .A2(G8), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT113), .ZN(new_n1071));
  INV_X1    g646(.A(G288), .ZN(new_n1072));
  XOR2_X1   g647(.A(KEYINPUT112), .B(G1976), .Z(new_n1073));
  NOR2_X1   g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1070), .B(new_n1071), .C1(KEYINPUT52), .C2(new_n1074), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1062), .A2(new_n1069), .A3(G8), .A4(new_n1074), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1062), .A2(new_n1069), .A3(new_n1071), .A4(G8), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1062), .A2(G8), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT114), .ZN(new_n1081));
  INV_X1    g656(.A(G1981), .ZN(new_n1082));
  INV_X1    g657(.A(new_n583), .ZN(new_n1083));
  INV_X1    g658(.A(new_n586), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1082), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NOR3_X1   g660(.A1(new_n583), .A2(new_n586), .A3(G1981), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1081), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n587), .A2(new_n1082), .ZN(new_n1088));
  OAI21_X1  g663(.A(G1981), .B1(new_n583), .B2(new_n586), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1088), .A2(KEYINPUT114), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT49), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1087), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1088), .A2(KEYINPUT49), .A3(new_n1089), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT115), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1080), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1087), .A2(new_n1090), .A3(new_n1094), .A4(new_n1091), .ZN(new_n1097));
  AOI22_X1  g672(.A1(new_n1075), .A2(new_n1079), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT110), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1059), .B1(new_n902), .B2(G1384), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT50), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n907), .A2(KEYINPUT109), .A3(new_n1024), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1100), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n504), .A2(new_n1024), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(KEYINPUT50), .ZN(new_n1106));
  AOI211_X1 g681(.A(G2090), .B(new_n1030), .C1(new_n1103), .C2(new_n1106), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n904), .A2(new_n908), .A3(KEYINPUT45), .A4(new_n1024), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1030), .B1(new_n1104), .B2(new_n1026), .ZN(new_n1109));
  AOI21_X1  g684(.A(G1971), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1099), .B1(new_n1107), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1112));
  INV_X1    g687(.A(G2090), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1112), .A2(new_n1113), .A3(new_n1031), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1110), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1114), .A2(new_n1115), .A3(KEYINPUT110), .ZN(new_n1116));
  NAND3_X1  g691(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT55), .ZN(new_n1118));
  INV_X1    g693(.A(G8), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1118), .B1(G166), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1117), .A2(new_n1120), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1111), .A2(G8), .A3(new_n1116), .A4(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1100), .A2(KEYINPUT50), .A3(new_n1102), .ZN(new_n1123));
  OAI21_X1  g698(.A(KEYINPUT116), .B1(new_n1104), .B2(KEYINPUT50), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT116), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n504), .A2(new_n1125), .A3(new_n1101), .A4(new_n1024), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1123), .A2(new_n1127), .A3(new_n1031), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1128), .A2(G2090), .ZN(new_n1129));
  OAI21_X1  g704(.A(G8), .B1(new_n1129), .B2(new_n1110), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1121), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  AND3_X1   g707(.A1(new_n1098), .A2(new_n1122), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT54), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1030), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(G1961), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT53), .ZN(new_n1138));
  INV_X1    g713(.A(G2078), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1108), .A2(new_n1139), .A3(new_n1109), .ZN(new_n1140));
  AOI22_X1  g715(.A1(new_n1136), .A2(new_n1137), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT122), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1100), .A2(new_n1026), .A3(new_n1102), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1030), .B1(new_n1105), .B2(KEYINPUT45), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1142), .B1(new_n1145), .B2(G2078), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1143), .A2(new_n1144), .A3(KEYINPUT122), .A4(new_n1139), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1146), .A2(KEYINPUT53), .A3(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(G301), .B1(new_n1141), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1140), .A2(new_n1138), .ZN(new_n1150));
  INV_X1    g725(.A(new_n470), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(KEYINPUT123), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1139), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT123), .ZN(new_n1154));
  AOI211_X1 g729(.A(new_n1153), .B(new_n465), .C1(new_n1154), .C2(new_n470), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1027), .A2(new_n1108), .A3(new_n1152), .A4(new_n1155), .ZN(new_n1156));
  OAI211_X1 g731(.A(new_n1150), .B(new_n1156), .C1(G1961), .C2(new_n1135), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1157), .A2(G171), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1134), .B1(new_n1149), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT121), .ZN(new_n1160));
  AOI21_X1  g735(.A(G1966), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1030), .A2(G2084), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1163), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n1161), .A2(new_n1164), .A3(G286), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n1160), .B(KEYINPUT51), .C1(new_n1165), .C2(new_n1119), .ZN(new_n1166));
  OAI211_X1 g741(.A(G8), .B(G286), .C1(new_n1161), .C2(new_n1164), .ZN(new_n1167));
  INV_X1    g742(.A(G1966), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1145), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1112), .A2(new_n1162), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1169), .A2(new_n1170), .A3(G168), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT51), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1119), .B1(KEYINPUT121), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1160), .A2(KEYINPUT51), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1171), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1166), .A2(new_n1167), .A3(new_n1175), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1134), .B1(new_n1157), .B2(G171), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1141), .A2(new_n1148), .A3(G301), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1133), .A2(new_n1159), .A3(new_n1176), .A4(new_n1179), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1030), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1181), .A2(new_n1037), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1182), .A2(KEYINPUT119), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT119), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1184), .B1(new_n1181), .B2(new_n1037), .ZN(new_n1185));
  OAI22_X1  g760(.A1(new_n1183), .A2(new_n1185), .B1(G1348), .B2(new_n1135), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1186), .A2(new_n613), .ZN(new_n1187));
  AND2_X1   g762(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1188));
  XNOR2_X1  g763(.A(KEYINPUT56), .B(G2072), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1128), .A2(new_n849), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g767(.A(new_n572), .B(KEYINPUT57), .ZN(new_n1193));
  INV_X1    g768(.A(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1192), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1187), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT118), .ZN(new_n1197));
  AOI22_X1  g772(.A1(new_n1188), .A2(new_n1189), .B1(new_n1128), .B2(new_n849), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1197), .B1(new_n1198), .B2(new_n1193), .ZN(new_n1199));
  AND4_X1   g774(.A1(new_n1197), .A2(new_n1190), .A3(new_n1191), .A4(new_n1193), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1196), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1195), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1202));
  INV_X1    g777(.A(KEYINPUT61), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  XOR2_X1   g779(.A(KEYINPUT120), .B(KEYINPUT60), .Z(new_n1205));
  INV_X1    g780(.A(new_n1205), .ZN(new_n1206));
  AOI21_X1  g781(.A(new_n613), .B1(new_n1186), .B2(KEYINPUT60), .ZN(new_n1207));
  XNOR2_X1  g782(.A(new_n1182), .B(KEYINPUT119), .ZN(new_n1208));
  OR2_X1    g783(.A1(new_n1135), .A2(G1348), .ZN(new_n1209));
  AOI21_X1  g784(.A(new_n605), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g785(.A(new_n1206), .B1(new_n1207), .B2(new_n1210), .ZN(new_n1211));
  INV_X1    g786(.A(KEYINPUT60), .ZN(new_n1212));
  AOI21_X1  g787(.A(new_n1212), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1213));
  OAI211_X1 g788(.A(new_n1187), .B(new_n1205), .C1(new_n1213), .C2(new_n613), .ZN(new_n1214));
  AOI21_X1  g789(.A(new_n1203), .B1(new_n1192), .B2(new_n1194), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1198), .A2(new_n1193), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1217));
  NOR2_X1   g792(.A1(new_n1217), .A2(G1996), .ZN(new_n1218));
  XNOR2_X1  g793(.A(KEYINPUT58), .B(G1341), .ZN(new_n1219));
  NOR2_X1   g794(.A1(new_n1181), .A2(new_n1219), .ZN(new_n1220));
  OAI21_X1  g795(.A(new_n558), .B1(new_n1218), .B2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1221), .A2(KEYINPUT59), .ZN(new_n1222));
  INV_X1    g797(.A(KEYINPUT59), .ZN(new_n1223));
  OAI211_X1 g798(.A(new_n1223), .B(new_n558), .C1(new_n1218), .C2(new_n1220), .ZN(new_n1224));
  AOI22_X1  g799(.A1(new_n1215), .A2(new_n1216), .B1(new_n1222), .B2(new_n1224), .ZN(new_n1225));
  NAND4_X1  g800(.A1(new_n1204), .A2(new_n1211), .A3(new_n1214), .A4(new_n1225), .ZN(new_n1226));
  AOI21_X1  g801(.A(new_n1180), .B1(new_n1201), .B2(new_n1226), .ZN(new_n1227));
  OAI211_X1 g802(.A(G8), .B(G168), .C1(new_n1161), .C2(new_n1164), .ZN(new_n1228));
  INV_X1    g803(.A(new_n1228), .ZN(new_n1229));
  NAND4_X1  g804(.A1(new_n1098), .A2(new_n1122), .A3(new_n1132), .A4(new_n1229), .ZN(new_n1230));
  INV_X1    g805(.A(KEYINPUT63), .ZN(new_n1231));
  NAND2_X1  g806(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  NAND3_X1  g807(.A1(new_n1111), .A2(G8), .A3(new_n1116), .ZN(new_n1233));
  INV_X1    g808(.A(KEYINPUT117), .ZN(new_n1234));
  NAND3_X1  g809(.A1(new_n1233), .A2(new_n1234), .A3(new_n1131), .ZN(new_n1235));
  NAND2_X1  g810(.A1(new_n1131), .A2(new_n1234), .ZN(new_n1236));
  NAND4_X1  g811(.A1(new_n1236), .A2(G8), .A3(new_n1111), .A4(new_n1116), .ZN(new_n1237));
  NOR2_X1   g812(.A1(new_n1228), .A2(new_n1231), .ZN(new_n1238));
  NAND4_X1  g813(.A1(new_n1235), .A2(new_n1098), .A3(new_n1237), .A4(new_n1238), .ZN(new_n1239));
  NAND2_X1  g814(.A1(new_n1232), .A2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g815(.A1(new_n1175), .A2(new_n1167), .ZN(new_n1241));
  AOI21_X1  g816(.A(new_n1174), .B1(new_n1171), .B2(new_n1173), .ZN(new_n1242));
  OAI21_X1  g817(.A(KEYINPUT62), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  INV_X1    g818(.A(KEYINPUT62), .ZN(new_n1244));
  NAND4_X1  g819(.A1(new_n1166), .A2(new_n1244), .A3(new_n1167), .A4(new_n1175), .ZN(new_n1245));
  NAND4_X1  g820(.A1(new_n1133), .A2(new_n1243), .A3(new_n1149), .A4(new_n1245), .ZN(new_n1246));
  NAND2_X1  g821(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1247));
  NAND3_X1  g822(.A1(new_n1247), .A2(new_n1063), .A3(new_n1072), .ZN(new_n1248));
  NAND2_X1  g823(.A1(new_n1248), .A2(new_n1088), .ZN(new_n1249));
  INV_X1    g824(.A(new_n1080), .ZN(new_n1250));
  INV_X1    g825(.A(new_n1122), .ZN(new_n1251));
  AOI22_X1  g826(.A1(new_n1249), .A2(new_n1250), .B1(new_n1251), .B2(new_n1098), .ZN(new_n1252));
  NAND3_X1  g827(.A1(new_n1240), .A2(new_n1246), .A3(new_n1252), .ZN(new_n1253));
  OAI21_X1  g828(.A(new_n1058), .B1(new_n1227), .B2(new_n1253), .ZN(new_n1254));
  NAND4_X1  g829(.A1(new_n1035), .A2(new_n1043), .A3(new_n1046), .A4(new_n1045), .ZN(new_n1255));
  AOI21_X1  g830(.A(new_n1050), .B1(new_n1255), .B2(new_n1038), .ZN(new_n1256));
  INV_X1    g831(.A(new_n1256), .ZN(new_n1257));
  NAND3_X1  g832(.A1(new_n1036), .A2(new_n1051), .A3(new_n834), .ZN(new_n1258));
  XNOR2_X1  g833(.A(new_n1258), .B(KEYINPUT48), .ZN(new_n1259));
  XNOR2_X1  g834(.A(KEYINPUT124), .B(KEYINPUT47), .ZN(new_n1260));
  XNOR2_X1  g835(.A(new_n1032), .B(KEYINPUT46), .ZN(new_n1261));
  OAI21_X1  g836(.A(new_n1036), .B1(new_n770), .B2(new_n1040), .ZN(new_n1262));
  AOI21_X1  g837(.A(new_n1260), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  INV_X1    g838(.A(new_n1263), .ZN(new_n1264));
  NAND3_X1  g839(.A1(new_n1261), .A2(new_n1262), .A3(new_n1260), .ZN(new_n1265));
  AOI22_X1  g840(.A1(new_n1049), .A2(new_n1259), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  NAND3_X1  g841(.A1(new_n1257), .A2(new_n1266), .A3(KEYINPUT125), .ZN(new_n1267));
  INV_X1    g842(.A(KEYINPUT125), .ZN(new_n1268));
  INV_X1    g843(.A(new_n1259), .ZN(new_n1269));
  INV_X1    g844(.A(new_n1265), .ZN(new_n1270));
  OAI22_X1  g845(.A1(new_n1056), .A2(new_n1269), .B1(new_n1270), .B2(new_n1263), .ZN(new_n1271));
  OAI21_X1  g846(.A(new_n1268), .B1(new_n1271), .B2(new_n1256), .ZN(new_n1272));
  NAND2_X1  g847(.A1(new_n1267), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g848(.A1(new_n1254), .A2(new_n1273), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g849(.A(KEYINPUT126), .B1(new_n685), .B2(G319), .ZN(new_n1276));
  INV_X1    g850(.A(KEYINPUT126), .ZN(new_n1277));
  AOI211_X1 g851(.A(new_n1277), .B(new_n460), .C1(new_n683), .C2(new_n684), .ZN(new_n1278));
  NOR2_X1   g852(.A1(new_n1276), .A2(new_n1278), .ZN(new_n1279));
  OAI21_X1  g853(.A(new_n1279), .B1(new_n715), .B2(new_n716), .ZN(new_n1280));
  AOI21_X1  g854(.A(new_n1280), .B1(new_n666), .B2(new_n669), .ZN(new_n1281));
  NAND2_X1  g855(.A1(new_n1281), .A2(new_n948), .ZN(new_n1282));
  INV_X1    g856(.A(new_n1282), .ZN(new_n1283));
  AOI21_X1  g857(.A(KEYINPUT127), .B1(new_n1015), .B2(new_n1283), .ZN(new_n1284));
  INV_X1    g858(.A(KEYINPUT127), .ZN(new_n1285));
  AOI211_X1 g859(.A(new_n1285), .B(new_n1282), .C1(new_n1010), .C2(new_n1014), .ZN(new_n1286));
  NOR2_X1   g860(.A1(new_n1284), .A2(new_n1286), .ZN(G308));
  NAND2_X1  g861(.A1(new_n1015), .A2(new_n1283), .ZN(G225));
endmodule


