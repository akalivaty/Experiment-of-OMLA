//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 0 0 0 0 1 0 0 1 0 1 0 0 0 0 1 1 1 1 1 0 0 0 0 0 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 1 0 1 1 0 0 1 1 1 0 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:53 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n596,
    new_n597, new_n598, new_n599, new_n600, new_n601, new_n602, new_n603,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n652, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920;
  INV_X1    g000(.A(G104), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT82), .B1(new_n187), .B2(G107), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT82), .ZN(new_n189));
  INV_X1    g003(.A(G107), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(G104), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n187), .A2(G107), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n188), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G101), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(KEYINPUT83), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT83), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n193), .A2(new_n196), .A3(G101), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  OAI21_X1  g012(.A(KEYINPUT3), .B1(new_n187), .B2(G107), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT3), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n200), .A2(new_n190), .A3(G104), .ZN(new_n201));
  INV_X1    g015(.A(G101), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n199), .A2(new_n201), .A3(new_n202), .A4(new_n192), .ZN(new_n203));
  XNOR2_X1  g017(.A(new_n203), .B(KEYINPUT81), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n198), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G146), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G143), .ZN(new_n207));
  INV_X1    g021(.A(G143), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g024(.A(KEYINPUT66), .B(G128), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT1), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n213), .B1(G143), .B2(new_n206), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n210), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(new_n210), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n216), .A2(new_n213), .A3(G128), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n205), .A2(KEYINPUT10), .A3(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT81), .ZN(new_n220));
  XNOR2_X1  g034(.A(new_n203), .B(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n199), .A2(new_n201), .A3(new_n192), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT80), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n199), .A2(new_n201), .A3(KEYINPUT80), .A4(new_n192), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n224), .A2(G101), .A3(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n221), .A2(KEYINPUT4), .A3(new_n226), .ZN(new_n227));
  OR2_X1    g041(.A1(new_n226), .A2(KEYINPUT4), .ZN(new_n228));
  NAND2_X1  g042(.A1(KEYINPUT0), .A2(G128), .ZN(new_n229));
  OR2_X1    g043(.A1(KEYINPUT0), .A2(G128), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n216), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n210), .B1(KEYINPUT0), .B2(G128), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n227), .A2(new_n228), .A3(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G128), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n210), .B1(new_n214), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n217), .A2(new_n237), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n221), .A2(new_n195), .A3(new_n197), .A4(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT10), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT11), .ZN(new_n242));
  INV_X1    g056(.A(G137), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G134), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT64), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n242), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  AOI211_X1 g060(.A(KEYINPUT64), .B(KEYINPUT11), .C1(new_n243), .C2(G134), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G131), .ZN(new_n249));
  INV_X1    g063(.A(G134), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G137), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n248), .A2(KEYINPUT65), .A3(new_n249), .A4(new_n251), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n245), .B1(new_n250), .B2(G137), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT11), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n244), .A2(new_n245), .A3(new_n242), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n254), .A2(new_n255), .A3(new_n249), .A4(new_n251), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT65), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n248), .A2(new_n251), .ZN(new_n259));
  AOI22_X1  g073(.A1(new_n252), .A2(new_n258), .B1(new_n259), .B2(G131), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n219), .A2(new_n235), .A3(new_n241), .A4(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(G110), .B(G140), .ZN(new_n262));
  INV_X1    g076(.A(G953), .ZN(new_n263));
  AND2_X1   g077(.A1(new_n263), .A2(G227), .ZN(new_n264));
  XOR2_X1   g078(.A(new_n262), .B(new_n264), .Z(new_n265));
  NAND2_X1  g079(.A1(new_n261), .A2(new_n265), .ZN(new_n266));
  OR2_X1    g080(.A1(new_n266), .A2(KEYINPUT85), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT84), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT12), .ZN(new_n269));
  INV_X1    g083(.A(new_n218), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n270), .B1(new_n198), .B2(new_n204), .ZN(new_n271));
  AND2_X1   g085(.A1(new_n271), .A2(new_n239), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n268), .B(new_n269), .C1(new_n272), .C2(new_n260), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n260), .B1(new_n271), .B2(new_n239), .ZN(new_n274));
  OAI21_X1  g088(.A(KEYINPUT84), .B1(new_n274), .B2(KEYINPUT12), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(KEYINPUT12), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n273), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n266), .A2(KEYINPUT85), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n267), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n219), .A2(new_n235), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n260), .B1(new_n280), .B2(new_n241), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  AND2_X1   g096(.A1(new_n282), .A2(new_n261), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n279), .B1(new_n283), .B2(new_n265), .ZN(new_n284));
  INV_X1    g098(.A(G469), .ZN(new_n285));
  INV_X1    g099(.A(G902), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n277), .A2(new_n261), .ZN(new_n288));
  INV_X1    g102(.A(new_n265), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n281), .A2(new_n266), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n290), .A2(G469), .A3(new_n292), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n287), .B(new_n293), .C1(new_n285), .C2(new_n286), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT86), .ZN(new_n295));
  XOR2_X1   g109(.A(KEYINPUT9), .B(G234), .Z(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(G221), .B1(new_n297), .B2(G902), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n294), .A2(new_n295), .A3(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n295), .B1(new_n294), .B2(new_n298), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT77), .B(G125), .ZN(new_n303));
  NOR3_X1   g117(.A1(new_n303), .A2(KEYINPUT16), .A3(G140), .ZN(new_n304));
  INV_X1    g118(.A(new_n303), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G140), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n306), .B1(G125), .B2(G140), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n304), .B1(new_n307), .B2(KEYINPUT16), .ZN(new_n308));
  AND2_X1   g122(.A1(new_n308), .A2(G146), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n308), .A2(G146), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  XOR2_X1   g125(.A(KEYINPUT69), .B(G237), .Z(new_n312));
  NOR2_X1   g126(.A1(new_n312), .A2(G953), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G214), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(new_n208), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n313), .A2(G143), .A3(G214), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n317), .A2(KEYINPUT17), .A3(G131), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT91), .B1(new_n317), .B2(G131), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n317), .A2(G131), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT91), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n315), .A2(new_n321), .A3(new_n249), .A4(new_n316), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n319), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n311), .B(new_n318), .C1(new_n323), .C2(KEYINPUT17), .ZN(new_n324));
  XNOR2_X1  g138(.A(G113), .B(G122), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n325), .B(new_n187), .ZN(new_n326));
  XOR2_X1   g140(.A(G125), .B(G140), .Z(new_n327));
  OR2_X1    g141(.A1(new_n327), .A2(G146), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n328), .B1(new_n307), .B2(new_n206), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT18), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n330), .A2(new_n249), .ZN(new_n331));
  OAI221_X1 g145(.A(new_n329), .B1(new_n317), .B2(new_n331), .C1(new_n320), .C2(new_n330), .ZN(new_n332));
  AND3_X1   g146(.A1(new_n324), .A2(new_n326), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n326), .B1(new_n324), .B2(new_n332), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n286), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT92), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT92), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n337), .B(new_n286), .C1(new_n333), .C2(new_n334), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n336), .A2(G475), .A3(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n309), .ZN(new_n340));
  MUX2_X1   g154(.A(new_n327), .B(new_n307), .S(KEYINPUT19), .Z(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n323), .B(new_n340), .C1(G146), .C2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n332), .ZN(new_n344));
  INV_X1    g158(.A(new_n326), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n324), .A2(new_n326), .A3(new_n332), .ZN(new_n347));
  AOI21_X1  g161(.A(G475), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n286), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT20), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n348), .A2(KEYINPUT20), .A3(new_n286), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n339), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n211), .A2(new_n208), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n354), .B1(G128), .B2(new_n208), .ZN(new_n355));
  OAI21_X1  g169(.A(G134), .B1(new_n354), .B2(KEYINPUT13), .ZN(new_n356));
  XOR2_X1   g170(.A(new_n355), .B(new_n356), .Z(new_n357));
  XNOR2_X1  g171(.A(G116), .B(G122), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n358), .B(new_n190), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  OR2_X1    g174(.A1(new_n355), .A2(G134), .ZN(new_n361));
  INV_X1    g175(.A(G116), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(KEYINPUT14), .A3(G122), .ZN(new_n363));
  INV_X1    g177(.A(new_n358), .ZN(new_n364));
  OAI211_X1 g178(.A(G107), .B(new_n363), .C1(new_n364), .C2(KEYINPUT14), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n355), .A2(G134), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n358), .A2(new_n190), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n361), .A2(new_n365), .A3(new_n366), .A4(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n360), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(G217), .ZN(new_n370));
  NOR3_X1   g184(.A1(new_n297), .A2(new_n370), .A3(G953), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n360), .A2(new_n368), .A3(new_n371), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT93), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(new_n376), .A3(new_n286), .ZN(new_n377));
  INV_X1    g191(.A(G478), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n378), .A2(KEYINPUT15), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n377), .B(new_n379), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n353), .A2(new_n380), .ZN(new_n381));
  AND2_X1   g195(.A1(new_n302), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n313), .A2(G210), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n383), .B(G101), .ZN(new_n384));
  XNOR2_X1  g198(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n384), .B(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n252), .A2(new_n258), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n259), .A2(G131), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n234), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT68), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n392), .B1(new_n362), .B2(G119), .ZN(new_n393));
  INV_X1    g207(.A(G119), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n394), .A2(KEYINPUT68), .A3(G116), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n393), .B(new_n395), .C1(G116), .C2(new_n394), .ZN(new_n396));
  XNOR2_X1  g210(.A(KEYINPUT2), .B(G113), .ZN(new_n397));
  XOR2_X1   g211(.A(new_n396), .B(new_n397), .Z(new_n398));
  AOI21_X1  g212(.A(new_n249), .B1(new_n251), .B2(new_n244), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n399), .B1(new_n215), .B2(new_n217), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n388), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n391), .A2(new_n398), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n403), .A2(KEYINPUT28), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT67), .ZN(new_n405));
  INV_X1    g219(.A(new_n258), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n256), .A2(new_n257), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n400), .B(new_n405), .C1(new_n406), .C2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n233), .B1(new_n388), .B2(new_n389), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n405), .B1(new_n388), .B2(new_n400), .ZN(new_n411));
  NOR3_X1   g225(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(KEYINPUT71), .B1(new_n412), .B2(new_n398), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n401), .A2(KEYINPUT67), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n391), .A2(new_n414), .A3(new_n408), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT71), .ZN(new_n416));
  INV_X1    g230(.A(new_n398), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n413), .A2(new_n402), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n404), .B1(new_n419), .B2(KEYINPUT28), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT29), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n387), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT28), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n391), .A2(new_n401), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n417), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n423), .B1(new_n425), .B2(new_n402), .ZN(new_n426));
  OR2_X1    g240(.A1(new_n426), .A2(KEYINPUT75), .ZN(new_n427));
  OAI21_X1  g241(.A(KEYINPUT75), .B1(new_n426), .B2(new_n404), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n422), .B1(new_n421), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT30), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n415), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n391), .A2(KEYINPUT30), .A3(new_n401), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n433), .A2(new_n417), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(new_n402), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n436), .A2(new_n386), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n431), .B1(KEYINPUT29), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(G472), .B1(new_n439), .B2(G902), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT32), .ZN(new_n441));
  OAI21_X1  g255(.A(KEYINPUT72), .B1(new_n420), .B2(new_n386), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n386), .A2(new_n402), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(KEYINPUT70), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT70), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n386), .A2(new_n445), .A3(new_n402), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n435), .A2(new_n444), .A3(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT31), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n435), .A2(new_n444), .A3(KEYINPUT31), .A4(new_n446), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT72), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n415), .A2(new_n417), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n403), .B1(new_n453), .B2(KEYINPUT71), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n423), .B1(new_n454), .B2(new_n418), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n452), .B(new_n387), .C1(new_n455), .C2(new_n404), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n442), .A2(new_n451), .A3(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT73), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n442), .A2(new_n456), .A3(new_n451), .A4(KEYINPUT73), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g275(.A1(G472), .A2(G902), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n462), .B(KEYINPUT74), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n441), .B1(new_n461), .B2(new_n464), .ZN(new_n465));
  AOI211_X1 g279(.A(KEYINPUT32), .B(new_n463), .C1(new_n459), .C2(new_n460), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n440), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  XNOR2_X1  g281(.A(KEYINPUT22), .B(G137), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n263), .A2(G221), .A3(G234), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n468), .B(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n394), .A2(G128), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n472), .B1(new_n211), .B2(new_n394), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n473), .B(KEYINPUT76), .ZN(new_n474));
  XOR2_X1   g288(.A(KEYINPUT24), .B(G110), .Z(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(G110), .ZN(new_n477));
  AOI21_X1  g291(.A(KEYINPUT23), .B1(new_n236), .B2(G119), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n478), .B1(new_n473), .B2(KEYINPUT23), .ZN(new_n479));
  OAI221_X1 g293(.A(new_n476), .B1(new_n477), .B2(new_n479), .C1(new_n309), .C2(new_n310), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n477), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n481), .B1(new_n474), .B2(new_n475), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n340), .A2(new_n482), .A3(new_n328), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n484), .A2(KEYINPUT78), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n484), .A2(KEYINPUT78), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n471), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n480), .A2(new_n483), .A3(new_n470), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n487), .A2(new_n286), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT25), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n370), .B1(G234), .B2(new_n286), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT25), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n487), .A2(new_n492), .A3(new_n286), .A4(new_n488), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n490), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  AND2_X1   g308(.A1(new_n487), .A2(new_n488), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n491), .A2(G902), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n496), .B(KEYINPUT79), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  AND2_X1   g313(.A1(new_n494), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(G952), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n501), .A2(G953), .ZN(new_n502));
  NAND2_X1  g316(.A1(G234), .A2(G237), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(KEYINPUT21), .B(G898), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n505), .B(KEYINPUT94), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n503), .A2(G902), .A3(G953), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n504), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(G214), .B1(G237), .B2(G902), .ZN(new_n510));
  XOR2_X1   g324(.A(new_n510), .B(KEYINPUT87), .Z(new_n511));
  NAND2_X1  g325(.A1(new_n218), .A2(new_n303), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n512), .B1(new_n303), .B2(new_n233), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n263), .A2(G224), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n513), .B(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n417), .A2(new_n227), .A3(new_n228), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT5), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n517), .A2(new_n394), .A3(G116), .ZN(new_n518));
  OAI211_X1 g332(.A(G113), .B(new_n518), .C1(new_n396), .C2(new_n517), .ZN(new_n519));
  OR2_X1    g333(.A1(new_n396), .A2(new_n397), .ZN(new_n520));
  AND2_X1   g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n205), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n516), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT88), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  XOR2_X1   g339(.A(G110), .B(G122), .Z(new_n526));
  NAND3_X1  g340(.A1(new_n516), .A2(KEYINPUT88), .A3(new_n522), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  OR2_X1    g342(.A1(new_n523), .A2(new_n526), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n528), .A2(KEYINPUT6), .A3(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT6), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n525), .A2(new_n531), .A3(new_n526), .A4(new_n527), .ZN(new_n532));
  AND2_X1   g346(.A1(new_n532), .A2(KEYINPUT89), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n532), .A2(KEYINPUT89), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n515), .B(new_n530), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(KEYINPUT7), .B1(new_n263), .B2(G224), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n515), .B(new_n536), .ZN(new_n537));
  XOR2_X1   g351(.A(new_n205), .B(new_n521), .Z(new_n538));
  XNOR2_X1  g352(.A(new_n526), .B(KEYINPUT8), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n537), .B(new_n529), .C1(new_n538), .C2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n535), .A2(new_n286), .A3(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(G210), .B1(G237), .B2(G902), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n535), .A2(new_n286), .A3(new_n542), .A4(new_n540), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n511), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(KEYINPUT90), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT90), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n509), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n382), .A2(new_n467), .A3(new_n500), .A4(new_n551), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n552), .B(G101), .ZN(G3));
  AOI21_X1  g367(.A(new_n463), .B1(new_n459), .B2(new_n460), .ZN(new_n554));
  AOI21_X1  g368(.A(G902), .B1(new_n459), .B2(new_n460), .ZN(new_n555));
  OR2_X1    g369(.A1(new_n555), .A2(KEYINPUT95), .ZN(new_n556));
  INV_X1    g370(.A(G472), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n557), .B1(new_n555), .B2(KEYINPUT95), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n554), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n559), .A2(new_n500), .A3(new_n302), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n546), .A2(new_n508), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n375), .A2(KEYINPUT33), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT33), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n373), .A2(new_n564), .A3(new_n374), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n563), .A2(G478), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(G478), .A2(G902), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n375), .A2(new_n378), .A3(new_n286), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n353), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n562), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n561), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n573), .B(G104), .ZN(new_n574));
  XOR2_X1   g388(.A(KEYINPUT96), .B(KEYINPUT34), .Z(new_n575));
  XNOR2_X1  g389(.A(new_n574), .B(new_n575), .ZN(G6));
  INV_X1    g390(.A(new_n353), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n380), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n562), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n561), .A2(new_n579), .ZN(new_n580));
  XOR2_X1   g394(.A(KEYINPUT35), .B(G107), .Z(new_n581));
  XNOR2_X1  g395(.A(new_n580), .B(new_n581), .ZN(G9));
  INV_X1    g396(.A(new_n301), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n485), .A2(new_n486), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n471), .A2(KEYINPUT36), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n585), .B(KEYINPUT97), .ZN(new_n586));
  AND2_X1   g400(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n584), .A2(new_n586), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n498), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n494), .A2(new_n589), .ZN(new_n590));
  AND4_X1   g404(.A1(new_n583), .A2(new_n299), .A3(new_n381), .A4(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n559), .A2(new_n591), .A3(new_n551), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(G110), .ZN(new_n593));
  XOR2_X1   g407(.A(KEYINPUT98), .B(KEYINPUT37), .Z(new_n594));
  XNOR2_X1  g408(.A(new_n593), .B(new_n594), .ZN(G12));
  INV_X1    g409(.A(new_n590), .ZN(new_n596));
  NOR3_X1   g410(.A1(new_n300), .A2(new_n596), .A3(new_n301), .ZN(new_n597));
  XOR2_X1   g411(.A(new_n504), .B(KEYINPUT99), .Z(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n599), .B1(G900), .B2(new_n507), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n578), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n467), .A2(new_n597), .A3(new_n546), .A4(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(G128), .ZN(G30));
  INV_X1    g418(.A(KEYINPUT101), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT100), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n461), .A2(new_n464), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(KEYINPUT32), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n554), .A2(new_n441), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n425), .A2(new_n402), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(new_n387), .ZN(new_n612));
  AND2_X1   g426(.A1(new_n447), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g427(.A(G472), .B1(new_n613), .B2(G902), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n606), .B1(new_n610), .B2(new_n614), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n606), .B(new_n614), .C1(new_n465), .C2(new_n466), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n605), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n614), .B1(new_n465), .B2(new_n466), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(KEYINPUT100), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n620), .A2(KEYINPUT101), .A3(new_n616), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  XOR2_X1   g437(.A(new_n600), .B(KEYINPUT39), .Z(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n302), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(KEYINPUT40), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n544), .A2(new_n545), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(KEYINPUT38), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n511), .ZN(new_n632));
  AND3_X1   g446(.A1(new_n353), .A2(new_n632), .A3(new_n380), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n596), .ZN(new_n634));
  XOR2_X1   g448(.A(new_n634), .B(KEYINPUT102), .Z(new_n635));
  NAND3_X1  g449(.A1(new_n623), .A2(new_n631), .A3(new_n635), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT103), .B(G143), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G45));
  NOR2_X1   g452(.A1(new_n571), .A2(new_n601), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n467), .A2(new_n597), .A3(new_n546), .A4(new_n639), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT104), .B(G146), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G48));
  INV_X1    g456(.A(new_n287), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n285), .B1(new_n284), .B2(new_n286), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n298), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n467), .A2(new_n500), .A3(new_n572), .A4(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(KEYINPUT105), .ZN(new_n649));
  XNOR2_X1  g463(.A(KEYINPUT41), .B(G113), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G15));
  NAND4_X1  g465(.A1(new_n467), .A2(new_n500), .A3(new_n579), .A4(new_n647), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G116), .ZN(G18));
  AND2_X1   g467(.A1(new_n381), .A2(new_n590), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n646), .A2(new_n509), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n467), .A2(new_n546), .A3(new_n654), .A4(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G119), .ZN(G21));
  INV_X1    g471(.A(new_n555), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n386), .B1(new_n429), .B2(KEYINPUT106), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n659), .B1(KEYINPUT106), .B2(new_n429), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n451), .ZN(new_n661));
  AOI22_X1  g475(.A1(new_n658), .A2(G472), .B1(new_n464), .B2(new_n661), .ZN(new_n662));
  AND2_X1   g476(.A1(new_n633), .A2(new_n628), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n662), .A2(new_n500), .A3(new_n663), .A4(new_n655), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G122), .ZN(G24));
  NOR2_X1   g479(.A1(new_n547), .A2(new_n646), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n662), .A2(new_n590), .A3(new_n639), .A4(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G125), .ZN(G27));
  INV_X1    g482(.A(new_n639), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n628), .A2(new_n511), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n294), .A2(new_n298), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n672), .A2(new_n500), .A3(new_n467), .A4(new_n674), .ZN(new_n675));
  OR2_X1    g489(.A1(KEYINPUT107), .A2(KEYINPUT42), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(new_n249), .ZN(G33));
  NAND4_X1  g492(.A1(new_n467), .A2(new_n500), .A3(new_n674), .A4(new_n670), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT108), .ZN(new_n680));
  INV_X1    g494(.A(new_n602), .ZN(new_n681));
  OR3_X1    g495(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n680), .B1(new_n679), .B2(new_n681), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(new_n250), .ZN(G36));
  NOR2_X1   g499(.A1(new_n285), .A2(new_n286), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n290), .A2(KEYINPUT45), .A3(new_n292), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT45), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n265), .B1(new_n277), .B2(new_n261), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n688), .B1(new_n689), .B2(new_n291), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n687), .A2(new_n690), .A3(G469), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(KEYINPUT109), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT109), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n687), .A2(new_n690), .A3(new_n693), .A4(G469), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n686), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n287), .B1(new_n695), .B2(KEYINPUT46), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT46), .ZN(new_n697));
  AOI211_X1 g511(.A(new_n697), .B(new_n686), .C1(new_n692), .C2(new_n694), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n298), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  OR2_X1    g513(.A1(new_n699), .A2(new_n624), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n559), .A2(new_n596), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n351), .A2(new_n352), .ZN(new_n703));
  XOR2_X1   g517(.A(KEYINPUT110), .B(KEYINPUT43), .Z(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n703), .A2(new_n339), .A3(new_n570), .A4(new_n705), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n339), .A2(new_n351), .A3(new_n570), .A4(new_n352), .ZN(new_n707));
  NAND2_X1  g521(.A1(KEYINPUT110), .A2(KEYINPUT43), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  AND2_X1   g524(.A1(new_n702), .A2(new_n710), .ZN(new_n711));
  OR2_X1    g525(.A1(new_n711), .A2(KEYINPUT44), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n702), .A2(KEYINPUT44), .A3(new_n710), .ZN(new_n713));
  OR2_X1    g527(.A1(new_n713), .A2(KEYINPUT111), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(KEYINPUT111), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n714), .A2(new_n670), .A3(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT112), .ZN(new_n717));
  AND2_X1   g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n716), .A2(new_n717), .ZN(new_n719));
  OAI211_X1 g533(.A(new_n701), .B(new_n712), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G137), .ZN(G39));
  INV_X1    g535(.A(KEYINPUT47), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n699), .A2(new_n722), .ZN(new_n723));
  OAI211_X1 g537(.A(KEYINPUT47), .B(new_n298), .C1(new_n696), .C2(new_n698), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(new_n672), .ZN(new_n726));
  OR3_X1    g540(.A1(new_n726), .A2(new_n500), .A3(new_n467), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G140), .ZN(G42));
  NAND2_X1  g542(.A1(new_n710), .A2(new_n598), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n647), .A2(new_n670), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n731), .A2(new_n590), .A3(new_n662), .ZN(new_n732));
  INV_X1    g546(.A(new_n298), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n645), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n723), .A2(new_n724), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n661), .A2(new_n464), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n500), .B(new_n736), .C1(new_n555), .C2(new_n557), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n729), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n735), .A2(new_n670), .A3(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT119), .ZN(new_n740));
  INV_X1    g554(.A(new_n737), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n741), .A2(new_n598), .A3(new_n647), .A4(new_n710), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n629), .A2(new_n632), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n740), .B(KEYINPUT50), .C1(new_n742), .C2(new_n744), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n729), .A2(new_n737), .A3(new_n646), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n740), .A2(KEYINPUT50), .ZN(new_n747));
  OR2_X1    g561(.A1(new_n740), .A2(KEYINPUT50), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n746), .A2(new_n747), .A3(new_n748), .A4(new_n743), .ZN(new_n749));
  AND3_X1   g563(.A1(new_n739), .A2(new_n745), .A3(new_n749), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n730), .A2(new_n504), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n622), .A2(new_n500), .A3(new_n577), .A4(new_n751), .ZN(new_n752));
  OAI211_X1 g566(.A(new_n732), .B(new_n750), .C1(new_n752), .C2(new_n570), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT51), .ZN(new_n754));
  AND3_X1   g568(.A1(new_n753), .A2(KEYINPUT118), .A3(new_n754), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n754), .B1(new_n753), .B2(KEYINPUT118), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n467), .A2(new_n500), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n731), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(KEYINPUT48), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n622), .A2(new_n500), .A3(new_n751), .ZN(new_n761));
  OAI211_X1 g575(.A(new_n760), .B(new_n502), .C1(new_n761), .C2(new_n571), .ZN(new_n762));
  NOR3_X1   g576(.A1(new_n755), .A2(new_n756), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n738), .A2(new_n666), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT53), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n671), .A2(new_n601), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n591), .A2(new_n467), .A3(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT115), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n591), .A2(new_n467), .A3(KEYINPUT115), .A4(new_n766), .ZN(new_n770));
  AOI22_X1  g584(.A1(new_n682), .A2(new_n683), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n662), .A2(new_n590), .ZN(new_n772));
  NOR4_X1   g586(.A1(new_n772), .A2(new_n673), .A3(new_n669), .A4(new_n671), .ZN(new_n773));
  INV_X1    g587(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n596), .A2(new_n600), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n663), .A2(new_n674), .ZN(new_n776));
  AOI211_X1 g590(.A(new_n775), .B(new_n776), .C1(new_n620), .C2(new_n616), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n603), .A2(new_n640), .A3(new_n667), .ZN(new_n778));
  OAI21_X1  g592(.A(KEYINPUT52), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  AND3_X1   g593(.A1(new_n603), .A2(new_n640), .A3(new_n667), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n781));
  INV_X1    g595(.A(new_n775), .ZN(new_n782));
  INV_X1    g596(.A(new_n776), .ZN(new_n783));
  OAI211_X1 g597(.A(new_n782), .B(new_n783), .C1(new_n615), .C2(new_n617), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n780), .A2(new_n781), .A3(new_n784), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n771), .A2(new_n774), .A3(new_n779), .A4(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n677), .ZN(new_n787));
  INV_X1    g601(.A(new_n571), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n551), .A2(KEYINPUT114), .A3(new_n788), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n546), .A2(new_n549), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n546), .A2(new_n549), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n508), .B(new_n788), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT114), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n789), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n552), .B1(new_n795), .B2(new_n560), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n559), .A2(new_n500), .A3(new_n551), .A4(new_n302), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n592), .B1(new_n797), .B2(new_n578), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n648), .A2(new_n652), .A3(new_n656), .A4(new_n664), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n787), .A2(new_n799), .A3(new_n801), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n765), .B1(new_n786), .B2(new_n802), .ZN(new_n803));
  NOR4_X1   g617(.A1(new_n677), .A2(new_n796), .A3(new_n798), .A4(new_n800), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n779), .A2(new_n785), .ZN(new_n805));
  AOI221_X4 g619(.A(new_n773), .B1(new_n769), .B2(new_n770), .C1(new_n682), .C2(new_n683), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n804), .A2(new_n805), .A3(new_n806), .A4(KEYINPUT53), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n803), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(KEYINPUT54), .ZN(new_n809));
  XNOR2_X1  g623(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  XOR2_X1   g625(.A(new_n800), .B(KEYINPUT116), .Z(new_n812));
  NAND4_X1  g626(.A1(new_n812), .A2(KEYINPUT53), .A3(new_n787), .A4(new_n799), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n803), .B(new_n811), .C1(new_n786), .C2(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n763), .A2(new_n764), .A3(new_n809), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n501), .A2(new_n263), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT113), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(KEYINPUT49), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n818), .A2(KEYINPUT49), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n500), .B(new_n819), .C1(new_n645), .C2(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n821), .A2(new_n629), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n645), .A2(new_n820), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n707), .A2(new_n511), .A3(new_n733), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n622), .A2(new_n822), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n817), .A2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT120), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n817), .A2(KEYINPUT120), .A3(new_n825), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(G75));
  OR2_X1    g644(.A1(new_n813), .A2(new_n786), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n286), .B1(new_n831), .B2(new_n803), .ZN(new_n832));
  AOI21_X1  g646(.A(KEYINPUT56), .B1(new_n832), .B2(G210), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n530), .B1(new_n533), .B2(new_n534), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(new_n515), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n835), .B(KEYINPUT55), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n836), .B1(KEYINPUT121), .B2(KEYINPUT56), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n833), .A2(new_n838), .ZN(new_n839));
  AOI211_X1 g653(.A(KEYINPUT56), .B(new_n837), .C1(new_n832), .C2(G210), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n263), .A2(G952), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(G51));
  NOR2_X1   g656(.A1(new_n813), .A2(new_n786), .ZN(new_n843));
  INV_X1    g657(.A(new_n803), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n810), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n845), .A2(KEYINPUT122), .A3(new_n814), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT122), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n847), .B(new_n810), .C1(new_n843), .C2(new_n844), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n686), .B(KEYINPUT57), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n846), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(new_n284), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n832), .A2(new_n694), .A3(new_n692), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n841), .B1(new_n851), .B2(new_n852), .ZN(G54));
  NAND3_X1  g667(.A1(new_n832), .A2(KEYINPUT58), .A3(G475), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n346), .A2(new_n347), .ZN(new_n855));
  INV_X1    g669(.A(new_n855), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n854), .A2(new_n856), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n857), .A2(new_n858), .A3(new_n841), .ZN(G60));
  NAND2_X1  g673(.A1(new_n563), .A2(new_n565), .ZN(new_n860));
  XOR2_X1   g674(.A(new_n567), .B(KEYINPUT59), .Z(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  AND4_X1   g676(.A1(new_n860), .A2(new_n846), .A3(new_n848), .A4(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n841), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n861), .B1(new_n809), .B2(new_n814), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n864), .B1(new_n865), .B2(new_n860), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n863), .A2(new_n866), .ZN(G63));
  NOR2_X1   g681(.A1(new_n587), .A2(new_n588), .ZN(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(G217), .A2(G902), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(KEYINPUT125), .ZN(new_n871));
  XNOR2_X1  g685(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n872));
  XOR2_X1   g686(.A(new_n871), .B(new_n872), .Z(new_n873));
  OAI211_X1 g687(.A(new_n869), .B(new_n873), .C1(new_n843), .C2(new_n844), .ZN(new_n874));
  INV_X1    g688(.A(new_n873), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n875), .B1(new_n831), .B2(new_n803), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n495), .B(KEYINPUT126), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n874), .B(new_n864), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT123), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n878), .A2(new_n879), .A3(KEYINPUT61), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT61), .B1(new_n878), .B2(new_n879), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n880), .A2(new_n881), .ZN(G66));
  AOI21_X1  g696(.A(new_n263), .B1(new_n506), .B2(G224), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n799), .A2(new_n801), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n883), .B1(new_n884), .B2(new_n263), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n834), .B1(G898), .B2(new_n263), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n885), .B(new_n886), .Z(G69));
  INV_X1    g701(.A(KEYINPUT62), .ZN(new_n888));
  INV_X1    g702(.A(new_n636), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n888), .B1(new_n889), .B2(new_n778), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n636), .A2(KEYINPUT62), .A3(new_n780), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AOI211_X1 g706(.A(new_n626), .B(new_n757), .C1(new_n571), .C2(new_n578), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(new_n670), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n720), .A2(new_n892), .A3(new_n727), .A4(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(new_n263), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n433), .A2(new_n434), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(new_n342), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n898), .B(KEYINPUT127), .Z(new_n899));
  NAND2_X1  g713(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(G900), .A2(G953), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n701), .A2(new_n758), .A3(new_n663), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n684), .A2(new_n778), .A3(new_n902), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n720), .A2(new_n787), .A3(new_n727), .A4(new_n903), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n901), .B(new_n898), .C1(new_n904), .C2(G953), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n900), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n263), .B1(G227), .B2(G900), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(new_n907), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n900), .A2(new_n909), .A3(new_n905), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n908), .A2(new_n910), .ZN(G72));
  NAND2_X1  g725(.A1(G472), .A2(G902), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(KEYINPUT63), .Z(new_n913));
  OAI21_X1  g727(.A(new_n913), .B1(new_n895), .B2(new_n884), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n914), .A2(new_n386), .A3(new_n436), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n913), .B1(new_n904), .B2(new_n884), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(new_n437), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n436), .A2(new_n387), .ZN(new_n918));
  AOI22_X1  g732(.A1(new_n803), .A2(new_n807), .B1(new_n447), .B2(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n841), .B1(new_n919), .B2(new_n913), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n915), .A2(new_n917), .A3(new_n920), .ZN(G57));
endmodule


