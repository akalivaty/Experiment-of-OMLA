//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 0 0 0 0 1 0 0 1 0 0 1 1 1 0 1 1 0 1 1 0 0 0 1 1 1 1 1 1 0 0 1 0 0 0 0 0 1 0 0 0 0 0 1 1 0 0 1 1 0 0 1 0 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:32 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(new_n201), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G1), .A2(G13), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n207), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(G1), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n209), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(G13), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n216), .B(G250), .C1(G257), .C2(G264), .ZN(new_n217));
  INV_X1    g0017(.A(KEYINPUT0), .ZN(new_n218));
  AOI21_X1  g0018(.A(new_n212), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G87), .ZN(new_n221));
  INV_X1    g0021(.A(G250), .ZN(new_n222));
  INV_X1    g0022(.A(G97), .ZN(new_n223));
  INV_X1    g0023(.A(G257), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n215), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n219), .B1(new_n218), .B2(new_n217), .C1(new_n229), .C2(KEYINPUT1), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XOR2_X1   g0035(.A(G250), .B(G257), .Z(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G68), .B(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT64), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G50), .ZN(new_n242));
  INV_X1    g0042(.A(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n244), .B(new_n248), .ZN(G351));
  NAND2_X1  g0049(.A1(new_n213), .A2(G13), .ZN(new_n250));
  NOR3_X1   g0050(.A1(new_n250), .A2(new_n209), .A3(G68), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(KEYINPUT12), .ZN(new_n252));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n208), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n254), .B1(new_n213), .B2(G20), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n252), .B1(G68), .B2(new_n255), .ZN(new_n256));
  NOR2_X1   g0056(.A1(G20), .A2(G33), .ZN(new_n257));
  INV_X1    g0057(.A(G68), .ZN(new_n258));
  AOI22_X1  g0058(.A1(new_n257), .A2(G50), .B1(G20), .B2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  OAI21_X1  g0060(.A(KEYINPUT66), .B1(new_n260), .B2(G20), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT66), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n262), .A2(new_n209), .A3(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G77), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n259), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(new_n254), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT11), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n266), .A2(KEYINPUT11), .A3(new_n254), .ZN(new_n270));
  AND3_X1   g0070(.A1(new_n256), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G41), .ZN(new_n273));
  INV_X1    g0073(.A(G45), .ZN(new_n274));
  AOI21_X1  g0074(.A(G1), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(KEYINPUT65), .B1(new_n275), .B2(G274), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n213), .B(G274), .C1(G41), .C2(G45), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT65), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n208), .B1(G33), .B2(G41), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n281), .A2(new_n275), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n280), .B1(G238), .B2(new_n282), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT3), .B(G33), .ZN(new_n284));
  INV_X1    g0084(.A(G1698), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n284), .A2(G226), .A3(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n284), .A2(G232), .A3(G1698), .ZN(new_n287));
  NAND2_X1  g0087(.A1(G33), .A2(G97), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  AND3_X1   g0089(.A1(new_n289), .A2(KEYINPUT70), .A3(new_n281), .ZN(new_n290));
  AOI21_X1  g0090(.A(KEYINPUT70), .B1(new_n289), .B2(new_n281), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n283), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT71), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n292), .A2(new_n293), .A3(KEYINPUT13), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT13), .ZN(new_n295));
  OAI221_X1 g0095(.A(new_n283), .B1(KEYINPUT71), .B2(new_n295), .C1(new_n290), .C2(new_n291), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n294), .A2(new_n296), .A3(G179), .ZN(new_n297));
  XNOR2_X1  g0097(.A(new_n297), .B(KEYINPUT74), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n292), .A2(new_n295), .ZN(new_n299));
  OAI211_X1 g0099(.A(KEYINPUT13), .B(new_n283), .C1(new_n290), .C2(new_n291), .ZN(new_n300));
  INV_X1    g0100(.A(G169), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT73), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n301), .B1(new_n302), .B2(KEYINPUT14), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n299), .A2(new_n300), .A3(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n302), .A2(KEYINPUT14), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n304), .B(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n272), .B1(new_n298), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n294), .A2(new_n296), .A3(G190), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n299), .A2(G200), .A3(new_n300), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n310), .A2(new_n311), .A3(new_n271), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT72), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n310), .A2(new_n311), .A3(KEYINPUT72), .A4(new_n271), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT3), .ZN(new_n318));
  OAI21_X1  g0118(.A(KEYINPUT75), .B1(new_n318), .B2(G33), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT75), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n320), .A2(new_n260), .A3(KEYINPUT3), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n318), .A2(G33), .ZN(new_n322));
  AND3_X1   g0122(.A1(new_n319), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(KEYINPUT7), .B1(new_n323), .B2(G20), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n319), .A2(new_n321), .A3(new_n322), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT7), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n325), .A2(new_n326), .A3(new_n209), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n324), .A2(G68), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(G58), .A2(G68), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  OAI21_X1  g0130(.A(G20), .B1(new_n330), .B2(new_n201), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT76), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  OAI211_X1 g0133(.A(KEYINPUT76), .B(G20), .C1(new_n330), .C2(new_n201), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n257), .A2(G159), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n328), .A2(KEYINPUT16), .A3(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT16), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n326), .B1(new_n284), .B2(G20), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(new_n322), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n342), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n258), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n339), .B1(new_n344), .B2(new_n336), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n338), .A2(new_n345), .A3(new_n254), .ZN(new_n346));
  NAND2_X1  g0146(.A1(G226), .A2(G1698), .ZN(new_n347));
  INV_X1    g0147(.A(G223), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n347), .B1(new_n348), .B2(G1698), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n349), .A2(new_n319), .A3(new_n321), .A4(new_n322), .ZN(new_n350));
  NAND2_X1  g0150(.A1(G33), .A2(G87), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n281), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n275), .A2(KEYINPUT65), .A3(G274), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n277), .A2(new_n278), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n282), .A2(G232), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(G200), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(new_n357), .B2(G190), .ZN(new_n360));
  INV_X1    g0160(.A(G13), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n361), .A2(G1), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(G20), .ZN(new_n363));
  XNOR2_X1  g0163(.A(KEYINPUT8), .B(G58), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n365), .B1(new_n255), .B2(new_n364), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n346), .A2(new_n360), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(KEYINPUT78), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT78), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n346), .A2(new_n360), .A3(new_n369), .A4(new_n366), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n368), .A2(KEYINPUT17), .A3(new_n370), .ZN(new_n371));
  OR2_X1    g0171(.A1(new_n367), .A2(KEYINPUT17), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n346), .A2(new_n366), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT77), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n301), .B1(new_n353), .B2(new_n356), .ZN(new_n376));
  OAI211_X1 g0176(.A(G1), .B(G13), .C1(new_n260), .C2(new_n273), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n377), .B1(new_n350), .B2(new_n351), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n213), .B1(G41), .B2(G45), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n377), .A2(G232), .A3(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(new_n276), .B2(new_n279), .ZN(new_n381));
  INV_X1    g0181(.A(G179), .ZN(new_n382));
  NOR3_X1   g0182(.A1(new_n378), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n375), .B1(new_n376), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(G169), .B1(new_n378), .B2(new_n381), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n385), .B(KEYINPUT77), .C1(new_n357), .C2(new_n382), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n374), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(KEYINPUT18), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n346), .A2(new_n366), .B1(new_n384), .B2(new_n386), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT18), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AND2_X1   g0192(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n373), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n363), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n395), .A2(G77), .ZN(new_n396));
  INV_X1    g0196(.A(new_n255), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n396), .B1(new_n397), .B2(G77), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n257), .ZN(new_n400));
  OAI22_X1  g0200(.A1(new_n364), .A2(new_n400), .B1(new_n209), .B2(new_n265), .ZN(new_n401));
  XOR2_X1   g0201(.A(KEYINPUT15), .B(G87), .Z(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(KEYINPUT67), .ZN(new_n403));
  XNOR2_X1  g0203(.A(KEYINPUT15), .B(G87), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT67), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AND2_X1   g0206(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n264), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n401), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n254), .ZN(new_n410));
  OAI211_X1 g0210(.A(KEYINPUT68), .B(new_n399), .C1(new_n409), .C2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT68), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n409), .A2(new_n410), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n412), .B1(new_n413), .B2(new_n398), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n284), .A2(G232), .A3(new_n285), .ZN(new_n415));
  INV_X1    g0215(.A(G107), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n284), .A2(G1698), .ZN(new_n417));
  INV_X1    g0217(.A(G238), .ZN(new_n418));
  OAI221_X1 g0218(.A(new_n415), .B1(new_n416), .B2(new_n284), .C1(new_n417), .C2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n281), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n280), .B1(G244), .B2(new_n282), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(G190), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n422), .A2(new_n358), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n411), .A2(new_n414), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n413), .A2(new_n398), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n423), .A2(G179), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n422), .A2(G169), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n428), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n427), .A2(new_n431), .ZN(new_n432));
  MUX2_X1   g0232(.A(new_n395), .B(new_n255), .S(G50), .Z(new_n433));
  INV_X1    g0233(.A(new_n364), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n408), .A2(new_n434), .ZN(new_n435));
  AOI22_X1  g0235(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n257), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n410), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n433), .A2(new_n437), .ZN(new_n438));
  XOR2_X1   g0238(.A(new_n438), .B(KEYINPUT9), .Z(new_n439));
  NAND3_X1  g0239(.A1(new_n284), .A2(G222), .A3(new_n285), .ZN(new_n440));
  OAI221_X1 g0240(.A(new_n440), .B1(new_n265), .B2(new_n284), .C1(new_n417), .C2(new_n348), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n281), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n280), .B1(G226), .B2(new_n282), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n358), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n445), .B1(G190), .B2(new_n444), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n439), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(KEYINPUT10), .B1(new_n446), .B2(KEYINPUT69), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n439), .B(new_n446), .C1(KEYINPUT69), .C2(KEYINPUT10), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n444), .A2(G169), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n451), .B1(new_n382), .B2(new_n444), .ZN(new_n452));
  INV_X1    g0252(.A(new_n438), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n432), .A2(new_n449), .A3(new_n450), .A4(new_n454), .ZN(new_n455));
  NOR4_X1   g0255(.A1(new_n309), .A2(new_n317), .A3(new_n394), .A4(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n363), .A2(G116), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n410), .B(new_n363), .C1(G1), .C2(new_n260), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n457), .B1(new_n459), .B2(G116), .ZN(new_n460));
  INV_X1    g0260(.A(G116), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(G20), .ZN(new_n462));
  AOI21_X1  g0262(.A(KEYINPUT86), .B1(new_n254), .B2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n254), .A2(KEYINPUT86), .A3(new_n462), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(G33), .A2(G283), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n467), .B(new_n209), .C1(G33), .C2(new_n223), .ZN(new_n468));
  AOI21_X1  g0268(.A(KEYINPUT20), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  AND3_X1   g0269(.A1(new_n254), .A2(KEYINPUT86), .A3(new_n462), .ZN(new_n470));
  OAI211_X1 g0270(.A(KEYINPUT20), .B(new_n468), .C1(new_n470), .C2(new_n463), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n460), .B1(new_n469), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n213), .A2(G45), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT5), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n475), .A2(G41), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n474), .B1(new_n476), .B2(KEYINPUT81), .ZN(new_n477));
  OAI21_X1  g0277(.A(KEYINPUT81), .B1(new_n273), .B2(KEYINPUT5), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n273), .A2(KEYINPUT5), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n477), .A2(G274), .A3(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n281), .B1(new_n477), .B2(new_n480), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n482), .B1(G270), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(G264), .A2(G1698), .ZN(new_n485));
  INV_X1    g0285(.A(G303), .ZN(new_n486));
  OAI22_X1  g0286(.A1(new_n325), .A2(new_n485), .B1(new_n486), .B2(new_n284), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n323), .A2(KEYINPUT85), .A3(G257), .A4(new_n285), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT85), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n319), .A2(new_n321), .A3(new_n285), .A4(new_n322), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n489), .B1(new_n490), .B2(new_n224), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n487), .B1(new_n488), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n484), .B1(new_n492), .B2(new_n377), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n473), .A2(new_n493), .A3(G169), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT21), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n473), .A2(new_n493), .A3(KEYINPUT21), .A4(G169), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n484), .B(G179), .C1(new_n492), .C2(new_n377), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(new_n473), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n496), .A2(new_n497), .A3(new_n500), .ZN(new_n501));
  OR2_X1    g0301(.A1(new_n493), .A2(G190), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n493), .A2(new_n358), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n473), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT6), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n223), .A2(new_n416), .ZN(new_n507));
  NOR2_X1   g0307(.A1(G97), .A2(G107), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n416), .A2(KEYINPUT6), .A3(G97), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n511), .A2(G20), .B1(G77), .B2(new_n257), .ZN(new_n512));
  NOR3_X1   g0312(.A1(new_n284), .A2(new_n326), .A3(G20), .ZN(new_n513));
  AOI21_X1  g0313(.A(KEYINPUT7), .B1(new_n342), .B2(new_n209), .ZN(new_n514));
  OAI21_X1  g0314(.A(G107), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n410), .B1(new_n512), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n395), .A2(KEYINPUT79), .A3(new_n223), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT79), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(new_n363), .B2(G97), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n517), .B(new_n519), .C1(new_n458), .C2(new_n223), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT4), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n319), .A2(new_n321), .A3(G244), .A4(new_n322), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n522), .B1(new_n523), .B2(G1698), .ZN(new_n524));
  AND2_X1   g0324(.A1(KEYINPUT4), .A2(G244), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n341), .A2(new_n322), .A3(new_n525), .A4(new_n285), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT80), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n341), .A2(new_n322), .A3(G250), .A4(G1698), .ZN(new_n529));
  AND2_X1   g0329(.A1(new_n529), .A2(new_n467), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n284), .A2(KEYINPUT80), .A3(new_n285), .A4(new_n525), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n524), .A2(new_n528), .A3(new_n530), .A4(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n281), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n477), .A2(new_n480), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n534), .A2(G257), .A3(new_n377), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n481), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n533), .A2(new_n537), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n538), .A2(G190), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n536), .B1(new_n532), .B2(new_n281), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n540), .A2(G200), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n521), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n467), .B(new_n529), .C1(new_n526), .C2(new_n527), .ZN(new_n543));
  AND2_X1   g0343(.A1(new_n526), .A2(new_n527), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n377), .B1(new_n545), .B2(new_n524), .ZN(new_n546));
  OAI21_X1  g0346(.A(G169), .B1(new_n546), .B2(new_n536), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n533), .A2(new_n537), .A3(G179), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OR2_X1    g0349(.A1(new_n516), .A2(new_n520), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n363), .B1(new_n403), .B2(new_n406), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n323), .A2(KEYINPUT84), .A3(new_n209), .A4(G68), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT84), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n319), .A2(new_n321), .A3(new_n209), .A4(new_n322), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n554), .B1(new_n555), .B2(new_n258), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n261), .A2(new_n263), .A3(G97), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT19), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n209), .B1(new_n288), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(G87), .A2(G97), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n416), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n557), .A2(new_n558), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n553), .A2(new_n556), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n552), .B1(new_n563), .B2(new_n254), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n407), .A2(new_n459), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n323), .A2(KEYINPUT83), .A3(G238), .A4(new_n285), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT83), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(new_n490), .B2(new_n418), .ZN(new_n569));
  NAND2_X1  g0369(.A1(G33), .A2(G116), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n571), .B1(KEYINPUT75), .B2(new_n341), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n572), .A2(G244), .A3(G1698), .A4(new_n321), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n567), .A2(new_n569), .A3(new_n570), .A4(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n281), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT82), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n474), .A2(new_n576), .A3(G250), .ZN(new_n577));
  AOI21_X1  g0377(.A(G274), .B1(KEYINPUT82), .B2(G250), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n577), .B1(new_n474), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n377), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n575), .A2(new_n382), .A3(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n580), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n582), .B1(new_n574), .B2(new_n281), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n566), .B(new_n581), .C1(G169), .C2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n575), .A2(G190), .A3(new_n580), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n458), .A2(new_n221), .ZN(new_n586));
  AOI211_X1 g0386(.A(new_n552), .B(new_n586), .C1(new_n563), .C2(new_n254), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n585), .B(new_n587), .C1(new_n358), .C2(new_n583), .ZN(new_n588));
  AND4_X1   g0388(.A1(new_n542), .A2(new_n551), .A3(new_n584), .A4(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n362), .A2(G20), .A3(new_n416), .ZN(new_n590));
  XNOR2_X1  g0390(.A(new_n590), .B(KEYINPUT25), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n591), .B1(G107), .B2(new_n459), .ZN(new_n592));
  INV_X1    g0392(.A(G264), .ZN(new_n593));
  AOI211_X1 g0393(.A(new_n593), .B(new_n281), .C1(new_n477), .C2(new_n480), .ZN(new_n594));
  NAND2_X1  g0394(.A1(G257), .A2(G1698), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(new_n222), .B2(G1698), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n596), .A2(new_n319), .A3(new_n321), .A4(new_n322), .ZN(new_n597));
  NAND2_X1  g0397(.A1(G33), .A2(G294), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n377), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NOR3_X1   g0399(.A1(new_n594), .A2(new_n482), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n424), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n601), .B1(new_n600), .B2(G200), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT87), .ZN(new_n603));
  NAND2_X1  g0403(.A1(KEYINPUT22), .A2(G87), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n555), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n221), .A2(G20), .ZN(new_n606));
  AOI21_X1  g0406(.A(KEYINPUT22), .B1(new_n284), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n603), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT22), .ZN(new_n609));
  INV_X1    g0409(.A(new_n606), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n609), .B1(new_n342), .B2(new_n610), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n611), .B(KEYINPUT87), .C1(new_n555), .C2(new_n604), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n570), .A2(G20), .ZN(new_n614));
  AOI21_X1  g0414(.A(KEYINPUT23), .B1(new_n416), .B2(G20), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n416), .A2(KEYINPUT23), .A3(G20), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n614), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n613), .A2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT24), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n254), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n618), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n622), .B1(new_n608), .B2(new_n612), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n623), .A2(KEYINPUT24), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n592), .B(new_n602), .C1(new_n621), .C2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n594), .A2(new_n599), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n301), .B1(new_n627), .B2(new_n481), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n628), .B1(G179), .B2(new_n600), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n619), .A2(new_n620), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n410), .B1(new_n623), .B2(KEYINPUT24), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n629), .B1(new_n632), .B2(new_n592), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n626), .A2(new_n633), .ZN(new_n634));
  AND4_X1   g0434(.A1(new_n456), .A2(new_n505), .A3(new_n589), .A4(new_n634), .ZN(G372));
  INV_X1    g0435(.A(KEYINPUT74), .ZN(new_n636));
  XNOR2_X1  g0436(.A(new_n297), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g0437(.A(new_n304), .B(new_n305), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n639), .A2(new_n272), .B1(new_n312), .B2(new_n431), .ZN(new_n640));
  INV_X1    g0440(.A(new_n373), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n393), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n449), .A2(new_n450), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n642), .A2(new_n643), .B1(new_n453), .B2(new_n452), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n625), .A2(new_n542), .A3(new_n551), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n382), .A2(new_n583), .B1(new_n564), .B2(new_n565), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT88), .ZN(new_n647));
  XNOR2_X1  g0447(.A(new_n580), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n575), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n301), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n649), .A2(G200), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n652), .A2(new_n585), .A3(new_n587), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n645), .A2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n592), .B1(new_n621), .B2(new_n624), .ZN(new_n656));
  INV_X1    g0456(.A(new_n629), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n500), .A2(new_n497), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(new_n496), .A3(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(KEYINPUT89), .B1(new_n655), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n538), .A2(new_n358), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n540), .A2(new_n424), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n550), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n521), .B1(new_n547), .B2(new_n548), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n585), .A2(new_n587), .ZN(new_n667));
  AOI22_X1  g0467(.A1(new_n667), .A2(new_n652), .B1(new_n646), .B2(new_n650), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n666), .A2(new_n668), .A3(new_n625), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n501), .A2(new_n633), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT89), .ZN(new_n671));
  NOR3_X1   g0471(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT90), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n584), .A2(new_n588), .A3(new_n665), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(KEYINPUT26), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT26), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n651), .A2(new_n653), .A3(new_n676), .A4(new_n665), .ZN(new_n677));
  AND4_X1   g0477(.A1(new_n673), .A2(new_n675), .A3(new_n651), .A4(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n651), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n679), .B1(new_n674), .B2(KEYINPUT26), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n673), .B1(new_n680), .B2(new_n677), .ZN(new_n681));
  OAI22_X1  g0481(.A1(new_n661), .A2(new_n672), .B1(new_n678), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n456), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n644), .A2(new_n683), .ZN(G369));
  INV_X1    g0484(.A(KEYINPUT27), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n685), .B1(new_n362), .B2(new_n209), .ZN(new_n686));
  NOR3_X1   g0486(.A1(new_n250), .A2(KEYINPUT27), .A3(G20), .ZN(new_n687));
  INV_X1    g0487(.A(G213), .ZN(new_n688));
  NOR3_X1   g0488(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(G343), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n473), .A2(new_n691), .ZN(new_n692));
  MUX2_X1   g0492(.A(new_n501), .B(new_n505), .S(new_n692), .Z(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(G330), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n658), .A2(new_n691), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n656), .A2(new_n691), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(new_n625), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n695), .B1(new_n658), .B2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n694), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n697), .A2(new_n658), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n691), .B1(new_n659), .B2(new_n496), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n695), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n701), .A2(new_n704), .ZN(G399));
  INV_X1    g0505(.A(new_n216), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(G41), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n560), .A2(new_n416), .A3(new_n461), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n708), .A2(G1), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(new_n207), .B2(new_n708), .ZN(new_n712));
  XNOR2_X1  g0512(.A(new_n712), .B(KEYINPUT28), .ZN(new_n713));
  OAI21_X1  g0513(.A(KEYINPUT26), .B1(new_n654), .B2(new_n551), .ZN(new_n714));
  OAI211_X1 g0514(.A(new_n714), .B(new_n651), .C1(KEYINPUT26), .C2(new_n674), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n669), .A2(new_n670), .ZN(new_n716));
  OAI211_X1 g0516(.A(KEYINPUT29), .B(new_n690), .C1(new_n715), .C2(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n675), .A2(new_n651), .A3(new_n677), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(KEYINPUT90), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n680), .A2(new_n673), .A3(new_n677), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n671), .B1(new_n669), .B2(new_n670), .ZN(new_n722));
  AND3_X1   g0522(.A1(new_n625), .A2(new_n542), .A3(new_n551), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n660), .A2(new_n723), .A3(KEYINPUT89), .A4(new_n668), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n691), .B1(new_n721), .B2(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n717), .B1(new_n726), .B2(KEYINPUT29), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT92), .ZN(new_n728));
  INV_X1    g0528(.A(G330), .ZN(new_n729));
  NAND2_X1  g0529(.A1(KEYINPUT91), .A2(KEYINPUT30), .ZN(new_n730));
  NOR2_X1   g0530(.A1(KEYINPUT91), .A2(KEYINPUT30), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n583), .A2(new_n540), .A3(new_n627), .A4(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n730), .B1(new_n733), .B2(new_n498), .ZN(new_n734));
  AND4_X1   g0534(.A1(new_n533), .A2(new_n537), .A3(new_n627), .A4(new_n732), .ZN(new_n735));
  INV_X1    g0535(.A(new_n730), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n735), .A2(new_n499), .A3(new_n583), .A4(new_n736), .ZN(new_n737));
  NOR3_X1   g0537(.A1(new_n540), .A2(G179), .A3(new_n600), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n738), .A2(new_n493), .A3(new_n649), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n734), .A2(new_n737), .A3(new_n739), .ZN(new_n740));
  AND3_X1   g0540(.A1(new_n740), .A2(KEYINPUT31), .A3(new_n691), .ZN(new_n741));
  AOI21_X1  g0541(.A(KEYINPUT31), .B1(new_n740), .B2(new_n691), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n634), .A2(new_n589), .A3(new_n505), .A4(new_n690), .ZN(new_n744));
  AOI211_X1 g0544(.A(new_n728), .B(new_n729), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n742), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n740), .A2(KEYINPUT31), .A3(new_n691), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n744), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(KEYINPUT92), .B1(new_n748), .B2(G330), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  AND2_X1   g0550(.A1(new_n727), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n713), .B1(new_n751), .B2(G1), .ZN(G364));
  NOR2_X1   g0552(.A1(G13), .A2(G33), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(G20), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n693), .A2(new_n756), .ZN(new_n757));
  OR2_X1    g0557(.A1(new_n301), .A2(KEYINPUT93), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n301), .A2(KEYINPUT93), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n209), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(new_n208), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n755), .ZN(new_n762));
  XNOR2_X1  g0562(.A(new_n762), .B(KEYINPUT94), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n706), .A2(new_n323), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n244), .A2(G45), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n207), .A2(new_n274), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n216), .A2(new_n284), .ZN(new_n769));
  INV_X1    g0569(.A(G355), .ZN(new_n770));
  OAI22_X1  g0570(.A1(new_n769), .A2(new_n770), .B1(G116), .B2(new_n216), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n763), .B1(new_n768), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n361), .A2(G20), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G45), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n708), .A2(G1), .A3(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n761), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n382), .A2(new_n358), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n209), .A2(new_n424), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(G326), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n342), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n382), .A2(G200), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n779), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n209), .A2(G190), .ZN(new_n786));
  NOR2_X1   g0586(.A1(G179), .A2(G200), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI22_X1  g0589(.A1(G322), .A2(new_n785), .B1(new_n789), .B2(G329), .ZN(new_n790));
  INV_X1    g0590(.A(G311), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n786), .A2(new_n783), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n778), .A2(new_n786), .ZN(new_n793));
  XOR2_X1   g0593(.A(KEYINPUT33), .B(G317), .Z(new_n794));
  OAI221_X1 g0594(.A(new_n790), .B1(new_n791), .B2(new_n792), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n787), .A2(G190), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(G20), .ZN(new_n797));
  AOI211_X1 g0597(.A(new_n782), .B(new_n795), .C1(G294), .C2(new_n797), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n779), .A2(new_n382), .A3(G200), .ZN(new_n799));
  OR2_X1    g0599(.A1(new_n799), .A2(KEYINPUT95), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(KEYINPUT95), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n786), .A2(new_n382), .A3(G200), .ZN(new_n804));
  XOR2_X1   g0604(.A(new_n804), .B(KEYINPUT96), .Z(new_n805));
  AOI22_X1  g0605(.A1(new_n803), .A2(G303), .B1(new_n805), .B2(G283), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n784), .A2(new_n243), .B1(new_n792), .B2(new_n265), .ZN(new_n807));
  INV_X1    g0607(.A(new_n797), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n284), .B1(new_n780), .B2(new_n202), .C1(new_n808), .C2(new_n223), .ZN(new_n809));
  INV_X1    g0609(.A(new_n793), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n807), .B(new_n809), .C1(G68), .C2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n803), .A2(G87), .ZN(new_n812));
  INV_X1    g0612(.A(G159), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n788), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT32), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n805), .A2(G107), .ZN(new_n816));
  AND3_X1   g0616(.A1(new_n812), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n798), .A2(new_n806), .B1(new_n811), .B2(new_n817), .ZN(new_n818));
  OAI211_X1 g0618(.A(new_n772), .B(new_n776), .C1(new_n777), .C2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n757), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT97), .ZN(new_n821));
  INV_X1    g0621(.A(new_n694), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n822), .A2(new_n776), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(G330), .B2(new_n693), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n821), .A2(new_n824), .ZN(G396));
  NOR2_X1   g0625(.A1(new_n761), .A2(new_n753), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n776), .B1(G77), .B2(new_n827), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT98), .ZN(new_n829));
  INV_X1    g0629(.A(G132), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n323), .B1(new_n830), .B2(new_n788), .ZN(new_n831));
  INV_X1    g0631(.A(new_n805), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n832), .A2(new_n258), .B1(new_n202), .B2(new_n802), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n831), .B(new_n833), .C1(G58), .C2(new_n797), .ZN(new_n834));
  INV_X1    g0634(.A(new_n780), .ZN(new_n835));
  INV_X1    g0635(.A(new_n792), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n835), .A2(G137), .B1(new_n836), .B2(G159), .ZN(new_n837));
  INV_X1    g0637(.A(G143), .ZN(new_n838));
  INV_X1    g0638(.A(G150), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n837), .B1(new_n838), .B2(new_n784), .C1(new_n839), .C2(new_n793), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n840), .B(KEYINPUT34), .ZN(new_n841));
  INV_X1    g0641(.A(G294), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n342), .B1(new_n788), .B2(new_n791), .C1(new_n842), .C2(new_n784), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n805), .A2(G87), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n844), .B1(new_n416), .B2(new_n802), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n843), .B(new_n845), .C1(G97), .C2(new_n797), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n780), .A2(new_n486), .B1(new_n792), .B2(new_n461), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n847), .B1(G283), .B2(new_n810), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT99), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n834), .A2(new_n841), .B1(new_n846), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n431), .A2(new_n691), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n428), .A2(new_n690), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(KEYINPUT100), .B1(new_n432), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT100), .ZN(new_n855));
  NOR4_X1   g0655(.A1(new_n427), .A2(new_n431), .A3(new_n855), .A4(new_n852), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n851), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n829), .B1(new_n777), .B2(new_n850), .C1(new_n857), .C2(new_n754), .ZN(new_n858));
  OR2_X1    g0658(.A1(new_n726), .A2(new_n857), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n682), .A2(new_n690), .A3(new_n857), .ZN(new_n860));
  AND2_X1   g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n748), .A2(G330), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n728), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n748), .A2(KEYINPUT92), .A3(G330), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n776), .B1(new_n861), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n861), .A2(new_n865), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n858), .B1(new_n867), .B2(new_n868), .ZN(G384));
  NAND2_X1  g0669(.A1(new_n329), .A2(G77), .ZN(new_n870));
  OAI22_X1  g0670(.A1(new_n207), .A2(new_n870), .B1(G50), .B2(new_n258), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n871), .A2(G1), .A3(new_n361), .ZN(new_n872));
  INV_X1    g0672(.A(new_n511), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT35), .ZN(new_n874));
  AOI211_X1 g0674(.A(new_n461), .B(new_n211), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n875), .B1(new_n874), .B2(new_n873), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT36), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n872), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n878), .B1(new_n877), .B2(new_n876), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT38), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT102), .ZN(new_n881));
  INV_X1    g0681(.A(new_n367), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n881), .B1(new_n882), .B2(new_n390), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n689), .B(KEYINPUT101), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n884), .B1(new_n346), .B2(new_n366), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n388), .A2(KEYINPUT102), .A3(new_n367), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n883), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  AND2_X1   g0688(.A1(new_n368), .A2(new_n370), .ZN(new_n889));
  NOR3_X1   g0689(.A1(new_n390), .A2(new_n885), .A3(KEYINPUT37), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n888), .A2(KEYINPUT37), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n886), .B1(new_n373), .B2(new_n393), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n880), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT39), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n338), .A2(new_n254), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT16), .B1(new_n328), .B2(new_n337), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n366), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n897), .B1(new_n387), .B2(new_n689), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n898), .A2(new_n368), .A3(new_n370), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(KEYINPUT37), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n890), .A2(new_n368), .A3(new_n370), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n389), .A2(new_n392), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n903), .B1(new_n372), .B2(new_n371), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n897), .A2(new_n689), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n902), .B(KEYINPUT38), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n893), .A2(new_n894), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n905), .B1(new_n373), .B2(new_n393), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n889), .A2(new_n890), .B1(new_n899), .B2(KEYINPUT37), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n880), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n910), .A2(new_n906), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n907), .B1(new_n911), .B2(new_n894), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n308), .A2(new_n691), .ZN(new_n913));
  AOI22_X1  g0713(.A1(new_n912), .A2(new_n913), .B1(new_n903), .B2(new_n884), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n316), .A2(new_n637), .A3(new_n638), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n272), .A2(new_n691), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n312), .A2(new_n916), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n915), .A2(new_n917), .B1(new_n308), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n431), .A2(new_n690), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n920), .B1(new_n860), .B2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n911), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n914), .A2(new_n924), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n456), .B(new_n717), .C1(new_n726), .C2(KEYINPUT29), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n644), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n925), .B(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT40), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n298), .A2(new_n307), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n916), .B1(new_n930), .B2(new_n316), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n918), .B1(new_n639), .B2(new_n272), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n748), .B(new_n857), .C1(new_n931), .C2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n929), .B1(new_n911), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n893), .A2(new_n906), .ZN(new_n935));
  INV_X1    g0735(.A(new_n920), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n748), .A2(new_n857), .ZN(new_n937));
  NAND4_X1  g0737(.A1(new_n935), .A2(new_n936), .A3(new_n937), .A4(KEYINPUT40), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n934), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n456), .A2(new_n748), .ZN(new_n940));
  XOR2_X1   g0740(.A(new_n939), .B(new_n940), .Z(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(G330), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n928), .A2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT103), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OAI221_X1 g0745(.A(new_n945), .B1(new_n213), .B2(new_n773), .C1(new_n928), .C2(new_n942), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n943), .A2(new_n944), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n879), .B1(new_n946), .B2(new_n947), .ZN(G367));
  OAI21_X1  g0748(.A(new_n666), .B1(new_n521), .B2(new_n690), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n551), .B2(new_n690), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n698), .A2(new_n703), .A3(new_n950), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n951), .A2(KEYINPUT42), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(KEYINPUT42), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n551), .B1(new_n949), .B2(new_n658), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n690), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n952), .A2(new_n953), .A3(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n587), .A2(new_n690), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n668), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n958), .B1(new_n651), .B2(new_n957), .ZN(new_n959));
  XOR2_X1   g0759(.A(KEYINPUT104), .B(KEYINPUT43), .Z(new_n960));
  NOR2_X1   g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n956), .A2(new_n962), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n963), .A2(KEYINPUT105), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n961), .B1(KEYINPUT43), .B2(new_n959), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n963), .A2(KEYINPUT105), .B1(new_n956), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n700), .A2(new_n950), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT106), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n967), .B(new_n969), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n707), .B(KEYINPUT41), .Z(new_n971));
  NAND2_X1  g0771(.A1(new_n704), .A2(new_n950), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n972), .A2(KEYINPUT107), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(KEYINPUT107), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT45), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n973), .A2(KEYINPUT45), .A3(new_n974), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n704), .A2(new_n950), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT44), .ZN(new_n980));
  AND3_X1   g0780(.A1(new_n977), .A2(new_n978), .A3(new_n980), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n698), .B(new_n703), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(new_n822), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n751), .A2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT109), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n981), .A2(new_n701), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n977), .A2(new_n978), .A3(new_n980), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n700), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(KEYINPUT108), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT108), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n987), .A2(new_n990), .A3(new_n700), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n751), .A2(KEYINPUT109), .A3(new_n983), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n986), .A2(new_n989), .A3(new_n991), .A4(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n971), .B1(new_n993), .B2(new_n751), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n774), .A2(G1), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n970), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n765), .A2(new_n238), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n407), .A2(new_n706), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n762), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n325), .B1(new_n784), .B2(new_n486), .C1(new_n791), .C2(new_n780), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n804), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n1001), .A2(G97), .B1(new_n789), .B2(G317), .ZN(new_n1002));
  INV_X1    g0802(.A(G283), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n1002), .B1(new_n1003), .B2(new_n792), .C1(new_n842), .C2(new_n793), .ZN(new_n1004));
  AOI211_X1 g0804(.A(new_n1000), .B(new_n1004), .C1(G107), .C2(new_n797), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT46), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n802), .B2(new_n461), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n803), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1005), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n1009), .B(KEYINPUT110), .Z(new_n1010));
  OAI22_X1  g0810(.A1(new_n838), .A2(new_n780), .B1(new_n804), .B2(new_n265), .ZN(new_n1011));
  AOI211_X1 g0811(.A(new_n342), .B(new_n1011), .C1(G137), .C2(new_n789), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n803), .A2(G58), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n797), .A2(G68), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n784), .A2(new_n839), .B1(new_n792), .B2(new_n202), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(G159), .B2(new_n810), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .A4(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1010), .A2(KEYINPUT47), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(new_n761), .ZN(new_n1019));
  AOI21_X1  g0819(.A(KEYINPUT47), .B1(new_n1010), .B2(new_n1017), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n776), .B1(new_n997), .B2(new_n999), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1021), .B(KEYINPUT111), .Z(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n756), .B2(new_n959), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n996), .A2(new_n1023), .ZN(G387));
  NAND2_X1  g0824(.A1(new_n699), .A2(new_n755), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n803), .A2(G294), .B1(G283), .B2(new_n797), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT48), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n835), .A2(G322), .B1(new_n836), .B2(G303), .ZN(new_n1028));
  INV_X1    g0828(.A(G317), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1028), .B1(new_n791), .B2(new_n793), .C1(new_n1029), .C2(new_n784), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1026), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(KEYINPUT112), .B(KEYINPUT49), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n1001), .A2(G116), .B1(new_n789), .B2(G326), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1034), .A2(new_n325), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n780), .A2(new_n813), .B1(new_n793), .B2(new_n364), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n323), .B1(new_n258), .B2(new_n792), .C1(new_n839), .C2(new_n788), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n1038), .B(new_n1039), .C1(G50), .C2(new_n785), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n805), .A2(G97), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n407), .A2(new_n797), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n803), .A2(G77), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n777), .B1(new_n1037), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n434), .A2(new_n202), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT50), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n710), .B(new_n274), .C1(new_n258), .C2(new_n265), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n764), .B1(new_n1047), .B2(new_n1048), .C1(new_n235), .C2(new_n274), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1049), .B1(G107), .B2(new_n216), .C1(new_n710), .C2(new_n769), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n775), .B(new_n1045), .C1(new_n763), .C2(new_n1050), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n983), .A2(new_n995), .B1(new_n1025), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n984), .A2(new_n707), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n751), .A2(new_n983), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1052), .B1(new_n1053), .B2(new_n1054), .ZN(G393));
  NAND2_X1  g0855(.A1(new_n981), .A2(new_n701), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1056), .A2(new_n988), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n708), .B1(new_n1057), .B2(new_n984), .ZN(new_n1058));
  AND2_X1   g0858(.A1(new_n1058), .A2(new_n993), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n762), .B1(new_n223), .B2(new_n216), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n765), .A2(new_n248), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n776), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT52), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n780), .A2(new_n1029), .B1(new_n784), .B2(new_n791), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n805), .A2(G107), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1065), .B1(new_n1063), .B2(new_n1064), .C1(new_n1003), .C2(new_n802), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(G303), .A2(new_n810), .B1(new_n789), .B2(G322), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n284), .B1(new_n836), .B2(G294), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1067), .B(new_n1068), .C1(new_n461), .C2(new_n808), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n780), .A2(new_n839), .B1(new_n784), .B2(new_n813), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT51), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1071), .B(new_n844), .C1(new_n258), .C2(new_n802), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n810), .A2(G50), .B1(new_n836), .B2(new_n434), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n325), .B1(G77), .B2(new_n797), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1073), .B(new_n1074), .C1(new_n838), .C2(new_n788), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n1066), .A2(new_n1069), .B1(new_n1072), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1062), .B1(new_n1076), .B2(new_n761), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(new_n950), .B2(new_n756), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n995), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1078), .B1(new_n1057), .B2(new_n1079), .ZN(new_n1080));
  OR2_X1    g0880(.A1(new_n1059), .A2(new_n1080), .ZN(G390));
  NAND3_X1  g0881(.A1(new_n748), .A2(G330), .A3(new_n857), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1082), .A2(new_n920), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n894), .B1(new_n910), .B2(new_n906), .ZN(new_n1085));
  AND2_X1   g0885(.A1(new_n893), .A2(new_n906), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1085), .B1(new_n1086), .B2(new_n894), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n922), .B2(new_n913), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1086), .A2(new_n913), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n854), .A2(new_n856), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1090), .B(new_n690), .C1(new_n715), .C2(new_n716), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(new_n921), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n936), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1089), .A2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1084), .B1(new_n1088), .B2(new_n1094), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n857), .B(new_n936), .C1(new_n745), .C2(new_n749), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1088), .A2(new_n1094), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT113), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n913), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n921), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(new_n726), .B2(new_n857), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1100), .B1(new_n1102), .B2(new_n920), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n1103), .A2(new_n1087), .B1(new_n1093), .B2(new_n1089), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1104), .A2(KEYINPUT113), .A3(new_n1096), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1095), .B1(new_n1099), .B2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n456), .A2(G330), .A3(new_n748), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n926), .A2(new_n644), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1102), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n936), .B1(new_n865), .B2(new_n857), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1109), .B1(new_n1110), .B2(new_n1083), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1092), .B1(new_n920), .B2(new_n1082), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n1096), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1108), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n707), .B1(new_n1106), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1095), .ZN(new_n1116));
  AOI21_X1  g0916(.A(KEYINPUT113), .B1(new_n1104), .B2(new_n1096), .ZN(new_n1117));
  AND4_X1   g0917(.A1(KEYINPUT113), .A2(new_n1088), .A3(new_n1094), .A4(new_n1096), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1116), .B(new_n1114), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  OR2_X1    g0920(.A1(new_n1115), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1087), .A2(new_n753), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n802), .A2(new_n839), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1123), .B(KEYINPUT53), .ZN(new_n1124));
  INV_X1    g0924(.A(G137), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(KEYINPUT54), .B(G143), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n793), .A2(new_n1125), .B1(new_n792), .B2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1127), .B1(G159), .B2(new_n797), .ZN(new_n1128));
  XOR2_X1   g0928(.A(new_n1128), .B(KEYINPUT114), .Z(new_n1129));
  AOI21_X1  g0929(.A(new_n342), .B1(new_n835), .B2(G128), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n202), .A2(new_n804), .B1(new_n784), .B2(new_n830), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(G125), .B2(new_n789), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1124), .A2(new_n1129), .A3(new_n1130), .A4(new_n1132), .ZN(new_n1133));
  OAI221_X1 g0933(.A(new_n342), .B1(new_n793), .B2(new_n416), .C1(new_n808), .C2(new_n265), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n784), .A2(new_n461), .B1(new_n788), .B2(new_n842), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n780), .A2(new_n1003), .B1(new_n792), .B2(new_n223), .ZN(new_n1136));
  NOR3_X1   g0936(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1137), .B(new_n812), .C1(new_n258), .C2(new_n832), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n777), .B1(new_n1133), .B2(new_n1138), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n775), .B(new_n1139), .C1(new_n364), .C2(new_n826), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n1106), .A2(new_n995), .B1(new_n1122), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1121), .A2(new_n1141), .ZN(G378));
  AOI21_X1  g0942(.A(new_n1108), .B1(new_n1106), .B2(new_n1114), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n934), .A2(new_n938), .A3(G330), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n914), .A2(new_n1144), .A3(new_n924), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1144), .B1(new_n914), .B2(new_n924), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT119), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n643), .A2(new_n454), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1148), .B(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n453), .A2(new_n689), .ZN(new_n1151));
  XOR2_X1   g0951(.A(new_n1151), .B(KEYINPUT55), .Z(new_n1152));
  XNOR2_X1  g0952(.A(new_n1150), .B(new_n1152), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n1145), .A2(new_n1146), .B1(new_n1147), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1144), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n925), .A2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1153), .A2(new_n1147), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n914), .A2(new_n1144), .A3(new_n924), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  AND2_X1   g0959(.A1(new_n1154), .A2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(KEYINPUT57), .B1(new_n1143), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1108), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1119), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT57), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1154), .A2(new_n1159), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n708), .B1(new_n1161), .B2(new_n1166), .ZN(new_n1167));
  OR2_X1    g0967(.A1(new_n1153), .A2(new_n754), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(G116), .A2(new_n835), .B1(new_n785), .B2(G107), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1169), .B(new_n1014), .C1(new_n223), .C2(new_n793), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1001), .A2(G58), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1043), .B(new_n1171), .C1(new_n1003), .C2(new_n788), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n325), .A2(new_n273), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  XOR2_X1   g0974(.A(new_n1174), .B(KEYINPUT115), .Z(new_n1175));
  AOI211_X1 g0975(.A(new_n1170), .B(new_n1175), .C1(new_n407), .C2(new_n836), .ZN(new_n1176));
  AOI21_X1  g0976(.A(G50), .B1(new_n260), .B2(new_n273), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n1176), .A2(KEYINPUT58), .B1(new_n1173), .B2(new_n1177), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n835), .A2(G125), .B1(new_n797), .B2(G150), .ZN(new_n1179));
  XOR2_X1   g0979(.A(new_n1179), .B(KEYINPUT116), .Z(new_n1180));
  AOI22_X1  g0980(.A1(G128), .A2(new_n785), .B1(new_n836), .B2(G137), .ZN(new_n1181));
  OAI221_X1 g0981(.A(new_n1181), .B1(new_n830), .B2(new_n793), .C1(new_n802), .C2(new_n1126), .ZN(new_n1182));
  OR2_X1    g0982(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  OR2_X1    g0983(.A1(new_n1183), .A2(KEYINPUT59), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(KEYINPUT59), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n260), .B(new_n273), .C1(new_n804), .C2(new_n813), .ZN(new_n1186));
  XOR2_X1   g0986(.A(KEYINPUT117), .B(G124), .Z(new_n1187));
  AOI21_X1  g0987(.A(new_n1186), .B1(new_n789), .B2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1184), .A2(new_n1185), .A3(new_n1188), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1178), .B(new_n1189), .C1(KEYINPUT58), .C2(new_n1176), .ZN(new_n1190));
  AND2_X1   g0990(.A1(new_n1190), .A2(new_n761), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n775), .B(new_n1191), .C1(new_n202), .C2(new_n826), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n1165), .A2(new_n995), .B1(new_n1168), .B2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  NOR3_X1   g0994(.A1(new_n1167), .A2(KEYINPUT120), .A3(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT120), .ZN(new_n1196));
  AOI221_X4 g0996(.A(KEYINPUT57), .B1(new_n1154), .B2(new_n1159), .C1(new_n1119), .C2(new_n1162), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1164), .B1(new_n1163), .B2(new_n1165), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n707), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1196), .B1(new_n1199), .B2(new_n1193), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1195), .A2(new_n1200), .ZN(G375));
  INV_X1    g1001(.A(new_n1114), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n857), .B1(new_n745), .B2(new_n749), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1083), .B1(new_n1203), .B2(new_n920), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1113), .B(new_n1108), .C1(new_n1204), .C2(new_n1102), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n971), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1202), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1079), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n920), .A2(new_n753), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n776), .B1(new_n827), .B2(G68), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1042), .B1(new_n223), .B2(new_n802), .C1(new_n832), .C2(new_n265), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(G116), .A2(new_n810), .B1(new_n785), .B2(G283), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(G107), .A2(new_n836), .B1(new_n789), .B2(G303), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n284), .B1(new_n835), .B2(G294), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n836), .A2(G150), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n797), .A2(G50), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1171), .A2(new_n1216), .A3(new_n1217), .A4(new_n323), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1126), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(G137), .A2(new_n785), .B1(new_n810), .B2(new_n1219), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n835), .A2(G132), .B1(new_n789), .B2(G128), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1220), .B(new_n1221), .C1(new_n802), .C2(new_n813), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n1211), .A2(new_n1215), .B1(new_n1218), .B2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1210), .B1(new_n1223), .B2(new_n761), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1208), .B1(new_n1209), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1207), .A2(new_n1225), .ZN(G381));
  INV_X1    g1026(.A(G378), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n1195), .B2(new_n1200), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1059), .A2(new_n1080), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1229), .A2(new_n996), .A3(new_n1023), .ZN(new_n1230));
  OR2_X1    g1030(.A1(G393), .A2(G396), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(G384), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  OR4_X1    g1034(.A1(G381), .A2(new_n1228), .A3(new_n1230), .A4(new_n1234), .ZN(G407));
  OAI211_X1 g1035(.A(G407), .B(G213), .C1(G343), .C2(new_n1228), .ZN(G409));
  NOR2_X1   g1036(.A1(new_n688), .A2(G343), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1193), .B(new_n1141), .C1(new_n1120), .C2(new_n1115), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1163), .A2(new_n1206), .A3(new_n1165), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1237), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(G378), .B1(new_n1167), .B2(new_n1194), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  OR2_X1    g1043(.A1(new_n1243), .A2(KEYINPUT123), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT125), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1205), .B(KEYINPUT60), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT121), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1114), .A2(new_n708), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1246), .A2(new_n1247), .A3(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(new_n1225), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1247), .B1(new_n1246), .B2(new_n1248), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1233), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT122), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1246), .A2(new_n1248), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(KEYINPUT121), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1255), .A2(G384), .A3(new_n1225), .A4(new_n1249), .ZN(new_n1256));
  AND3_X1   g1056(.A1(new_n1252), .A2(new_n1253), .A3(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1253), .B1(new_n1252), .B2(new_n1256), .ZN(new_n1258));
  XOR2_X1   g1058(.A(KEYINPUT124), .B(G2897), .Z(new_n1259));
  NOR3_X1   g1059(.A1(new_n1259), .A2(new_n688), .A3(G343), .ZN(new_n1260));
  NOR3_X1   g1060(.A1(new_n1257), .A2(new_n1258), .A3(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1252), .A2(new_n1256), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1262), .A2(G2897), .A3(new_n1237), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1245), .B1(new_n1261), .B2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1262), .A2(KEYINPUT122), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1252), .A2(new_n1253), .A3(new_n1256), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  OAI211_X1 g1068(.A(KEYINPUT125), .B(new_n1263), .C1(new_n1268), .C2(new_n1260), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1243), .A2(KEYINPUT123), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1244), .A2(new_n1265), .A3(new_n1269), .A4(new_n1270), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1241), .A2(new_n1242), .A3(new_n1266), .A4(new_n1267), .ZN(new_n1272));
  XNOR2_X1  g1072(.A(new_n1272), .B(KEYINPUT63), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT61), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(G387), .A2(G390), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(new_n1230), .ZN(new_n1276));
  XNOR2_X1  g1076(.A(G393), .B(G396), .ZN(new_n1277));
  OR2_X1    g1077(.A1(new_n1277), .A2(KEYINPUT126), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(KEYINPUT126), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1276), .A2(new_n1278), .A3(new_n1279), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1275), .A2(new_n1277), .A3(KEYINPUT126), .A4(new_n1230), .ZN(new_n1281));
  AND2_X1   g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1271), .A2(new_n1273), .A3(new_n1274), .A4(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1265), .A2(new_n1269), .A3(new_n1243), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1272), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT62), .ZN(new_n1286));
  AOI21_X1  g1086(.A(KEYINPUT61), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1272), .A2(KEYINPUT62), .ZN(new_n1288));
  AND3_X1   g1088(.A1(new_n1284), .A2(new_n1287), .A3(new_n1288), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1283), .B1(new_n1289), .B2(new_n1282), .ZN(G405));
  NAND3_X1  g1090(.A1(new_n1228), .A2(new_n1242), .A3(new_n1268), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1262), .ZN(new_n1292));
  OAI21_X1  g1092(.A(KEYINPUT120), .B1(new_n1167), .B2(new_n1194), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1199), .A2(new_n1196), .A3(new_n1193), .ZN(new_n1294));
  AOI21_X1  g1094(.A(G378), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1242), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1292), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1291), .A2(new_n1297), .A3(new_n1282), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1282), .B1(new_n1291), .B2(new_n1297), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1298), .B1(new_n1299), .B2(KEYINPUT127), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT127), .ZN(new_n1301));
  AOI211_X1 g1101(.A(new_n1301), .B(new_n1282), .C1(new_n1297), .C2(new_n1291), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1300), .A2(new_n1302), .ZN(G402));
endmodule


