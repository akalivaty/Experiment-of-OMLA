//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 1 1 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 0 1 0 0 0 0 1 0 0 0 0 0 1 0 1 1 1 1 0 0 0 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:38 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n555, new_n556, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n618, new_n619, new_n622, new_n624, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1173, new_n1174, new_n1175, new_n1176;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT66), .Z(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n452), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n452), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  OR2_X1    g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(G2105), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  AOI22_X1  g041(.A1(new_n464), .A2(G137), .B1(G101), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G125), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n468), .B1(new_n462), .B2(new_n463), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(KEYINPUT67), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT67), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n472), .A2(G113), .A3(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g049(.A(G2105), .B1(new_n469), .B2(new_n474), .ZN(new_n475));
  AND2_X1   g050(.A1(new_n467), .A2(new_n475), .ZN(G160));
  NAND2_X1  g051(.A1(new_n464), .A2(G136), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n465), .B1(new_n462), .B2(new_n463), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n477), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  AND2_X1   g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  NOR2_X1   g059(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n485));
  OAI211_X1 g060(.A(G126), .B(G2105), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  OR2_X1    g061(.A1(G102), .A2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G114), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n487), .A2(new_n489), .A3(G2104), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n493), .B1(new_n484), .B2(new_n485), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n493), .B(new_n496), .C1(new_n485), .C2(new_n484), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n491), .B1(new_n495), .B2(new_n497), .ZN(G164));
  INV_X1    g073(.A(G543), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n499), .A2(KEYINPUT5), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT69), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n501), .B1(new_n502), .B2(G543), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n499), .A2(KEYINPUT69), .A3(KEYINPUT5), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n500), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n506), .A2(KEYINPUT6), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT68), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n508), .B1(new_n509), .B2(G651), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n506), .A2(KEYINPUT68), .A3(KEYINPUT6), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n507), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n505), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G50), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n513), .A2(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n505), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n518), .A2(new_n506), .ZN(new_n519));
  OR2_X1    g094(.A1(new_n517), .A2(new_n519), .ZN(G303));
  INV_X1    g095(.A(G303), .ZN(G166));
  AND2_X1   g096(.A1(G63), .A2(G651), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n523), .A2(KEYINPUT7), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(KEYINPUT7), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n505), .A2(new_n522), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n505), .A2(new_n512), .A3(G89), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n512), .A2(G51), .A3(G543), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT70), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g106(.A1(new_n526), .A2(new_n527), .A3(KEYINPUT70), .A4(new_n528), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(G168));
  INV_X1    g108(.A(G90), .ZN(new_n534));
  INV_X1    g109(.A(G52), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n513), .A2(new_n534), .B1(new_n515), .B2(new_n535), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n505), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n506), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n536), .A2(new_n538), .ZN(G171));
  NAND2_X1  g114(.A1(G68), .A2(G543), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n502), .A2(G543), .ZN(new_n541));
  AND3_X1   g116(.A1(new_n499), .A2(KEYINPUT69), .A3(KEYINPUT5), .ZN(new_n542));
  AOI21_X1  g117(.A(KEYINPUT69), .B1(new_n499), .B2(KEYINPUT5), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(G56), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n540), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT71), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n506), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n548), .B1(new_n547), .B2(new_n546), .ZN(new_n549));
  INV_X1    g124(.A(new_n513), .ZN(new_n550));
  INV_X1    g125(.A(new_n515), .ZN(new_n551));
  AOI22_X1  g126(.A1(G81), .A2(new_n550), .B1(new_n551), .B2(G43), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n549), .A2(G860), .A3(new_n552), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  OAI211_X1 g132(.A(G65), .B(new_n541), .C1(new_n542), .C2(new_n543), .ZN(new_n558));
  AND2_X1   g133(.A1(G78), .A2(G543), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT72), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n506), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  AND3_X1   g136(.A1(new_n505), .A2(new_n512), .A3(G91), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n510), .A2(new_n511), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n509), .A2(G651), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n564), .A2(G53), .A3(G543), .A4(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(KEYINPUT9), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT9), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n512), .A2(new_n568), .A3(G53), .A4(G543), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n563), .A2(new_n570), .ZN(G299));
  INV_X1    g146(.A(G171), .ZN(G301));
  INV_X1    g147(.A(G168), .ZN(G286));
  NAND2_X1  g148(.A1(new_n550), .A2(G87), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n551), .A2(G49), .ZN(new_n575));
  OAI21_X1  g150(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(G288));
  NAND2_X1  g152(.A1(new_n505), .A2(G61), .ZN(new_n578));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(G651), .ZN(new_n581));
  AND2_X1   g156(.A1(G48), .A2(G543), .ZN(new_n582));
  AND3_X1   g157(.A1(new_n506), .A2(KEYINPUT68), .A3(KEYINPUT6), .ZN(new_n583));
  AOI21_X1  g158(.A(KEYINPUT68), .B1(new_n506), .B2(KEYINPUT6), .ZN(new_n584));
  OAI211_X1 g159(.A(new_n565), .B(new_n582), .C1(new_n583), .C2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT73), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n512), .A2(KEYINPUT73), .A3(new_n582), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n505), .A2(new_n512), .A3(G86), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n581), .A2(new_n589), .A3(new_n590), .ZN(G305));
  NAND2_X1  g166(.A1(G72), .A2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G60), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n544), .B2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT74), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n506), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n596), .B1(new_n595), .B2(new_n594), .ZN(new_n597));
  AOI22_X1  g172(.A1(G85), .A2(new_n550), .B1(new_n551), .B2(G47), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(G290));
  NAND2_X1  g174(.A1(G301), .A2(G868), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT75), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n550), .A2(new_n601), .A3(G92), .ZN(new_n602));
  INV_X1    g177(.A(G92), .ZN(new_n603));
  OAI21_X1  g178(.A(KEYINPUT75), .B1(new_n513), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n602), .A2(KEYINPUT10), .A3(new_n604), .ZN(new_n608));
  NAND2_X1  g183(.A1(G79), .A2(G543), .ZN(new_n609));
  INV_X1    g184(.A(G66), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n544), .B2(new_n610), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n611), .A2(G651), .B1(new_n551), .B2(G54), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n607), .A2(new_n608), .A3(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n600), .B1(new_n614), .B2(G868), .ZN(G284));
  OAI21_X1  g190(.A(new_n600), .B1(new_n614), .B2(G868), .ZN(G321));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  NOR2_X1   g192(.A1(G286), .A2(new_n617), .ZN(new_n618));
  XOR2_X1   g193(.A(G299), .B(KEYINPUT76), .Z(new_n619));
  AOI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(new_n617), .ZN(G297));
  AOI21_X1  g195(.A(new_n618), .B1(new_n619), .B2(new_n617), .ZN(G280));
  INV_X1    g196(.A(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n614), .B1(new_n622), .B2(G860), .ZN(G148));
  NAND2_X1  g198(.A1(new_n549), .A2(new_n552), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(new_n617), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n613), .A2(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(new_n617), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g203(.A(KEYINPUT3), .B(G2104), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(new_n466), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(KEYINPUT12), .Z(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT13), .Z(new_n632));
  XOR2_X1   g207(.A(KEYINPUT77), .B(G2100), .Z(new_n633));
  OR2_X1    g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n464), .A2(G135), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n478), .A2(G123), .ZN(new_n637));
  OR2_X1    g212(.A1(G99), .A2(G2105), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n638), .B(G2104), .C1(G111), .C2(new_n465), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n636), .A2(new_n637), .A3(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(G2096), .Z(new_n641));
  NAND3_X1  g216(.A1(new_n634), .A2(new_n635), .A3(new_n641), .ZN(G156));
  XNOR2_X1  g217(.A(G2427), .B(G2438), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2430), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2435), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n646), .A2(new_n647), .A3(KEYINPUT14), .ZN(new_n648));
  XOR2_X1   g223(.A(G1341), .B(G1348), .Z(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n648), .B(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2451), .B(G2454), .Z(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n652), .A2(new_n655), .ZN(new_n657));
  AND3_X1   g232(.A1(new_n656), .A2(G14), .A3(new_n657), .ZN(G401));
  INV_X1    g233(.A(KEYINPUT18), .ZN(new_n659));
  XOR2_X1   g234(.A(G2084), .B(G2090), .Z(new_n660));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n662), .A2(KEYINPUT17), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n660), .A2(new_n661), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n659), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G2100), .ZN(new_n666));
  XOR2_X1   g241(.A(G2072), .B(G2078), .Z(new_n667));
  AOI21_X1  g242(.A(new_n667), .B1(new_n662), .B2(KEYINPUT18), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G2096), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n666), .B(new_n669), .ZN(G227));
  XNOR2_X1  g245(.A(G1956), .B(G2474), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT79), .ZN(new_n672));
  XOR2_X1   g247(.A(G1961), .B(G1966), .Z(new_n673));
  OR2_X1    g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1971), .B(G1976), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT19), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n672), .A2(new_n673), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n674), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n677), .A2(new_n676), .ZN(new_n679));
  INV_X1    g254(.A(KEYINPUT20), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NOR3_X1   g256(.A1(new_n677), .A2(KEYINPUT20), .A3(new_n676), .ZN(new_n682));
  OAI221_X1 g257(.A(new_n678), .B1(new_n676), .B2(new_n674), .C1(new_n681), .C2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT80), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n685));
  AND2_X1   g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n684), .A2(new_n685), .ZN(new_n687));
  XOR2_X1   g262(.A(G1991), .B(G1996), .Z(new_n688));
  OR3_X1    g263(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1981), .B(G1986), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n688), .B1(new_n686), .B2(new_n687), .ZN(new_n691));
  AND3_X1   g266(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n690), .B1(new_n689), .B2(new_n691), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n692), .A2(new_n693), .ZN(G229));
  XOR2_X1   g269(.A(KEYINPUT95), .B(KEYINPUT23), .Z(new_n695));
  INV_X1    g270(.A(G16), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G20), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n695), .B(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(G299), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n698), .B1(new_n699), .B2(new_n696), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT96), .B(G1956), .Z(new_n701));
  XOR2_X1   g276(.A(new_n700), .B(new_n701), .Z(new_n702));
  AND2_X1   g277(.A1(new_n696), .A2(G19), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(new_n624), .B2(G16), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  AND2_X1   g280(.A1(new_n705), .A2(G1341), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n705), .A2(G1341), .ZN(new_n707));
  NOR3_X1   g282(.A1(new_n702), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n696), .A2(G4), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(new_n614), .B2(new_n696), .ZN(new_n710));
  INV_X1    g285(.A(G1348), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  AND3_X1   g287(.A1(G168), .A2(KEYINPUT90), .A3(G16), .ZN(new_n713));
  AOI21_X1  g288(.A(KEYINPUT90), .B1(G168), .B2(G16), .ZN(new_n714));
  OAI22_X1  g289(.A1(new_n713), .A2(new_n714), .B1(G16), .B2(G21), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(G1966), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n708), .A2(new_n712), .A3(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G29), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G26), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT28), .ZN(new_n720));
  AOI22_X1  g295(.A1(G128), .A2(new_n478), .B1(new_n464), .B2(G140), .ZN(new_n721));
  INV_X1    g296(.A(G104), .ZN(new_n722));
  AND3_X1   g297(.A1(new_n722), .A2(new_n465), .A3(KEYINPUT84), .ZN(new_n723));
  AOI21_X1  g298(.A(KEYINPUT84), .B1(new_n722), .B2(new_n465), .ZN(new_n724));
  OAI221_X1 g299(.A(G2104), .B1(G116), .B2(new_n465), .C1(new_n723), .C2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n721), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n720), .B1(new_n727), .B2(new_n718), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(G2067), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n718), .A2(G27), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G164), .B2(new_n718), .ZN(new_n731));
  INV_X1    g306(.A(G2078), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n718), .A2(G32), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n478), .A2(G129), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT88), .ZN(new_n736));
  NAND3_X1  g311(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT26), .Z(new_n738));
  NAND2_X1  g313(.A1(new_n464), .A2(G141), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n466), .A2(G105), .ZN(new_n740));
  AND3_X1   g315(.A1(new_n738), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n736), .A2(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n734), .B1(new_n742), .B2(new_n718), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT27), .B(G1996), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT89), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n733), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n718), .A2(G35), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G162), .B2(new_n718), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT29), .Z(new_n749));
  INV_X1    g324(.A(G2090), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AOI211_X1 g326(.A(new_n729), .B(new_n746), .C1(new_n751), .C2(KEYINPUT94), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(KEYINPUT94), .B2(new_n751), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n743), .A2(new_n745), .ZN(new_n754));
  NAND2_X1  g329(.A1(G160), .A2(G29), .ZN(new_n755));
  INV_X1    g330(.A(G34), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n756), .A2(KEYINPUT24), .ZN(new_n757));
  AOI21_X1  g332(.A(G29), .B1(new_n756), .B2(KEYINPUT24), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n757), .B1(new_n758), .B2(KEYINPUT87), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(KEYINPUT87), .B2(new_n758), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n755), .A2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(G2084), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n696), .A2(G5), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G171), .B2(new_n696), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n754), .B(new_n763), .C1(G1961), .C2(new_n765), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT93), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n765), .A2(G1961), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT92), .Z(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT31), .B(G11), .ZN(new_n770));
  XOR2_X1   g345(.A(KEYINPUT30), .B(G28), .Z(new_n771));
  OAI21_X1  g346(.A(new_n770), .B1(new_n771), .B2(G29), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n640), .A2(new_n718), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n772), .B1(new_n773), .B2(KEYINPUT91), .ZN(new_n774));
  OAI221_X1 g349(.A(new_n774), .B1(KEYINPUT91), .B2(new_n773), .C1(new_n761), .C2(new_n762), .ZN(new_n775));
  INV_X1    g350(.A(G2072), .ZN(new_n776));
  AND2_X1   g351(.A1(new_n718), .A2(G33), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT85), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT25), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n464), .A2(G139), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT86), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n629), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n780), .B(new_n782), .C1(new_n465), .C2(new_n783), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n777), .B1(new_n784), .B2(G29), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n775), .B1(new_n776), .B2(new_n785), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n749), .A2(new_n750), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n785), .A2(new_n776), .ZN(new_n788));
  NAND4_X1  g363(.A1(new_n769), .A2(new_n786), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  NOR4_X1   g364(.A1(new_n717), .A2(new_n753), .A3(new_n767), .A4(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  MUX2_X1   g366(.A(G6), .B(G305), .S(G16), .Z(new_n792));
  XOR2_X1   g367(.A(KEYINPUT32), .B(G1981), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n696), .A2(G22), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G166), .B2(new_n696), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n796), .A2(G1971), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n796), .A2(G1971), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n696), .A2(G23), .ZN(new_n799));
  AND3_X1   g374(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(new_n696), .ZN(new_n801));
  XNOR2_X1  g376(.A(KEYINPUT33), .B(G1976), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n794), .A2(new_n797), .A3(new_n798), .A4(new_n803), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT83), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT34), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n805), .A2(new_n806), .ZN(new_n808));
  MUX2_X1   g383(.A(G24), .B(G290), .S(G16), .Z(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(G1986), .Z(new_n810));
  NAND2_X1  g385(.A1(new_n718), .A2(G25), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT81), .ZN(new_n812));
  NOR2_X1   g387(.A1(G95), .A2(G2105), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT82), .Z(new_n814));
  OAI21_X1  g389(.A(G2104), .B1(new_n465), .B2(G107), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n464), .A2(G131), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n478), .A2(G119), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n812), .B1(new_n821), .B2(new_n718), .ZN(new_n822));
  XOR2_X1   g397(.A(KEYINPUT35), .B(G1991), .Z(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n807), .A2(new_n808), .A3(new_n810), .A4(new_n824), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n825), .A2(KEYINPUT36), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(KEYINPUT36), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n791), .B1(new_n826), .B2(new_n827), .ZN(G311));
  NAND2_X1  g403(.A1(new_n826), .A2(new_n827), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(new_n790), .ZN(G150));
  NAND2_X1  g405(.A1(new_n614), .A2(G559), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT38), .ZN(new_n832));
  INV_X1    g407(.A(G93), .ZN(new_n833));
  INV_X1    g408(.A(G55), .ZN(new_n834));
  OAI22_X1  g409(.A1(new_n513), .A2(new_n833), .B1(new_n515), .B2(new_n834), .ZN(new_n835));
  AOI22_X1  g410(.A1(new_n505), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n836), .A2(new_n506), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n624), .B(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n832), .B(new_n839), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n840), .A2(KEYINPUT39), .ZN(new_n841));
  INV_X1    g416(.A(G860), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n840), .A2(KEYINPUT39), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n838), .A2(new_n842), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT37), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n844), .A2(new_n846), .ZN(G145));
  XNOR2_X1  g422(.A(KEYINPUT100), .B(G37), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n742), .B(new_n727), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n495), .A2(new_n497), .ZN(new_n851));
  INV_X1    g426(.A(new_n491), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n742), .B(new_n726), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(G164), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n784), .A2(KEYINPUT98), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n854), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n784), .A2(KEYINPUT98), .ZN(new_n859));
  OR2_X1    g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n858), .A2(new_n859), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n820), .B(KEYINPUT99), .ZN(new_n863));
  INV_X1    g438(.A(new_n631), .ZN(new_n864));
  AND2_X1   g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n863), .A2(new_n864), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n464), .A2(G142), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n478), .A2(G130), .ZN(new_n868));
  OR2_X1    g443(.A1(G106), .A2(G2105), .ZN(new_n869));
  OAI211_X1 g444(.A(new_n869), .B(G2104), .C1(G118), .C2(new_n465), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n867), .A2(new_n868), .A3(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  OR3_X1    g447(.A1(new_n865), .A2(new_n866), .A3(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n872), .B1(new_n865), .B2(new_n866), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n862), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g451(.A1(new_n860), .A2(new_n874), .A3(new_n873), .A4(new_n861), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  XOR2_X1   g453(.A(G160), .B(KEYINPUT97), .Z(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(new_n482), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(new_n640), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n878), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n876), .A2(new_n881), .A3(new_n877), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n849), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n885), .B(KEYINPUT40), .Z(G395));
  INV_X1    g461(.A(new_n838), .ZN(new_n887));
  AOI21_X1  g462(.A(KEYINPUT101), .B1(new_n887), .B2(new_n617), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n839), .B1(G559), .B2(new_n613), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n624), .B(new_n887), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(new_n626), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n614), .A2(new_n699), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n613), .A2(G299), .ZN(new_n894));
  AOI21_X1  g469(.A(KEYINPUT41), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AND3_X1   g470(.A1(new_n893), .A2(KEYINPUT41), .A3(new_n894), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n892), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n893), .A2(new_n894), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n889), .A2(new_n898), .A3(new_n891), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  OR2_X1    g475(.A1(new_n900), .A2(KEYINPUT42), .ZN(new_n901));
  XNOR2_X1  g476(.A(G290), .B(G305), .ZN(new_n902));
  XNOR2_X1  g477(.A(G303), .B(new_n800), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n902), .B(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n900), .A2(KEYINPUT42), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n901), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(G868), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n905), .B1(new_n901), .B2(new_n906), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n888), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n909), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n911), .A2(KEYINPUT101), .A3(G868), .A4(new_n907), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n910), .A2(new_n912), .ZN(G295));
  AND2_X1   g488(.A1(new_n910), .A2(new_n912), .ZN(G331));
  XNOR2_X1  g489(.A(G168), .B(G171), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n839), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n890), .A2(new_n915), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n919), .B1(new_n896), .B2(new_n895), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n917), .A2(new_n918), .A3(new_n898), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(new_n904), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n920), .A2(new_n905), .A3(new_n921), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n849), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT43), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(G37), .B1(new_n923), .B2(new_n924), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n927), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n925), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT103), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n932), .A2(new_n933), .A3(KEYINPUT43), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT103), .B1(new_n925), .B2(new_n926), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n934), .A2(KEYINPUT44), .A3(new_n935), .ZN(new_n936));
  AND3_X1   g511(.A1(new_n928), .A2(KEYINPUT102), .A3(new_n926), .ZN(new_n937));
  AOI21_X1  g512(.A(KEYINPUT102), .B1(new_n928), .B2(new_n926), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n931), .B1(new_n936), .B2(new_n939), .ZN(G397));
  INV_X1    g515(.A(KEYINPUT45), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n941), .B1(G164), .B2(G1384), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n467), .A2(new_n475), .A3(G40), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n944), .B(KEYINPUT104), .ZN(new_n945));
  INV_X1    g520(.A(new_n742), .ZN(new_n946));
  INV_X1    g521(.A(G2067), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n726), .B(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n945), .B1(new_n946), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(G1996), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n944), .A2(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n952), .B(KEYINPUT46), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n950), .A2(new_n953), .ZN(new_n954));
  XOR2_X1   g529(.A(new_n954), .B(KEYINPUT47), .Z(new_n955));
  NOR2_X1   g530(.A1(G290), .A2(G1986), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(new_n944), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n957), .B(KEYINPUT126), .ZN(new_n958));
  XOR2_X1   g533(.A(KEYINPUT125), .B(KEYINPUT48), .Z(new_n959));
  OR2_X1    g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n948), .B1(new_n951), .B2(new_n742), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n945), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n962), .B1(new_n946), .B2(new_n952), .ZN(new_n963));
  XOR2_X1   g538(.A(new_n820), .B(new_n823), .Z(new_n964));
  AOI21_X1  g539(.A(new_n963), .B1(new_n964), .B2(new_n945), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n958), .A2(new_n959), .ZN(new_n966));
  AND3_X1   g541(.A1(new_n960), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n821), .A2(new_n823), .ZN(new_n968));
  OAI22_X1  g543(.A1(new_n963), .A2(new_n968), .B1(G2067), .B2(new_n726), .ZN(new_n969));
  AOI211_X1 g544(.A(new_n955), .B(new_n967), .C1(new_n945), .C2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT124), .ZN(new_n971));
  AND2_X1   g546(.A1(G290), .A2(G1986), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n944), .B1(new_n972), .B2(new_n956), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n965), .A2(new_n973), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n467), .A2(new_n475), .A3(G40), .ZN(new_n975));
  AOI21_X1  g550(.A(G1384), .B1(new_n851), .B2(new_n852), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(G1976), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n977), .B(G8), .C1(G288), .C2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(KEYINPUT52), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT52), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n981), .B1(new_n800), .B2(G1976), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n980), .B1(new_n979), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT109), .ZN(new_n984));
  INV_X1    g559(.A(new_n977), .ZN(new_n985));
  INV_X1    g560(.A(G8), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n585), .A2(new_n586), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT73), .B1(new_n512), .B2(new_n582), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n590), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n506), .B1(new_n578), .B2(new_n579), .ZN(new_n991));
  OAI21_X1  g566(.A(G1981), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(G1981), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n581), .A2(new_n993), .A3(new_n590), .A4(new_n589), .ZN(new_n994));
  AOI21_X1  g569(.A(KEYINPUT108), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT49), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n987), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  AOI211_X1 g572(.A(KEYINPUT108), .B(KEYINPUT49), .C1(new_n992), .C2(new_n994), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n984), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT108), .ZN(new_n1000));
  AOI22_X1  g575(.A1(new_n550), .A2(G86), .B1(new_n587), .B2(new_n588), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n993), .B1(new_n1001), .B2(new_n581), .ZN(new_n1002));
  NOR3_X1   g577(.A1(new_n990), .A2(G1981), .A3(new_n991), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1000), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(KEYINPUT49), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n995), .A2(new_n996), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n1005), .A2(KEYINPUT109), .A3(new_n1006), .A4(new_n987), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n983), .B1(new_n999), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(G8), .B1(new_n517), .B2(new_n519), .ZN(new_n1009));
  XNOR2_X1  g584(.A(KEYINPUT106), .B(KEYINPUT55), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  OAI221_X1 g586(.A(G8), .B1(KEYINPUT106), .B2(KEYINPUT55), .C1(new_n517), .C2(new_n519), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G1384), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n853), .A2(KEYINPUT45), .A3(new_n1014), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n942), .A2(new_n1015), .A3(new_n975), .ZN(new_n1016));
  XOR2_X1   g591(.A(KEYINPUT105), .B(G1971), .Z(new_n1017));
  OAI21_X1  g592(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT50), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n853), .A2(new_n1019), .A3(new_n1014), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1018), .A2(new_n1020), .A3(new_n975), .ZN(new_n1021));
  OAI22_X1  g596(.A1(new_n1016), .A2(new_n1017), .B1(new_n1021), .B2(G2090), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1013), .B1(new_n1022), .B2(G8), .ZN(new_n1023));
  INV_X1    g598(.A(new_n497), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n496), .B1(new_n629), .B2(new_n493), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1014), .B1(new_n1026), .B2(new_n491), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n943), .B1(new_n1027), .B2(new_n941), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1017), .B1(new_n1028), .B2(new_n1015), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n975), .B1(new_n976), .B2(new_n1019), .ZN(new_n1030));
  NOR3_X1   g605(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1031));
  NOR3_X1   g606(.A1(new_n1030), .A2(new_n1031), .A3(G2090), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n1013), .B(G8), .C1(new_n1029), .C2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT107), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1022), .A2(KEYINPUT107), .A3(G8), .A4(new_n1013), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1023), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(G1966), .B1(new_n1028), .B2(new_n1015), .ZN(new_n1038));
  NOR3_X1   g613(.A1(new_n1030), .A2(new_n1031), .A3(G2084), .ZN(new_n1039));
  OAI21_X1  g614(.A(G8), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n531), .A2(G8), .A3(new_n532), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT119), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n531), .A2(KEYINPUT119), .A3(G8), .A4(new_n532), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  XOR2_X1   g621(.A(KEYINPUT120), .B(KEYINPUT51), .Z(new_n1047));
  NAND3_X1  g622(.A1(new_n1040), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n942), .A2(new_n1015), .A3(new_n975), .ZN(new_n1049));
  INV_X1    g624(.A(G1966), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n943), .B1(new_n1027), .B2(KEYINPUT50), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1052), .A2(new_n762), .A3(new_n1020), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1045), .B1(G8), .B2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g630(.A1(KEYINPUT120), .A2(KEYINPUT51), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1056), .B1(new_n1054), .B2(new_n1045), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1048), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n1008), .A2(new_n1037), .A3(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n942), .A2(new_n1015), .A3(new_n732), .A4(new_n975), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT53), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1028), .A2(KEYINPUT53), .A3(new_n732), .A4(new_n1015), .ZN(new_n1064));
  INV_X1    g639(.A(G1961), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1021), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1063), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(G171), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT123), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1067), .A2(G171), .ZN(new_n1071));
  AOI22_X1  g646(.A1(new_n1069), .A2(new_n1070), .B1(new_n1071), .B2(KEYINPUT122), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1068), .A2(KEYINPUT123), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1060), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(KEYINPUT122), .A2(KEYINPUT54), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1075), .B1(new_n1067), .B2(G171), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n1067), .A2(KEYINPUT121), .A3(G171), .ZN(new_n1077));
  AOI21_X1  g652(.A(KEYINPUT121), .B1(new_n1067), .B2(G171), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1076), .B1(new_n1079), .B2(new_n1060), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1059), .B1(new_n1074), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT57), .ZN(new_n1082));
  AND3_X1   g657(.A1(new_n563), .A2(new_n1082), .A3(new_n570), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1082), .B1(new_n563), .B2(new_n570), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(G1956), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1086), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1087));
  XNOR2_X1  g662(.A(KEYINPUT56), .B(G2072), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n942), .A2(new_n1015), .A3(new_n975), .A4(new_n1088), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n1085), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1084), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n563), .A2(new_n1082), .A3(new_n570), .ZN(new_n1092));
  AOI22_X1  g667(.A1(new_n1087), .A2(new_n1089), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT116), .ZN(new_n1095));
  OAI21_X1  g670(.A(KEYINPUT61), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1098));
  AOI21_X1  g673(.A(G1956), .B1(new_n1052), .B2(new_n1020), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1089), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1098), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1085), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT61), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1101), .B(new_n1102), .C1(KEYINPUT116), .C2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1016), .A2(KEYINPUT112), .A3(new_n951), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT112), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1107), .B1(new_n1049), .B2(G1996), .ZN(new_n1108));
  XOR2_X1   g683(.A(KEYINPUT58), .B(G1341), .Z(new_n1109));
  NAND2_X1  g684(.A1(new_n977), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT113), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n977), .A2(KEYINPUT113), .A3(new_n1109), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1106), .A2(new_n1108), .A3(new_n1112), .A4(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT114), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1115), .A2(KEYINPUT59), .ZN(new_n1116));
  XNOR2_X1  g691(.A(new_n1116), .B(KEYINPUT115), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n624), .B1(new_n1115), .B2(KEYINPUT59), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1114), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1117), .B1(new_n1114), .B2(new_n1118), .ZN(new_n1120));
  OAI22_X1  g695(.A1(new_n1097), .A2(new_n1105), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT117), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  OAI221_X1 g698(.A(KEYINPUT117), .B1(new_n1119), .B2(new_n1120), .C1(new_n1097), .C2(new_n1105), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n614), .A2(KEYINPUT118), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n1021), .A2(new_n711), .B1(new_n985), .B2(new_n947), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT118), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n613), .A2(new_n1127), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1125), .A2(KEYINPUT60), .A3(new_n1126), .A4(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1126), .A2(KEYINPUT60), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1130), .A2(new_n1127), .A3(new_n613), .ZN(new_n1131));
  OR2_X1    g706(.A1(new_n1126), .A2(KEYINPUT60), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1129), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1123), .A2(new_n1124), .A3(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1126), .A2(new_n613), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1102), .B1(new_n1135), .B2(new_n1093), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1081), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1008), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n999), .A2(new_n1007), .ZN(new_n1140));
  NOR2_X1   g715(.A1(G288), .A2(G1976), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1003), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  XOR2_X1   g717(.A(new_n987), .B(KEYINPUT110), .Z(new_n1143));
  OAI21_X1  g718(.A(new_n1139), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT111), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1040), .A2(G286), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1008), .A2(new_n1037), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT63), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1008), .A2(new_n1037), .A3(KEYINPUT63), .A4(new_n1147), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  OAI211_X1 g727(.A(new_n1139), .B(KEYINPUT111), .C1(new_n1142), .C2(new_n1143), .ZN(new_n1153));
  AND3_X1   g728(.A1(new_n1079), .A2(new_n1008), .A3(new_n1037), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT62), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1058), .A2(new_n1155), .ZN(new_n1156));
  OAI211_X1 g731(.A(new_n1048), .B(KEYINPUT62), .C1(new_n1055), .C2(new_n1057), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1154), .A2(new_n1158), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1146), .A2(new_n1152), .A3(new_n1153), .A4(new_n1159), .ZN(new_n1160));
  OAI211_X1 g735(.A(new_n971), .B(new_n974), .C1(new_n1137), .C2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1161), .ZN(new_n1162));
  AND2_X1   g737(.A1(new_n1159), .A2(new_n1153), .ZN(new_n1163));
  AOI22_X1  g738(.A1(new_n1144), .A2(new_n1145), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1136), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1133), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1166), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1165), .B1(new_n1167), .B2(new_n1124), .ZN(new_n1168));
  OAI211_X1 g743(.A(new_n1163), .B(new_n1164), .C1(new_n1168), .C2(new_n1081), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n971), .B1(new_n1169), .B2(new_n974), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n970), .B1(new_n1162), .B2(new_n1170), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g746(.A1(G401), .A2(new_n460), .A3(G227), .ZN(new_n1173));
  INV_X1    g747(.A(new_n1173), .ZN(new_n1174));
  OAI21_X1  g748(.A(new_n1174), .B1(new_n692), .B2(new_n693), .ZN(new_n1175));
  NOR2_X1   g749(.A1(new_n1175), .A2(new_n885), .ZN(new_n1176));
  NAND2_X1  g750(.A1(new_n1176), .A2(new_n929), .ZN(G225));
  INV_X1    g751(.A(G225), .ZN(G308));
endmodule


