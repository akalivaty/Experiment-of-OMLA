//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0 1 0 1 1 0 0 1 0 1 0 1 1 1 0 1 0 1 0 0 0 1 1 0 0 0 1 0 0 1 0 1 0 1 1 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:26 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G143), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  AND2_X1   g004(.A1(KEYINPUT0), .A2(G128), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n188), .A2(new_n190), .A3(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(G143), .B(G146), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT0), .B(G128), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n192), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT66), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT66), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n192), .B(new_n197), .C1(new_n193), .C2(new_n194), .ZN(new_n198));
  OR2_X1    g012(.A1(KEYINPUT64), .A2(G134), .ZN(new_n199));
  INV_X1    g013(.A(G137), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(KEYINPUT11), .ZN(new_n201));
  NAND2_X1  g015(.A1(KEYINPUT64), .A2(G134), .ZN(new_n202));
  AND3_X1   g016(.A1(new_n199), .A2(new_n201), .A3(new_n202), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n200), .A2(KEYINPUT11), .A3(G134), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT11), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G137), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  NOR3_X1   g021(.A1(new_n203), .A2(G131), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G131), .ZN(new_n209));
  AND2_X1   g023(.A1(new_n204), .A2(new_n206), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n199), .A2(new_n201), .A3(new_n202), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  OAI211_X1 g026(.A(new_n196), .B(new_n198), .C1(new_n208), .C2(new_n212), .ZN(new_n213));
  AOI21_X1  g027(.A(G137), .B1(new_n199), .B2(new_n202), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT65), .B1(new_n200), .B2(G134), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT65), .ZN(new_n216));
  INV_X1    g030(.A(G134), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n216), .A2(new_n217), .A3(G137), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(G131), .B1(new_n214), .B2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n210), .A2(new_n209), .A3(new_n211), .ZN(new_n221));
  INV_X1    g035(.A(G128), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n188), .B(new_n190), .C1(KEYINPUT1), .C2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n188), .A2(new_n190), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT1), .B1(new_n189), .B2(G146), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n224), .A2(G128), .A3(new_n225), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n220), .A2(new_n221), .A3(new_n223), .A4(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n213), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G119), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G116), .ZN(new_n230));
  INV_X1    g044(.A(G116), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G119), .ZN(new_n232));
  INV_X1    g046(.A(G113), .ZN(new_n233));
  AND2_X1   g047(.A1(new_n233), .A2(KEYINPUT2), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n233), .A2(KEYINPUT2), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n230), .B(new_n232), .C1(new_n234), .C2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n230), .A2(new_n232), .ZN(new_n237));
  XNOR2_X1  g051(.A(KEYINPUT2), .B(G113), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n236), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n228), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT71), .ZN(new_n242));
  INV_X1    g056(.A(new_n240), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n213), .A2(new_n243), .A3(new_n227), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT70), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n213), .A2(new_n227), .A3(KEYINPUT70), .A4(new_n243), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT71), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n228), .A2(new_n248), .A3(new_n240), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n242), .A2(new_n246), .A3(new_n247), .A4(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT28), .ZN(new_n251));
  XOR2_X1   g065(.A(KEYINPUT67), .B(KEYINPUT27), .Z(new_n252));
  NOR2_X1   g066(.A1(G237), .A2(G953), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G210), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n252), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT26), .B(G101), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n255), .B(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT28), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n244), .A2(new_n259), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n251), .A2(KEYINPUT29), .A3(new_n258), .A4(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT30), .ZN(new_n262));
  AND4_X1   g076(.A1(new_n221), .A2(new_n220), .A3(new_n223), .A4(new_n226), .ZN(new_n263));
  OAI21_X1  g077(.A(G131), .B1(new_n203), .B2(new_n207), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n195), .B1(new_n264), .B2(new_n221), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n262), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n213), .A2(KEYINPUT30), .A3(new_n227), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n266), .A2(new_n240), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(new_n244), .ZN(new_n269));
  AOI21_X1  g083(.A(KEYINPUT29), .B1(new_n269), .B2(new_n257), .ZN(new_n270));
  XNOR2_X1  g084(.A(KEYINPUT68), .B(KEYINPUT28), .ZN(new_n271));
  AND3_X1   g085(.A1(new_n213), .A2(new_n243), .A3(new_n227), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n264), .A2(new_n221), .ZN(new_n273));
  INV_X1    g087(.A(new_n195), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n243), .B1(new_n275), .B2(new_n227), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n271), .B1(new_n272), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n277), .A2(new_n258), .A3(new_n260), .ZN(new_n278));
  AOI21_X1  g092(.A(G902), .B1(new_n270), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n261), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G472), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT32), .ZN(new_n282));
  NOR2_X1   g096(.A1(G472), .A2(G902), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT31), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n268), .A2(new_n284), .A3(new_n244), .A4(new_n258), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n258), .B1(new_n277), .B2(new_n260), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n285), .B1(new_n286), .B2(KEYINPUT69), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n268), .A2(new_n244), .A3(new_n258), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(KEYINPUT31), .ZN(new_n289));
  INV_X1    g103(.A(new_n271), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n240), .B1(new_n263), .B2(new_n265), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n290), .B1(new_n291), .B2(new_n244), .ZN(new_n292));
  AND2_X1   g106(.A1(new_n244), .A2(new_n259), .ZN(new_n293));
  OAI211_X1 g107(.A(KEYINPUT69), .B(new_n257), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n289), .A2(new_n294), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n282), .B(new_n283), .C1(new_n287), .C2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n257), .B1(new_n292), .B2(new_n293), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT69), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n300), .A2(new_n289), .A3(new_n294), .A4(new_n285), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n282), .B1(new_n301), .B2(new_n283), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n281), .B1(new_n297), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G469), .ZN(new_n304));
  INV_X1    g118(.A(G902), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT81), .ZN(new_n306));
  INV_X1    g120(.A(G107), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n306), .B1(new_n307), .B2(G104), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(G104), .ZN(new_n309));
  INV_X1    g123(.A(G104), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n310), .A2(KEYINPUT81), .A3(G107), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n308), .A2(new_n309), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G101), .ZN(new_n313));
  INV_X1    g127(.A(G101), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n310), .A2(G107), .ZN(new_n315));
  AND3_X1   g129(.A1(new_n307), .A2(KEYINPUT3), .A3(G104), .ZN(new_n316));
  AOI21_X1  g130(.A(KEYINPUT3), .B1(new_n307), .B2(G104), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n314), .B(new_n315), .C1(new_n316), .C2(new_n317), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n313), .A2(new_n318), .A3(new_n223), .A4(new_n226), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT10), .ZN(new_n320));
  AOI21_X1  g134(.A(KEYINPUT82), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n319), .A2(KEYINPUT82), .A3(new_n320), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n273), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT4), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n326), .A2(new_n327), .A3(G101), .ZN(new_n328));
  AND3_X1   g142(.A1(new_n196), .A2(new_n198), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n326), .A2(G101), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n330), .A2(KEYINPUT4), .A3(new_n318), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n313), .A2(new_n318), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n226), .A2(new_n223), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI22_X1  g148(.A1(new_n329), .A2(new_n331), .B1(KEYINPUT10), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n324), .A2(new_n325), .A3(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(G110), .B(G140), .ZN(new_n337));
  INV_X1    g151(.A(G227), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n338), .A2(G953), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n337), .B(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  AOI22_X1  g155(.A1(new_n313), .A2(new_n318), .B1(new_n226), .B2(new_n223), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n273), .B1(new_n334), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT12), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n332), .A2(new_n333), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n319), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n347), .A2(KEYINPUT12), .A3(new_n273), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n336), .A2(new_n341), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n334), .A2(KEYINPUT10), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n331), .A2(new_n198), .A3(new_n196), .A4(new_n328), .ZN(new_n352));
  AND3_X1   g166(.A1(new_n319), .A2(KEYINPUT82), .A3(new_n320), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n351), .B(new_n352), .C1(new_n353), .C2(new_n321), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n273), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n341), .B1(new_n355), .B2(new_n336), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n304), .B(new_n305), .C1(new_n350), .C2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(G469), .A2(G902), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n347), .A2(KEYINPUT12), .A3(new_n273), .ZN(new_n359));
  AOI21_X1  g173(.A(KEYINPUT12), .B1(new_n347), .B2(new_n273), .ZN(new_n360));
  OAI22_X1  g174(.A1(new_n354), .A2(new_n273), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n340), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n355), .A2(new_n336), .A3(new_n341), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n362), .A2(G469), .A3(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n357), .A2(new_n358), .A3(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(G214), .B1(G237), .B2(G902), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(G210), .B1(G237), .B2(G902), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT5), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n370), .A2(new_n229), .A3(G116), .ZN(new_n371));
  OAI211_X1 g185(.A(G113), .B(new_n371), .C1(new_n237), .C2(new_n370), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n372), .A2(new_n313), .A3(new_n236), .A4(new_n318), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n318), .A2(KEYINPUT4), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT3), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n375), .B1(new_n310), .B2(G107), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n307), .A2(KEYINPUT3), .A3(G104), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n314), .B1(new_n378), .B2(new_n315), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n374), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n328), .A2(new_n240), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n373), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  XNOR2_X1  g196(.A(G110), .B(G122), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n383), .B(new_n373), .C1(new_n380), .C2(new_n381), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT6), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n387), .A2(KEYINPUT83), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n385), .A2(new_n386), .A3(new_n388), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n382), .B(new_n384), .C1(KEYINPUT83), .C2(new_n387), .ZN(new_n390));
  INV_X1    g204(.A(G125), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n226), .A2(new_n391), .A3(new_n223), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n192), .B(G125), .C1(new_n193), .C2(new_n194), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(G953), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G224), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n394), .B(new_n396), .ZN(new_n397));
  AND3_X1   g211(.A1(new_n389), .A2(new_n390), .A3(new_n397), .ZN(new_n398));
  XOR2_X1   g212(.A(new_n383), .B(KEYINPUT8), .Z(new_n399));
  NAND2_X1  g213(.A1(new_n372), .A2(new_n236), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n332), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n399), .B1(new_n401), .B2(new_n373), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n396), .A2(KEYINPUT7), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n403), .B1(new_n392), .B2(new_n393), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n392), .A2(new_n393), .A3(new_n403), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT84), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n392), .A2(KEYINPUT84), .A3(new_n393), .A4(new_n403), .ZN(new_n409));
  AND2_X1   g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n405), .A2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n386), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n305), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n369), .B1(new_n398), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n408), .A2(new_n409), .ZN(new_n415));
  NOR3_X1   g229(.A1(new_n415), .A2(new_n404), .A3(new_n402), .ZN(new_n416));
  AOI21_X1  g230(.A(G902), .B1(new_n416), .B2(new_n386), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n389), .A2(new_n390), .A3(new_n397), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n417), .A2(new_n368), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n367), .B1(new_n414), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(G221), .ZN(new_n421));
  XOR2_X1   g235(.A(KEYINPUT9), .B(G234), .Z(new_n422));
  AOI21_X1  g236(.A(new_n421), .B1(new_n422), .B2(new_n305), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  AND3_X1   g238(.A1(new_n365), .A2(new_n420), .A3(new_n424), .ZN(new_n425));
  XOR2_X1   g239(.A(KEYINPUT72), .B(G217), .Z(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n427), .B1(G234), .B2(new_n305), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G140), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(G125), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n391), .A2(G140), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n431), .A2(new_n432), .A3(KEYINPUT74), .ZN(new_n433));
  OR3_X1    g247(.A1(new_n391), .A2(KEYINPUT74), .A3(G140), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n433), .A2(new_n434), .A3(KEYINPUT16), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n391), .A2(G140), .ZN(new_n436));
  OR2_X1    g250(.A1(new_n436), .A2(KEYINPUT16), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(G146), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT75), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n435), .A2(new_n187), .A3(new_n437), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n438), .A2(KEYINPUT75), .A3(G146), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n229), .A2(G128), .ZN(new_n444));
  OR2_X1    g258(.A1(new_n444), .A2(KEYINPUT73), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(KEYINPUT73), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n229), .A2(G128), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n445), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  XOR2_X1   g262(.A(KEYINPUT24), .B(G110), .Z(new_n449));
  NAND3_X1  g263(.A1(new_n222), .A2(KEYINPUT23), .A3(G119), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n447), .B(new_n450), .C1(new_n444), .C2(KEYINPUT23), .ZN(new_n451));
  AOI22_X1  g265(.A1(new_n448), .A2(new_n449), .B1(new_n451), .B2(G110), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n442), .A2(new_n443), .A3(new_n452), .ZN(new_n453));
  OAI22_X1  g267(.A1(new_n448), .A2(new_n449), .B1(new_n451), .B2(G110), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n430), .A2(G125), .ZN(new_n455));
  OAI21_X1  g269(.A(KEYINPUT76), .B1(new_n436), .B2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT76), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n431), .A2(new_n432), .A3(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n456), .A2(new_n187), .A3(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n454), .A2(new_n439), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n453), .A2(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(KEYINPUT22), .B(G137), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n395), .A2(G221), .A3(G234), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n462), .B(new_n463), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n464), .B(KEYINPUT77), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n461), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT78), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n453), .A2(new_n460), .A3(new_n464), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n461), .A2(KEYINPUT78), .A3(new_n466), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n469), .A2(new_n305), .A3(new_n470), .A4(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT25), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI211_X1 g288(.A(new_n468), .B(new_n465), .C1(new_n453), .C2(new_n460), .ZN(new_n475));
  INV_X1    g289(.A(new_n470), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n477), .A2(KEYINPUT25), .A3(new_n305), .A4(new_n469), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n429), .B1(new_n474), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(KEYINPUT78), .B1(new_n461), .B2(new_n466), .ZN(new_n480));
  NOR3_X1   g294(.A1(new_n480), .A2(new_n475), .A3(new_n476), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT80), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n428), .A2(G902), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n483), .B(KEYINPUT79), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n481), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n469), .A2(new_n470), .A3(new_n471), .A4(new_n484), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(KEYINPUT80), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n479), .A2(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(G116), .B(G122), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n490), .B(new_n307), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n189), .A2(G128), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT13), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n222), .A2(G143), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n492), .A2(new_n493), .ZN(new_n497));
  OAI21_X1  g311(.A(G134), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n199), .A2(new_n202), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n492), .A2(new_n495), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n491), .B(new_n498), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n499), .B(new_n500), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n490), .A2(new_n307), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n231), .A2(KEYINPUT14), .A3(G122), .ZN(new_n504));
  INV_X1    g318(.A(new_n490), .ZN(new_n505));
  OAI211_X1 g319(.A(G107), .B(new_n504), .C1(new_n505), .C2(KEYINPUT14), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n502), .A2(new_n503), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n501), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n426), .A2(new_n422), .A3(new_n395), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n508), .B(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n305), .ZN(new_n511));
  INV_X1    g325(.A(G478), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n512), .A2(KEYINPUT15), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n510), .B(new_n305), .C1(KEYINPUT15), .C2(new_n512), .ZN(new_n515));
  INV_X1    g329(.A(G952), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n516), .A2(G953), .ZN(new_n517));
  NAND2_X1  g331(.A1(G234), .A2(G237), .ZN(new_n518));
  AND2_X1   g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AND3_X1   g333(.A1(new_n518), .A2(G902), .A3(G953), .ZN(new_n520));
  XNOR2_X1  g334(.A(KEYINPUT21), .B(G898), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n514), .A2(new_n515), .A3(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(G475), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n441), .A2(new_n440), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n187), .B1(new_n435), .B2(new_n437), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n443), .ZN(new_n529));
  INV_X1    g343(.A(G237), .ZN(new_n530));
  AND4_X1   g344(.A1(G143), .A2(new_n530), .A3(new_n395), .A4(G214), .ZN(new_n531));
  AOI21_X1  g345(.A(G143), .B1(new_n253), .B2(G214), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n533), .A2(new_n209), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT17), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n533), .A2(new_n209), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n530), .A2(new_n395), .A3(G214), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(new_n189), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n253), .A2(G143), .A3(G214), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(G131), .ZN(new_n542));
  AOI21_X1  g356(.A(KEYINPUT17), .B1(new_n537), .B2(new_n542), .ZN(new_n543));
  OAI22_X1  g357(.A1(new_n528), .A2(new_n529), .B1(new_n536), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n433), .A2(new_n434), .A3(G146), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n459), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(KEYINPUT18), .A2(G131), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT85), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n548), .B1(new_n533), .B2(new_n549), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n539), .A2(new_n549), .A3(new_n548), .A4(new_n540), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n546), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT86), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n539), .A2(new_n549), .A3(new_n540), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n547), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n551), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n558), .A2(KEYINPUT86), .A3(new_n546), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n544), .A2(new_n560), .ZN(new_n561));
  XNOR2_X1  g375(.A(G113), .B(G122), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n562), .B(new_n310), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n544), .A2(new_n560), .A3(new_n563), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n525), .B1(new_n567), .B2(new_n305), .ZN(new_n568));
  NOR2_X1   g382(.A1(G475), .A2(G902), .ZN(new_n569));
  XOR2_X1   g383(.A(KEYINPUT87), .B(KEYINPUT19), .Z(new_n570));
  NAND3_X1  g384(.A1(new_n456), .A2(new_n458), .A3(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT19), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n433), .A2(new_n434), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n571), .B(new_n187), .C1(new_n572), .C2(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n541), .A2(G131), .ZN(new_n575));
  OAI211_X1 g389(.A(new_n574), .B(new_n439), .C1(new_n534), .C2(new_n575), .ZN(new_n576));
  AND3_X1   g390(.A1(new_n558), .A2(KEYINPUT86), .A3(new_n546), .ZN(new_n577));
  AOI21_X1  g391(.A(KEYINPUT86), .B1(new_n558), .B2(new_n546), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT88), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n579), .A2(new_n580), .A3(new_n564), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n566), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n580), .B1(new_n579), .B2(new_n564), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n569), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(KEYINPUT20), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT20), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n586), .B(new_n569), .C1(new_n582), .C2(new_n583), .ZN(new_n587));
  AOI211_X1 g401(.A(new_n524), .B(new_n568), .C1(new_n585), .C2(new_n587), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n303), .A2(new_n425), .A3(new_n489), .A4(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n589), .B(G101), .ZN(G3));
  AOI21_X1  g404(.A(new_n568), .B1(new_n585), .B2(new_n587), .ZN(new_n591));
  INV_X1    g405(.A(new_n419), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n368), .B1(new_n417), .B2(new_n418), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n366), .B(new_n523), .C1(new_n592), .C2(new_n593), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n509), .A2(KEYINPUT89), .ZN(new_n595));
  OR2_X1    g409(.A1(new_n508), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n508), .A2(new_n595), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n596), .A2(KEYINPUT33), .A3(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT90), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n596), .A2(KEYINPUT90), .A3(KEYINPUT33), .A4(new_n597), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT33), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n510), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n512), .A2(G902), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n600), .A2(new_n601), .A3(new_n603), .A4(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n511), .A2(new_n512), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NOR3_X1   g422(.A1(new_n591), .A2(new_n594), .A3(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n196), .A2(new_n328), .A3(new_n198), .ZN(new_n611));
  OAI22_X1  g425(.A1(new_n611), .A2(new_n380), .B1(new_n320), .B2(new_n319), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n612), .B1(new_n322), .B2(new_n323), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n340), .B1(new_n613), .B2(new_n325), .ZN(new_n614));
  AOI22_X1  g428(.A1(new_n614), .A2(new_n355), .B1(new_n361), .B2(new_n340), .ZN(new_n615));
  OAI21_X1  g429(.A(G469), .B1(new_n615), .B2(G902), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n423), .B1(new_n616), .B2(new_n357), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n301), .A2(new_n305), .ZN(new_n618));
  AOI22_X1  g432(.A1(new_n618), .A2(G472), .B1(new_n283), .B2(new_n301), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n489), .A2(new_n617), .A3(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n610), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(KEYINPUT34), .B(G104), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G6));
  INV_X1    g437(.A(new_n420), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT91), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n585), .A2(new_n625), .A3(new_n587), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n514), .A2(new_n515), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n628), .A2(new_n568), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n527), .B1(new_n542), .B2(new_n537), .ZN(new_n630));
  AOI22_X1  g444(.A1(new_n555), .A2(new_n559), .B1(new_n574), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g445(.A(KEYINPUT88), .B1(new_n631), .B2(new_n563), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n632), .A2(new_n566), .A3(new_n581), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n586), .B1(new_n633), .B2(new_n569), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(KEYINPUT91), .ZN(new_n635));
  AND4_X1   g449(.A1(new_n523), .A2(new_n626), .A3(new_n629), .A4(new_n635), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n624), .B1(new_n636), .B2(KEYINPUT92), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT92), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n626), .A2(new_n629), .A3(new_n635), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n638), .B1(new_n639), .B2(new_n522), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n641), .A2(new_n620), .ZN(new_n642));
  XNOR2_X1  g456(.A(KEYINPUT35), .B(G107), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G9));
  AOI21_X1  g458(.A(KEYINPUT25), .B1(new_n481), .B2(new_n305), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n471), .A2(new_n470), .ZN(new_n646));
  NOR4_X1   g460(.A1(new_n646), .A2(new_n480), .A3(new_n473), .A4(G902), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n428), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n466), .A2(KEYINPUT36), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(new_n461), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n484), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n652), .A2(new_n425), .A3(new_n588), .A4(new_n619), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT37), .B(G110), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(KEYINPUT93), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n653), .B(new_n655), .ZN(G12));
  INV_X1    g470(.A(new_n519), .ZN(new_n657));
  INV_X1    g471(.A(G900), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n520), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n639), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n662), .A2(new_n303), .A3(new_n425), .A4(new_n652), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G128), .ZN(G30));
  XNOR2_X1  g478(.A(new_n660), .B(KEYINPUT39), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n617), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT96), .B(KEYINPUT40), .Z(new_n667));
  OR2_X1    g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(KEYINPUT94), .B(KEYINPUT38), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n670), .B1(new_n592), .B2(new_n593), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n414), .A2(new_n419), .A3(new_n669), .ZN(new_n672));
  AND2_X1   g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n673), .A2(new_n367), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n666), .A2(new_n667), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n591), .A2(new_n628), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n668), .A2(new_n674), .A3(new_n675), .A4(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n250), .A2(new_n257), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n678), .A2(KEYINPUT95), .A3(new_n288), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n305), .ZN(new_n680));
  AOI21_X1  g494(.A(KEYINPUT95), .B1(new_n678), .B2(new_n288), .ZN(new_n681));
  OAI21_X1  g495(.A(G472), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n682), .B1(new_n297), .B2(new_n302), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n650), .A2(new_n484), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n479), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n677), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(new_n189), .ZN(G45));
  NOR3_X1   g502(.A1(new_n591), .A2(new_n608), .A3(new_n661), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n689), .A2(new_n303), .A3(new_n425), .A4(new_n652), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G146), .ZN(G48));
  OAI21_X1  g505(.A(new_n305), .B1(new_n350), .B2(new_n356), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT97), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n693), .A2(new_n304), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  OAI221_X1 g509(.A(new_n305), .B1(new_n693), .B2(new_n304), .C1(new_n350), .C2(new_n356), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n697), .A2(new_n423), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n609), .A2(new_n303), .A3(new_n489), .A4(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(KEYINPUT41), .B(G113), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G15));
  AND3_X1   g515(.A1(new_n303), .A2(new_n489), .A3(new_n698), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n637), .A2(new_n702), .A3(new_n640), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G116), .ZN(G18));
  AND4_X1   g518(.A1(new_n420), .A2(new_n695), .A3(new_n424), .A4(new_n696), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n303), .A2(new_n652), .A3(new_n705), .A4(new_n588), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(KEYINPUT98), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n420), .A2(new_n695), .A3(new_n424), .A4(new_n696), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n567), .A2(new_n305), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(G475), .ZN(new_n710));
  INV_X1    g524(.A(new_n587), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n710), .B1(new_n711), .B2(new_n634), .ZN(new_n712));
  NOR3_X1   g526(.A1(new_n708), .A2(new_n712), .A3(new_n524), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT98), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n713), .A2(new_n714), .A3(new_n303), .A4(new_n652), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n707), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(KEYINPUT99), .B(G119), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G21));
  AOI21_X1  g532(.A(new_n293), .B1(new_n250), .B2(KEYINPUT28), .ZN(new_n719));
  OAI211_X1 g533(.A(KEYINPUT100), .B(new_n289), .C1(new_n719), .C2(new_n258), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n285), .ZN(new_n721));
  AND2_X1   g535(.A1(new_n246), .A2(new_n247), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n248), .B1(new_n228), .B2(new_n240), .ZN(new_n723));
  AOI211_X1 g537(.A(KEYINPUT71), .B(new_n243), .C1(new_n213), .C2(new_n227), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n259), .B1(new_n722), .B2(new_n725), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n257), .B1(new_n726), .B2(new_n293), .ZN(new_n727));
  AOI21_X1  g541(.A(KEYINPUT100), .B1(new_n727), .B2(new_n289), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n283), .B1(new_n721), .B2(new_n728), .ZN(new_n729));
  AND4_X1   g543(.A1(new_n424), .A2(new_n695), .A3(new_n523), .A4(new_n696), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n618), .A2(G472), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n729), .A2(new_n489), .A3(new_n730), .A4(new_n731), .ZN(new_n732));
  OAI21_X1  g546(.A(KEYINPUT101), .B1(new_n591), .B2(new_n628), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT101), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n712), .A2(new_n734), .A3(new_n627), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n733), .A2(new_n420), .A3(new_n735), .ZN(new_n736));
  OR2_X1    g550(.A1(new_n732), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G122), .ZN(G24));
  OAI21_X1  g552(.A(new_n289), .B1(new_n719), .B2(new_n258), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT100), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n741), .A2(new_n285), .A3(new_n720), .ZN(new_n742));
  AOI22_X1  g556(.A1(new_n742), .A2(new_n283), .B1(G472), .B2(new_n618), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n712), .A2(new_n607), .A3(new_n660), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n744), .A2(new_n708), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n743), .A2(new_n745), .A3(new_n652), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G125), .ZN(G27));
  NAND3_X1  g561(.A1(new_n414), .A2(new_n366), .A3(new_n419), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT102), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n414), .A2(KEYINPUT102), .A3(new_n366), .A4(new_n419), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n750), .A2(new_n424), .A3(new_n365), .A4(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n753), .A2(new_n303), .A3(new_n489), .A4(new_n689), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT42), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n283), .B1(new_n287), .B2(new_n295), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(KEYINPUT32), .ZN(new_n758));
  AOI22_X1  g572(.A1(new_n758), .A2(new_n296), .B1(G472), .B2(new_n280), .ZN(new_n759));
  AND2_X1   g573(.A1(new_n485), .A2(new_n487), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n648), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n762), .A2(KEYINPUT42), .A3(new_n689), .A4(new_n753), .ZN(new_n763));
  AND3_X1   g577(.A1(new_n756), .A2(KEYINPUT103), .A3(new_n763), .ZN(new_n764));
  AOI21_X1  g578(.A(KEYINPUT103), .B1(new_n756), .B2(new_n763), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G131), .ZN(G33));
  AOI211_X1 g581(.A(new_n625), .B(new_n586), .C1(new_n633), .C2(new_n569), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n711), .A2(new_n634), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n768), .B1(new_n769), .B2(new_n625), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n770), .A2(KEYINPUT104), .A3(new_n629), .A4(new_n660), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT104), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n772), .B1(new_n639), .B2(new_n661), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n762), .A2(new_n771), .A3(new_n753), .A4(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G134), .ZN(G36));
  INV_X1    g589(.A(new_n665), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n615), .A2(KEYINPUT45), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n362), .A2(new_n363), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT45), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n777), .A2(new_n780), .A3(G469), .ZN(new_n781));
  AOI21_X1  g595(.A(KEYINPUT46), .B1(new_n781), .B2(new_n358), .ZN(new_n782));
  INV_X1    g596(.A(new_n357), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n781), .A2(KEYINPUT46), .A3(new_n358), .ZN(new_n785));
  AOI211_X1 g599(.A(new_n423), .B(new_n776), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT44), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n591), .A2(new_n607), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(KEYINPUT43), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT43), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n591), .A2(new_n790), .A3(new_n607), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(new_n619), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(new_n652), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n787), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n750), .A2(new_n751), .ZN(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n685), .A2(new_n619), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n798), .A2(KEYINPUT44), .A3(new_n789), .A4(new_n791), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n786), .A2(new_n795), .A3(new_n797), .A4(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G137), .ZN(G39));
  AOI21_X1  g615(.A(new_n423), .B1(new_n784), .B2(new_n785), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT47), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n803), .A2(KEYINPUT105), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  NOR4_X1   g620(.A1(new_n303), .A2(new_n744), .A3(new_n489), .A4(new_n796), .ZN(new_n807));
  XNOR2_X1  g621(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n806), .B(new_n807), .C1(new_n802), .C2(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(G140), .ZN(G42));
  NAND2_X1  g624(.A1(new_n617), .A2(new_n420), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n759), .A2(new_n811), .A3(new_n685), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n729), .A2(new_n652), .A3(new_n731), .ZN(new_n813));
  AOI22_X1  g627(.A1(new_n662), .A2(new_n812), .B1(new_n813), .B2(new_n745), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n683), .A2(new_n617), .A3(new_n685), .A4(new_n660), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n815), .A2(new_n736), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT52), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n814), .A2(new_n816), .A3(new_n817), .A4(new_n690), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n746), .A2(new_n663), .A3(new_n690), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n815), .A2(new_n736), .ZN(new_n820));
  OAI21_X1  g634(.A(KEYINPUT52), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  OAI21_X1  g636(.A(KEYINPUT107), .B1(new_n591), .B2(new_n608), .ZN(new_n823));
  INV_X1    g637(.A(new_n594), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT107), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n712), .A2(new_n825), .A3(new_n607), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n823), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n620), .B1(new_n827), .B2(KEYINPUT108), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT108), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n823), .A2(new_n826), .A3(new_n829), .A4(new_n824), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n710), .B(new_n627), .C1(new_n711), .C2(new_n634), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n832), .A2(new_n594), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n833), .A2(new_n489), .A3(new_n617), .A4(new_n619), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n589), .A2(new_n834), .A3(new_n653), .ZN(new_n835));
  INV_X1    g649(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n831), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n759), .A2(new_n685), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n568), .A2(new_n627), .A3(new_n661), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n770), .A2(KEYINPUT109), .A3(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n626), .A2(new_n839), .A3(new_n635), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT109), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n838), .A2(new_n840), .A3(new_n753), .A4(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n743), .A2(new_n652), .A3(new_n753), .A4(new_n689), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n774), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n837), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT110), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n716), .A2(new_n703), .A3(new_n737), .A4(new_n699), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n759), .A2(new_n752), .A3(new_n761), .ZN(new_n851));
  AOI21_X1  g665(.A(KEYINPUT42), .B1(new_n851), .B2(new_n689), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n303), .A2(new_n489), .ZN(new_n853));
  NOR4_X1   g667(.A1(new_n853), .A2(new_n755), .A3(new_n744), .A4(new_n752), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n849), .B1(new_n850), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n699), .B1(new_n732), .B2(new_n736), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n857), .B1(new_n715), .B2(new_n707), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n756), .A2(new_n763), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n858), .A2(KEYINPUT110), .A3(new_n703), .A4(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n822), .A2(new_n848), .A3(new_n856), .A4(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT54), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n818), .A2(new_n821), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT103), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n864), .B1(new_n852), .B2(new_n854), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n774), .A2(new_n844), .A3(new_n845), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n756), .A2(KEYINPUT103), .A3(new_n763), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n835), .B1(new_n830), .B2(new_n828), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n858), .A2(new_n869), .A3(new_n703), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n863), .A2(new_n868), .A3(new_n870), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n861), .B(new_n862), .C1(new_n871), .C2(KEYINPUT53), .ZN(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n850), .A2(new_n837), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n874), .A2(new_n766), .A3(new_n866), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n847), .B1(new_n875), .B2(new_n863), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n868), .A2(new_n870), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n877), .A2(KEYINPUT53), .A3(new_n822), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n862), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n873), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n806), .B1(new_n802), .B2(new_n808), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n881), .B1(new_n424), .B2(new_n697), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n743), .A2(new_n489), .ZN(new_n883));
  OAI21_X1  g697(.A(KEYINPUT111), .B1(new_n792), .B2(new_n657), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT111), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n789), .A2(new_n885), .A3(new_n519), .A4(new_n791), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n883), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n887), .A2(new_n797), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n882), .A2(new_n888), .A3(KEYINPUT112), .ZN(new_n889));
  AOI21_X1  g703(.A(KEYINPUT112), .B1(new_n882), .B2(new_n888), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n698), .A2(new_n367), .A3(new_n673), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n887), .A2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT50), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n887), .A2(KEYINPUT50), .A3(new_n892), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(new_n698), .ZN(new_n898));
  AOI211_X1 g712(.A(new_n898), .B(new_n796), .C1(new_n884), .C2(new_n886), .ZN(new_n899));
  OR2_X1    g713(.A1(new_n683), .A2(new_n761), .ZN(new_n900));
  NOR4_X1   g714(.A1(new_n900), .A2(new_n657), .A3(new_n898), .A4(new_n796), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n712), .A2(new_n607), .ZN(new_n902));
  AOI22_X1  g716(.A1(new_n899), .A2(new_n813), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n897), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(KEYINPUT51), .B1(new_n891), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n887), .A2(new_n705), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n591), .A2(new_n608), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n901), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n906), .A2(new_n517), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(KEYINPUT113), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT113), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n906), .A2(new_n911), .A3(new_n908), .A4(new_n517), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  OR2_X1    g727(.A1(KEYINPUT114), .A2(KEYINPUT48), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n853), .B1(KEYINPUT114), .B2(KEYINPUT48), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n899), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n914), .B1(new_n899), .B2(new_n915), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n897), .A2(new_n903), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n882), .A2(new_n888), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(KEYINPUT51), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n913), .B(new_n918), .C1(new_n919), .C2(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n905), .A2(new_n922), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n880), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(G952), .A2(G953), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n673), .A2(new_n366), .A3(new_n424), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n926), .B1(KEYINPUT49), .B2(new_n697), .ZN(new_n927));
  OR2_X1    g741(.A1(new_n697), .A2(KEYINPUT49), .ZN(new_n928));
  OR2_X1    g742(.A1(new_n928), .A2(KEYINPUT106), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n788), .B1(new_n928), .B2(KEYINPUT106), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n927), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  OAI22_X1  g745(.A1(new_n924), .A2(new_n925), .B1(new_n900), .B2(new_n931), .ZN(G75));
  NOR2_X1   g746(.A1(new_n395), .A2(G952), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(KEYINPUT53), .B1(new_n877), .B2(new_n822), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n856), .A2(new_n860), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n846), .A2(new_n847), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n937), .A2(new_n818), .A3(new_n821), .A4(new_n869), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  OAI211_X1 g753(.A(G210), .B(G902), .C1(new_n935), .C2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT56), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n389), .A2(new_n390), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(new_n397), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT55), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n934), .B1(new_n942), .B2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT117), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n945), .B(KEYINPUT116), .ZN(new_n948));
  XNOR2_X1  g762(.A(KEYINPUT115), .B(KEYINPUT56), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  AND3_X1   g764(.A1(new_n940), .A2(new_n947), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n947), .B1(new_n940), .B2(new_n950), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n946), .A2(new_n953), .ZN(G51));
  XOR2_X1   g768(.A(new_n358), .B(KEYINPUT57), .Z(new_n955));
  AOI21_X1  g769(.A(new_n862), .B1(new_n876), .B2(new_n861), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n955), .B1(new_n873), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n957), .B1(new_n356), .B2(new_n350), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n876), .A2(new_n861), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(G902), .ZN(new_n960));
  OR2_X1    g774(.A1(new_n960), .A2(new_n781), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n933), .B1(new_n958), .B2(new_n961), .ZN(G54));
  INV_X1    g776(.A(new_n633), .ZN(new_n963));
  NAND2_X1  g777(.A1(KEYINPUT58), .A2(G475), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n963), .B1(new_n960), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(new_n934), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n960), .A2(new_n963), .A3(new_n964), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n966), .A2(new_n967), .ZN(G60));
  NAND3_X1  g782(.A1(new_n600), .A2(new_n601), .A3(new_n603), .ZN(new_n969));
  XNOR2_X1  g783(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n512), .A2(new_n305), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n970), .B(new_n971), .Z(new_n972));
  NOR2_X1   g786(.A1(new_n969), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n973), .B1(new_n873), .B2(new_n956), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT119), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n974), .A2(new_n975), .A3(new_n934), .ZN(new_n976));
  INV_X1    g790(.A(new_n973), .ZN(new_n977));
  OAI21_X1  g791(.A(KEYINPUT54), .B1(new_n935), .B2(new_n939), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n977), .B1(new_n978), .B2(new_n872), .ZN(new_n979));
  OAI21_X1  g793(.A(KEYINPUT119), .B1(new_n979), .B2(new_n933), .ZN(new_n980));
  INV_X1    g794(.A(new_n972), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n981), .B1(new_n873), .B2(new_n879), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n969), .ZN(new_n983));
  AND3_X1   g797(.A1(new_n976), .A2(new_n980), .A3(new_n983), .ZN(G63));
  NAND2_X1  g798(.A1(G217), .A2(G902), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT60), .Z(new_n986));
  NAND2_X1  g800(.A1(new_n959), .A2(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(new_n481), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n959), .A2(new_n650), .A3(new_n986), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n989), .A2(new_n934), .A3(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT61), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n989), .A2(KEYINPUT61), .A3(new_n934), .A4(new_n990), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(G66));
  NAND2_X1  g809(.A1(new_n870), .A2(new_n395), .ZN(new_n996));
  INV_X1    g810(.A(G224), .ZN(new_n997));
  OAI21_X1  g811(.A(G953), .B1(new_n521), .B2(new_n997), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n996), .A2(KEYINPUT120), .A3(new_n998), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n999), .B1(KEYINPUT120), .B2(new_n996), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n943), .B1(G898), .B2(new_n395), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1001), .B(KEYINPUT121), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1000), .B(new_n1002), .ZN(G69));
  INV_X1    g817(.A(new_n819), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n800), .A2(KEYINPUT124), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(new_n1005), .ZN(new_n1006));
  AOI21_X1  g820(.A(KEYINPUT124), .B1(new_n800), .B2(new_n1004), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n736), .A2(new_n853), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n786), .A2(new_n1009), .ZN(new_n1010));
  AND3_X1   g824(.A1(new_n809), .A2(new_n774), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1011), .A2(new_n766), .ZN(new_n1012));
  OAI21_X1  g826(.A(KEYINPUT125), .B1(new_n1008), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(new_n1007), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1014), .A2(new_n1005), .ZN(new_n1015));
  INV_X1    g829(.A(KEYINPUT125), .ZN(new_n1016));
  NAND4_X1  g830(.A1(new_n1015), .A2(new_n1016), .A3(new_n766), .A4(new_n1011), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n1013), .A2(new_n1017), .A3(new_n395), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n266), .A2(new_n267), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n1020));
  XOR2_X1   g834(.A(new_n1019), .B(new_n1020), .Z(new_n1021));
  AOI21_X1  g835(.A(new_n1021), .B1(G900), .B2(G953), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1018), .A2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g837(.A(G953), .B1(new_n338), .B2(new_n658), .ZN(new_n1024));
  XNOR2_X1  g838(.A(new_n1024), .B(KEYINPUT123), .ZN(new_n1025));
  NOR2_X1   g839(.A1(new_n1025), .A2(KEYINPUT126), .ZN(new_n1026));
  AND2_X1   g840(.A1(new_n823), .A2(new_n826), .ZN(new_n1027));
  INV_X1    g841(.A(new_n832), .ZN(new_n1028));
  OAI211_X1 g842(.A(new_n851), .B(new_n665), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1029));
  AND3_X1   g843(.A1(new_n809), .A2(new_n1029), .A3(new_n800), .ZN(new_n1030));
  OAI21_X1  g844(.A(KEYINPUT62), .B1(new_n687), .B2(new_n819), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1031), .A2(KEYINPUT122), .ZN(new_n1032));
  INV_X1    g846(.A(KEYINPUT122), .ZN(new_n1033));
  OAI211_X1 g847(.A(new_n1033), .B(KEYINPUT62), .C1(new_n687), .C2(new_n819), .ZN(new_n1034));
  OR3_X1    g848(.A1(new_n687), .A2(KEYINPUT62), .A3(new_n819), .ZN(new_n1035));
  NAND4_X1  g849(.A1(new_n1030), .A2(new_n1032), .A3(new_n1034), .A4(new_n1035), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1036), .A2(new_n395), .ZN(new_n1037));
  AOI21_X1  g851(.A(new_n1026), .B1(new_n1037), .B2(new_n1021), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1025), .A2(KEYINPUT126), .ZN(new_n1039));
  AND3_X1   g853(.A1(new_n1023), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g854(.A(new_n1039), .B1(new_n1023), .B2(new_n1038), .ZN(new_n1041));
  NOR2_X1   g855(.A1(new_n1040), .A2(new_n1041), .ZN(G72));
  NAND3_X1  g856(.A1(new_n1013), .A2(new_n1017), .A3(new_n874), .ZN(new_n1043));
  NAND2_X1  g857(.A1(G472), .A2(G902), .ZN(new_n1044));
  XOR2_X1   g858(.A(new_n1044), .B(KEYINPUT63), .Z(new_n1045));
  NAND2_X1  g859(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g860(.A1(new_n269), .A2(new_n258), .ZN(new_n1047));
  NAND2_X1  g861(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g862(.A1(new_n876), .A2(new_n878), .ZN(new_n1049));
  INV_X1    g863(.A(new_n1047), .ZN(new_n1050));
  NAND2_X1  g864(.A1(new_n269), .A2(new_n258), .ZN(new_n1051));
  NAND4_X1  g865(.A1(new_n1049), .A2(new_n1045), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  OAI21_X1  g866(.A(new_n1045), .B1(new_n1036), .B2(new_n870), .ZN(new_n1053));
  INV_X1    g867(.A(new_n1051), .ZN(new_n1054));
  AOI21_X1  g868(.A(new_n933), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND4_X1  g869(.A1(new_n1048), .A2(KEYINPUT127), .A3(new_n1052), .A4(new_n1055), .ZN(new_n1056));
  INV_X1    g870(.A(KEYINPUT127), .ZN(new_n1057));
  NAND2_X1  g871(.A1(new_n1052), .A2(new_n1055), .ZN(new_n1058));
  AOI21_X1  g872(.A(new_n1050), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1059));
  OAI21_X1  g873(.A(new_n1057), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g874(.A1(new_n1056), .A2(new_n1060), .ZN(G57));
endmodule


