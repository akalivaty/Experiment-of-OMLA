//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 1 1 1 1 0 0 0 1 0 1 1 0 1 0 1 0 1 0 1 0 0 0 1 0 0 1 0 1 1 1 0 1 0 1 0 0 1 1 1 1 0 1 1 1 0 1 1 0 1 1 0 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:46 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1303,
    new_n1304, new_n1305, new_n1306, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1374, new_n1375, new_n1376, new_n1377,
    new_n1378, new_n1379, new_n1380, new_n1381, new_n1382, new_n1383,
    new_n1384, new_n1385, new_n1386, new_n1387;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n201), .A2(G77), .A3(new_n203), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  AND2_X1   g0012(.A1(KEYINPUT65), .A2(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(KEYINPUT65), .A2(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n203), .A2(G50), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  INV_X1    g0021(.A(G68), .ZN(new_n222));
  INV_X1    g0022(.A(G238), .ZN(new_n223));
  INV_X1    g0023(.A(G87), .ZN(new_n224));
  INV_X1    g0024(.A(G250), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n227));
  INV_X1    g0027(.A(G77), .ZN(new_n228));
  INV_X1    g0028(.A(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G107), .ZN(new_n230));
  INV_X1    g0030(.A(G264), .ZN(new_n231));
  OAI221_X1 g0031(.A(new_n227), .B1(new_n228), .B2(new_n229), .C1(new_n230), .C2(new_n231), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n209), .B1(new_n226), .B2(new_n232), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n212), .B(new_n220), .C1(KEYINPUT1), .C2(new_n233), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n233), .ZN(G361));
  XOR2_X1   g0035(.A(G238), .B(G244), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XOR2_X1   g0037(.A(KEYINPUT2), .B(G226), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G264), .B(G270), .Z(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XOR2_X1   g0044(.A(G107), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G68), .B(G77), .Z(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n246), .B(new_n249), .Z(G351));
  AOI21_X1  g0050(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT66), .ZN(new_n252));
  INV_X1    g0052(.A(G1698), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT3), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n259));
  NAND4_X1  g0059(.A1(new_n254), .A2(new_n256), .A3(new_n258), .A4(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G222), .ZN(new_n261));
  AND2_X1   g0061(.A1(new_n256), .A2(new_n258), .ZN(new_n262));
  OAI22_X1  g0062(.A1(new_n260), .A2(new_n261), .B1(new_n262), .B2(new_n228), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n256), .A2(new_n258), .ZN(new_n264));
  INV_X1    g0064(.A(G223), .ZN(new_n265));
  NOR3_X1   g0065(.A1(new_n264), .A2(new_n265), .A3(new_n253), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n251), .B1(new_n263), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G41), .ZN(new_n268));
  INV_X1    g0068(.A(G45), .ZN(new_n269));
  AOI21_X1  g0069(.A(G1), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(G33), .A2(G41), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n271), .A2(G1), .A3(G13), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n270), .A2(new_n272), .A3(G274), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n251), .A2(new_n270), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n274), .B1(G226), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n267), .A2(new_n276), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n277), .A2(G179), .ZN(new_n278));
  AND2_X1   g0078(.A1(new_n278), .A2(KEYINPUT69), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n278), .A2(KEYINPUT69), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n216), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n215), .A2(G33), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT8), .ZN(new_n285));
  INV_X1    g0085(.A(G58), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n285), .B1(new_n286), .B2(KEYINPUT67), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT67), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n288), .A2(KEYINPUT8), .A3(G58), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G150), .ZN(new_n291));
  NOR2_X1   g0091(.A1(G20), .A2(G33), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  OAI22_X1  g0093(.A1(new_n284), .A2(new_n290), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT68), .ZN(new_n295));
  AND2_X1   g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(G20), .B1(new_n201), .B2(new_n203), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n297), .B1(new_n294), .B2(new_n295), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n283), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G13), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n300), .A2(G1), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G20), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n302), .A2(G50), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n283), .B1(new_n206), .B2(G20), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n303), .B1(new_n304), .B2(G50), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n299), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n277), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n306), .B1(G169), .B2(new_n307), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n281), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G190), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n277), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n311), .B1(G200), .B2(new_n277), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n306), .A2(KEYINPUT9), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT9), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n314), .B1(new_n299), .B2(new_n305), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n312), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT10), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT10), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n318), .B(new_n312), .C1(new_n313), .C2(new_n315), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n309), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  AND2_X1   g0120(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n321));
  NOR2_X1   g0121(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n262), .A2(G232), .A3(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n262), .A2(G238), .A3(G1698), .ZN(new_n325));
  AND2_X1   g0125(.A1(KEYINPUT70), .A2(G107), .ZN(new_n326));
  NOR2_X1   g0126(.A1(KEYINPUT70), .A2(G107), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n324), .B(new_n325), .C1(new_n328), .C2(new_n262), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n251), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n274), .B1(G244), .B2(new_n275), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n330), .A2(KEYINPUT71), .A3(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(KEYINPUT71), .B1(new_n330), .B2(new_n331), .ZN(new_n334));
  OAI21_X1  g0134(.A(G190), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n334), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n336), .A2(G200), .A3(new_n332), .ZN(new_n337));
  XNOR2_X1  g0137(.A(KEYINPUT15), .B(G87), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n284), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g0139(.A(KEYINPUT8), .B(G58), .ZN(new_n340));
  OAI22_X1  g0140(.A1(new_n215), .A2(new_n228), .B1(new_n340), .B2(new_n293), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n283), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n302), .A2(G77), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n343), .B1(new_n304), .B2(G77), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n335), .A2(new_n337), .A3(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(G179), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n348), .B1(new_n333), .B2(new_n334), .ZN(new_n349));
  INV_X1    g0149(.A(G169), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n336), .A2(new_n350), .A3(new_n332), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n349), .A2(new_n351), .A3(new_n345), .ZN(new_n352));
  AND2_X1   g0152(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  AND3_X1   g0153(.A1(new_n320), .A2(KEYINPUT72), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(KEYINPUT72), .B1(new_n320), .B2(new_n353), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n292), .A2(G50), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n207), .A2(G68), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n357), .B1(KEYINPUT75), .B2(new_n358), .ZN(new_n359));
  OAI221_X1 g0159(.A(new_n359), .B1(KEYINPUT75), .B2(new_n357), .C1(new_n284), .C2(new_n228), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n283), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT11), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n360), .A2(KEYINPUT11), .A3(new_n283), .ZN(new_n364));
  OR3_X1    g0164(.A1(new_n302), .A2(KEYINPUT12), .A3(G68), .ZN(new_n365));
  OAI21_X1  g0165(.A(KEYINPUT12), .B1(new_n302), .B2(G68), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n365), .A2(new_n366), .B1(G68), .B2(new_n304), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n363), .A2(new_n364), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(G33), .A2(G97), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n256), .A2(new_n258), .A3(G232), .A4(G1698), .ZN(new_n370));
  INV_X1    g0170(.A(G226), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n369), .B(new_n370), .C1(new_n260), .C2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n251), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n272), .A2(G238), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n273), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n373), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(KEYINPUT13), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n376), .B1(new_n372), .B2(new_n251), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT13), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT74), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n378), .A2(KEYINPUT74), .A3(KEYINPUT13), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n368), .B1(new_n385), .B2(G190), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n380), .A2(new_n381), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n379), .A2(KEYINPUT73), .A3(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT73), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n380), .A2(new_n389), .A3(new_n381), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n388), .A2(G200), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n386), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT76), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n386), .A2(KEYINPUT76), .A3(new_n391), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n388), .A2(G169), .A3(new_n390), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n397), .A2(KEYINPUT14), .B1(new_n385), .B2(G179), .ZN(new_n398));
  OAI21_X1  g0198(.A(KEYINPUT73), .B1(new_n380), .B2(new_n381), .ZN(new_n399));
  XNOR2_X1  g0199(.A(new_n399), .B(new_n387), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT14), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n400), .A2(KEYINPUT77), .A3(new_n401), .A4(G169), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n388), .A2(new_n401), .A3(G169), .A4(new_n390), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT77), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n398), .A2(new_n402), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n368), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT18), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT16), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT7), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n410), .B1(new_n264), .B2(new_n215), .ZN(new_n411));
  AOI211_X1 g0211(.A(KEYINPUT7), .B(G20), .C1(new_n256), .C2(new_n258), .ZN(new_n412));
  NOR3_X1   g0212(.A1(new_n411), .A2(new_n412), .A3(new_n222), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n286), .A2(new_n222), .ZN(new_n414));
  OAI21_X1  g0214(.A(G20), .B1(new_n414), .B2(new_n202), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n292), .A2(G159), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n409), .B1(new_n413), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(KEYINPUT78), .B1(new_n257), .B2(G33), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT78), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n420), .A2(new_n255), .A3(KEYINPUT3), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n419), .A2(new_n421), .A3(new_n258), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n207), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n222), .B1(new_n423), .B2(KEYINPUT7), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT79), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n419), .A2(new_n421), .A3(KEYINPUT79), .A4(new_n258), .ZN(new_n427));
  OR2_X1    g0227(.A1(KEYINPUT65), .A2(G20), .ZN(new_n428));
  NAND2_X1  g0228(.A1(KEYINPUT65), .A2(G20), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n430), .A2(KEYINPUT7), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n426), .A2(new_n427), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n424), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n417), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n283), .B(new_n418), .C1(new_n435), .C2(new_n409), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n290), .A2(new_n302), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n437), .B1(new_n304), .B2(new_n290), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n274), .B1(G232), .B2(new_n275), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n254), .A2(new_n259), .ZN(new_n441));
  OAI22_X1  g0241(.A1(new_n441), .A2(new_n265), .B1(new_n371), .B2(new_n253), .ZN(new_n442));
  AND3_X1   g0242(.A1(new_n419), .A2(new_n421), .A3(new_n258), .ZN(new_n443));
  AOI22_X1  g0243(.A1(new_n442), .A2(new_n443), .B1(G33), .B2(G87), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n440), .B(G179), .C1(new_n444), .C2(new_n272), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n275), .A2(G232), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n273), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n323), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n448));
  OAI22_X1  g0248(.A1(new_n448), .A2(new_n422), .B1(new_n255), .B2(new_n224), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n447), .B1(new_n449), .B2(new_n251), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n445), .B1(new_n450), .B2(new_n350), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n408), .B1(new_n439), .B2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n438), .ZN(new_n453));
  INV_X1    g0253(.A(new_n283), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n417), .B1(new_n424), .B2(new_n432), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n454), .B1(new_n455), .B2(KEYINPUT16), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n453), .B1(new_n456), .B2(new_n418), .ZN(new_n457));
  INV_X1    g0257(.A(new_n451), .ZN(new_n458));
  NOR3_X1   g0258(.A1(new_n457), .A2(new_n458), .A3(KEYINPUT18), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n452), .A2(new_n459), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n440), .B(G190), .C1(new_n444), .C2(new_n272), .ZN(new_n461));
  INV_X1    g0261(.A(G200), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n461), .B1(new_n450), .B2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  AND3_X1   g0264(.A1(new_n457), .A2(KEYINPUT17), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(KEYINPUT17), .B1(new_n457), .B2(new_n464), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n396), .A2(new_n407), .A3(new_n460), .A4(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n356), .A2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT19), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n428), .A2(G33), .A3(G97), .A4(new_n429), .ZN(new_n471));
  NAND3_X1  g0271(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n428), .A2(new_n429), .A3(new_n472), .ZN(new_n473));
  OR2_X1    g0273(.A1(KEYINPUT70), .A2(G107), .ZN(new_n474));
  NOR2_X1   g0274(.A1(G87), .A2(G97), .ZN(new_n475));
  NAND2_X1  g0275(.A1(KEYINPUT70), .A2(G107), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n474), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n470), .A2(new_n471), .B1(new_n473), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n443), .A2(G68), .A3(new_n215), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n454), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n338), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n481), .A2(new_n302), .ZN(new_n482));
  OAI21_X1  g0282(.A(KEYINPUT81), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n471), .A2(new_n470), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n473), .A2(new_n477), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NOR3_X1   g0286(.A1(new_n422), .A2(new_n222), .A3(new_n430), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n283), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT81), .ZN(new_n489));
  INV_X1    g0289(.A(new_n482), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n483), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n272), .A2(G274), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n269), .A2(G1), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n495), .A2(new_n225), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n494), .A2(new_n495), .B1(new_n272), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(G33), .A2(G116), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  OAI22_X1  g0299(.A1(new_n441), .A2(new_n223), .B1(new_n229), .B2(new_n253), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n499), .B1(new_n500), .B2(new_n443), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n497), .B1(new_n501), .B2(new_n272), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G200), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n206), .A2(G33), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n454), .A2(new_n302), .A3(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n505), .A2(new_n224), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n496), .A2(new_n272), .ZN(new_n508));
  INV_X1    g0308(.A(new_n495), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n508), .B1(new_n509), .B2(new_n493), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n323), .A2(G238), .B1(G244), .B2(G1698), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n498), .B1(new_n511), .B2(new_n422), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n510), .B1(new_n512), .B2(new_n251), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(G190), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n492), .A2(new_n503), .A3(new_n507), .A4(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n502), .A2(G169), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n516), .B1(new_n348), .B2(new_n502), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n505), .A2(new_n338), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n518), .B1(new_n483), .B2(new_n491), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n517), .B1(new_n519), .B2(KEYINPUT82), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT82), .ZN(new_n521));
  AOI211_X1 g0321(.A(new_n521), .B(new_n518), .C1(new_n483), .C2(new_n491), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n515), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT83), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  OAI211_X1 g0325(.A(KEYINPUT83), .B(new_n515), .C1(new_n520), .C2(new_n522), .ZN(new_n526));
  XNOR2_X1  g0326(.A(KEYINPUT5), .B(G41), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n527), .A2(G274), .A3(new_n272), .A4(new_n495), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n251), .B1(new_n495), .B2(new_n527), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(G264), .ZN(new_n530));
  INV_X1    g0330(.A(G294), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n255), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(G257), .A2(G1698), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(new_n441), .B2(new_n225), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n532), .B1(new_n534), .B2(new_n443), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n528), .B(new_n530), .C1(new_n535), .C2(new_n272), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT85), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n536), .A2(new_n537), .A3(G169), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n323), .A2(G250), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n422), .B1(new_n539), .B2(new_n533), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n251), .B1(new_n540), .B2(new_n532), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n541), .A2(G179), .A3(new_n528), .A4(new_n530), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n537), .B1(new_n536), .B2(G169), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT22), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n428), .A2(G87), .A3(new_n429), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n545), .B1(new_n546), .B2(new_n264), .ZN(new_n547));
  NOR2_X1   g0347(.A1(KEYINPUT23), .A2(G107), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n430), .A2(new_n548), .B1(new_n207), .B2(new_n499), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n474), .A2(new_n476), .ZN(new_n550));
  OAI21_X1  g0350(.A(KEYINPUT23), .B1(new_n550), .B2(new_n207), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n547), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  NOR4_X1   g0352(.A1(new_n422), .A2(new_n430), .A3(new_n545), .A4(new_n224), .ZN(new_n553));
  OAI21_X1  g0353(.A(KEYINPUT24), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n548), .ZN(new_n555));
  OAI22_X1  g0355(.A1(new_n215), .A2(new_n555), .B1(G20), .B2(new_n498), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT23), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n557), .B1(new_n328), .B2(G20), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n443), .A2(KEYINPUT22), .A3(G87), .A4(new_n215), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT24), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n559), .A2(new_n560), .A3(new_n561), .A4(new_n547), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n454), .B1(new_n554), .B2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT25), .ZN(new_n564));
  NOR3_X1   g0364(.A1(new_n302), .A2(new_n564), .A3(G107), .ZN(new_n565));
  NOR3_X1   g0365(.A1(new_n300), .A2(new_n207), .A3(G1), .ZN(new_n566));
  AOI21_X1  g0366(.A(KEYINPUT25), .B1(new_n566), .B2(new_n230), .ZN(new_n567));
  OAI22_X1  g0367(.A1(new_n565), .A2(new_n567), .B1(new_n230), .B2(new_n505), .ZN(new_n568));
  OAI22_X1  g0368(.A1(new_n543), .A2(new_n544), .B1(new_n563), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n554), .A2(new_n562), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n568), .B1(new_n570), .B2(new_n283), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n536), .A2(new_n462), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n541), .A2(new_n310), .A3(new_n528), .A4(new_n530), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n572), .A2(KEYINPUT86), .A3(new_n573), .ZN(new_n574));
  OR3_X1    g0374(.A1(new_n536), .A2(KEYINPUT86), .A3(G190), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n571), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n254), .A2(G244), .A3(new_n259), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(KEYINPUT4), .B1(new_n443), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(G33), .A2(G283), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n256), .A2(new_n258), .A3(G250), .A4(G1698), .ZN(new_n581));
  NAND2_X1  g0381(.A1(KEYINPUT4), .A2(G244), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n580), .B(new_n581), .C1(new_n260), .C2(new_n582), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n251), .B1(new_n579), .B2(new_n583), .ZN(new_n584));
  AND2_X1   g0384(.A1(KEYINPUT5), .A2(G41), .ZN(new_n585));
  NOR2_X1   g0385(.A1(KEYINPUT5), .A2(G41), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n495), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n272), .ZN(new_n588));
  INV_X1    g0388(.A(G257), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n528), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n584), .A2(new_n591), .A3(G179), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT4), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n593), .B1(new_n422), .B2(new_n577), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n262), .A2(KEYINPUT4), .A3(G244), .A4(new_n323), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n594), .A2(new_n595), .A3(new_n580), .A4(new_n581), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n590), .B1(new_n596), .B2(new_n251), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n592), .B1(new_n597), .B2(new_n350), .ZN(new_n598));
  OAI21_X1  g0398(.A(KEYINPUT7), .B1(new_n262), .B2(new_n430), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n264), .A2(new_n410), .A3(new_n207), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n599), .A2(new_n550), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n292), .A2(G77), .ZN(new_n602));
  XNOR2_X1  g0402(.A(KEYINPUT80), .B(G107), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(G97), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n605), .A2(new_n230), .A3(KEYINPUT6), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(KEYINPUT6), .B2(new_n605), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n603), .B(new_n606), .C1(KEYINPUT6), .C2(new_n605), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n608), .A2(new_n609), .A3(new_n430), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n601), .A2(new_n602), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n283), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n302), .A2(G97), .ZN(new_n613));
  AND3_X1   g0413(.A1(new_n454), .A2(new_n302), .A3(new_n504), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n613), .B1(new_n614), .B2(G97), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n598), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n597), .A2(G190), .ZN(new_n618));
  INV_X1    g0418(.A(new_n615), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n619), .B1(new_n611), .B2(new_n283), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n618), .B(new_n620), .C1(new_n462), .C2(new_n597), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n569), .A2(new_n576), .A3(new_n617), .A4(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(G270), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n528), .B1(new_n588), .B2(new_n623), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n231), .A2(new_n253), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n443), .A2(KEYINPUT84), .A3(new_n625), .ZN(new_n626));
  NOR3_X1   g0426(.A1(new_n321), .A2(new_n322), .A3(new_n589), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n443), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT84), .ZN(new_n629));
  INV_X1    g0429(.A(new_n625), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n629), .B1(new_n422), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n264), .A2(G303), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n626), .A2(new_n628), .A3(new_n631), .A4(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n624), .B1(new_n633), .B2(new_n251), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n255), .A2(G97), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n428), .A2(new_n635), .A3(new_n429), .A4(new_n580), .ZN(new_n636));
  INV_X1    g0436(.A(G116), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n282), .A2(new_n216), .B1(G20), .B2(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(KEYINPUT20), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n636), .A2(KEYINPUT20), .A3(new_n638), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n302), .A2(G116), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n643), .B1(new_n614), .B2(G116), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n348), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n634), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT21), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n350), .B1(new_n642), .B2(new_n644), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n633), .A2(new_n251), .ZN(new_n649));
  OAI211_X1 g0449(.A(new_n647), .B(new_n648), .C1(new_n649), .C2(new_n624), .ZN(new_n650));
  INV_X1    g0450(.A(new_n641), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n651), .A2(new_n639), .ZN(new_n652));
  INV_X1    g0452(.A(new_n643), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n653), .B1(new_n505), .B2(new_n637), .ZN(new_n654));
  OAI21_X1  g0454(.A(G169), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(KEYINPUT21), .B1(new_n634), .B2(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n646), .B1(new_n650), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n634), .A2(G190), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n652), .A2(new_n654), .ZN(new_n659));
  OAI211_X1 g0459(.A(new_n658), .B(new_n659), .C1(new_n462), .C2(new_n634), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n622), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n469), .A2(new_n525), .A3(new_n526), .A4(new_n662), .ZN(new_n663));
  XNOR2_X1  g0463(.A(new_n663), .B(KEYINPUT87), .ZN(G372));
  NAND2_X1  g0464(.A1(new_n317), .A2(new_n319), .ZN(new_n665));
  INV_X1    g0465(.A(new_n467), .ZN(new_n666));
  INV_X1    g0466(.A(new_n352), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n396), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n666), .B1(new_n668), .B2(new_n407), .ZN(new_n669));
  INV_X1    g0469(.A(new_n460), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n665), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n309), .ZN(new_n672));
  AND2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n617), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n525), .A2(new_n526), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(KEYINPUT26), .ZN(new_n676));
  AOI221_X4 g0476(.A(new_n506), .B1(new_n513), .B2(G190), .C1(new_n483), .C2(new_n491), .ZN(new_n677));
  OAI21_X1  g0477(.A(KEYINPUT88), .B1(new_n513), .B2(new_n462), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT88), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n502), .A2(new_n679), .A3(G200), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n519), .ZN(new_n682));
  AOI22_X1  g0482(.A1(new_n677), .A2(new_n681), .B1(new_n682), .B2(new_n517), .ZN(new_n683));
  AND3_X1   g0483(.A1(new_n584), .A2(G179), .A3(new_n591), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n350), .B1(new_n584), .B2(new_n591), .ZN(new_n685));
  OAI21_X1  g0485(.A(KEYINPUT89), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT89), .ZN(new_n687));
  OAI211_X1 g0487(.A(new_n592), .B(new_n687), .C1(new_n597), .C2(new_n350), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n686), .A2(new_n616), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT90), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT26), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n686), .A2(KEYINPUT90), .A3(new_n616), .A4(new_n688), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n683), .A2(new_n691), .A3(new_n692), .A4(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n682), .A2(new_n517), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n657), .A2(new_n569), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n621), .A2(new_n617), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n681), .A2(new_n492), .A3(new_n507), .A4(new_n514), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n696), .A2(new_n576), .A3(new_n697), .A4(new_n698), .ZN(new_n699));
  AND3_X1   g0499(.A1(new_n694), .A2(new_n695), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n676), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n469), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n673), .A2(new_n702), .ZN(G369));
  NAND2_X1  g0503(.A1(new_n215), .A2(new_n301), .ZN(new_n704));
  OR2_X1    g0504(.A1(new_n704), .A2(KEYINPUT27), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(KEYINPUT27), .ZN(new_n706));
  AND3_X1   g0506(.A1(new_n705), .A2(G213), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(G343), .ZN(new_n708));
  XNOR2_X1  g0508(.A(new_n708), .B(KEYINPUT91), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n657), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n710), .B(KEYINPUT92), .ZN(new_n711));
  INV_X1    g0511(.A(new_n709), .ZN(new_n712));
  OAI211_X1 g0512(.A(new_n569), .B(new_n576), .C1(new_n712), .C2(new_n571), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(new_n569), .B2(new_n712), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n569), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n716), .B1(new_n717), .B2(new_n712), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n712), .A2(new_n659), .ZN(new_n719));
  INV_X1    g0519(.A(new_n657), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n721), .B1(new_n661), .B2(new_n719), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(G330), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(new_n714), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n718), .A2(new_n725), .ZN(G399));
  INV_X1    g0526(.A(new_n210), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(G41), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n328), .A2(new_n637), .A3(new_n475), .ZN(new_n729));
  NOR3_X1   g0529(.A1(new_n728), .A2(new_n206), .A3(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT93), .ZN(new_n731));
  AOI22_X1  g0531(.A1(new_n730), .A2(new_n731), .B1(new_n219), .B2(new_n728), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n732), .B1(new_n731), .B2(new_n730), .ZN(new_n733));
  XOR2_X1   g0533(.A(KEYINPUT94), .B(KEYINPUT28), .Z(new_n734));
  XNOR2_X1  g0534(.A(new_n733), .B(new_n734), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n662), .A2(new_n525), .A3(new_n526), .A4(new_n712), .ZN(new_n736));
  INV_X1    g0536(.A(new_n536), .ZN(new_n737));
  OAI21_X1  g0537(.A(KEYINPUT95), .B1(new_n737), .B2(new_n597), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n502), .A2(new_n348), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(new_n634), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n584), .A2(new_n591), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT95), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n741), .A2(new_n742), .A3(new_n536), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n738), .A2(new_n740), .A3(new_n743), .ZN(new_n744));
  AOI211_X1 g0544(.A(new_n348), .B(new_n510), .C1(new_n512), .C2(new_n251), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n588), .A2(new_n231), .ZN(new_n746));
  AOI22_X1  g0546(.A1(new_n323), .A2(G250), .B1(G257), .B2(G1698), .ZN(new_n747));
  OAI22_X1  g0547(.A1(new_n747), .A2(new_n422), .B1(new_n255), .B2(new_n531), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n746), .B1(new_n748), .B2(new_n251), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n745), .A2(new_n634), .A3(new_n749), .A4(new_n597), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT30), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  AND3_X1   g0552(.A1(new_n749), .A2(new_n513), .A3(G179), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n753), .A2(KEYINPUT30), .A3(new_n634), .A4(new_n597), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n744), .A2(new_n752), .A3(new_n754), .ZN(new_n755));
  AND3_X1   g0555(.A1(new_n755), .A2(KEYINPUT31), .A3(new_n709), .ZN(new_n756));
  AOI21_X1  g0556(.A(KEYINPUT31), .B1(new_n755), .B2(new_n709), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n736), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G330), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT96), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(G330), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n763), .B1(new_n736), .B2(new_n758), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(KEYINPUT96), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n701), .A2(new_n712), .ZN(new_n768));
  INV_X1    g0568(.A(KEYINPUT29), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g0570(.A1(new_n525), .A2(new_n692), .A3(new_n526), .A4(new_n674), .ZN(new_n771));
  AND4_X1   g0571(.A1(new_n576), .A2(new_n698), .A3(new_n617), .A4(new_n621), .ZN(new_n772));
  AOI22_X1  g0572(.A1(new_n772), .A2(new_n696), .B1(new_n682), .B2(new_n517), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n683), .A2(new_n691), .A3(new_n693), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(KEYINPUT26), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n771), .A2(new_n773), .A3(new_n775), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n776), .A2(KEYINPUT29), .A3(new_n712), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n767), .B1(new_n770), .B2(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n735), .B1(new_n778), .B2(G1), .ZN(G364));
  NOR2_X1   g0579(.A1(new_n430), .A2(new_n300), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G45), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G1), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n728), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n724), .A2(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n784), .B1(G330), .B2(new_n722), .ZN(new_n785));
  INV_X1    g0585(.A(new_n783), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n727), .A2(new_n264), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n787), .A2(G355), .B1(new_n637), .B2(new_n727), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n426), .A2(new_n427), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n727), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n219), .A2(new_n269), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n792), .B1(new_n249), .B2(new_n269), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n788), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(G13), .A2(G33), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(G20), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n216), .B1(G20), .B2(new_n350), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n786), .B1(new_n794), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n310), .A2(G200), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n215), .B1(new_n348), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(new_n605), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n430), .A2(G179), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(G200), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT97), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n807), .A2(G190), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n803), .B1(new_n808), .B2(G68), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT99), .ZN(new_n810));
  NOR2_X1   g0610(.A1(G190), .A2(G200), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n430), .A2(new_n348), .A3(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(G159), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  XOR2_X1   g0614(.A(KEYINPUT98), .B(KEYINPUT32), .Z(new_n815));
  XNOR2_X1  g0615(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n348), .A2(G20), .A3(G190), .A4(G200), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n262), .B1(new_n817), .B2(new_n224), .ZN(new_n818));
  NOR3_X1   g0618(.A1(new_n804), .A2(new_n310), .A3(G200), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n818), .B1(new_n819), .B2(G58), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n805), .A2(new_n811), .ZN(new_n821));
  NOR4_X1   g0621(.A1(new_n215), .A2(G179), .A3(G190), .A4(new_n462), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n820), .B1(new_n228), .B2(new_n821), .C1(new_n230), .C2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n807), .A2(new_n310), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n816), .B(new_n824), .C1(G50), .C2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(G303), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n264), .B1(new_n827), .B2(new_n817), .C1(new_n802), .C2(new_n531), .ZN(new_n828));
  INV_X1    g0628(.A(new_n812), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n819), .A2(G322), .B1(G329), .B2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(G283), .ZN(new_n831));
  INV_X1    g0631(.A(G311), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n830), .B1(new_n831), .B2(new_n823), .C1(new_n832), .C2(new_n821), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n828), .B(new_n833), .C1(G326), .C2(new_n825), .ZN(new_n834));
  XNOR2_X1  g0634(.A(KEYINPUT33), .B(G317), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n808), .A2(new_n835), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n810), .A2(new_n826), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n798), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n800), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  XOR2_X1   g0639(.A(new_n839), .B(KEYINPUT100), .Z(new_n840));
  INV_X1    g0640(.A(new_n797), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n722), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n785), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  XOR2_X1   g0643(.A(new_n843), .B(KEYINPUT101), .Z(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(G396));
  NOR2_X1   g0645(.A1(new_n798), .A2(new_n795), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n783), .B1(G77), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n819), .ZN(new_n849));
  OAI22_X1  g0649(.A1(new_n849), .A2(new_n531), .B1(new_n832), .B2(new_n812), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n823), .A2(new_n224), .B1(new_n821), .B2(new_n637), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n264), .B1(new_n817), .B2(new_n230), .ZN(new_n852));
  NOR4_X1   g0652(.A1(new_n850), .A2(new_n851), .A3(new_n803), .A4(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n808), .ZN(new_n854));
  INV_X1    g0654(.A(new_n825), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n853), .B1(new_n854), .B2(new_n831), .C1(new_n827), .C2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n821), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n857), .A2(G159), .B1(new_n819), .B2(G143), .ZN(new_n858));
  INV_X1    g0658(.A(G137), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n858), .B1(new_n854), .B2(new_n291), .C1(new_n859), .C2(new_n855), .ZN(new_n860));
  XOR2_X1   g0660(.A(new_n860), .B(KEYINPUT34), .Z(new_n861));
  NOR2_X1   g0661(.A1(new_n823), .A2(new_n222), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n862), .B1(G132), .B2(new_n829), .ZN(new_n863));
  INV_X1    g0663(.A(new_n802), .ZN(new_n864));
  INV_X1    g0664(.A(new_n817), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n864), .A2(G58), .B1(new_n865), .B2(G50), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n863), .A2(new_n789), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n856), .B1(new_n861), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n848), .B1(new_n868), .B2(new_n798), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n709), .A2(new_n345), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n347), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n352), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n667), .A2(new_n712), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n795), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n869), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n768), .A2(new_n874), .ZN(new_n877));
  INV_X1    g0677(.A(new_n874), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n701), .A2(new_n712), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n881), .A2(new_n767), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  OR2_X1    g0683(.A1(new_n883), .A2(KEYINPUT102), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n786), .B1(new_n880), .B2(new_n766), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n885), .B1(new_n883), .B2(KEYINPUT102), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n876), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(G384));
  NOR2_X1   g0688(.A1(new_n780), .A2(new_n206), .ZN(new_n889));
  INV_X1    g0689(.A(new_n873), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n709), .B1(new_n676), .B2(new_n700), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n890), .B1(new_n891), .B2(new_n878), .ZN(new_n892));
  AND3_X1   g0692(.A1(new_n406), .A2(KEYINPUT103), .A3(new_n368), .ZN(new_n893));
  AOI21_X1  g0693(.A(KEYINPUT103), .B1(new_n406), .B2(new_n368), .ZN(new_n894));
  INV_X1    g0694(.A(new_n368), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n712), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n385), .A2(G190), .ZN(new_n898));
  AND4_X1   g0698(.A1(KEYINPUT76), .A2(new_n898), .A3(new_n895), .A4(new_n391), .ZN(new_n899));
  AOI21_X1  g0699(.A(KEYINPUT76), .B1(new_n386), .B2(new_n391), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n897), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NOR3_X1   g0701(.A1(new_n893), .A2(new_n894), .A3(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n406), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n897), .B1(new_n396), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n892), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n707), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT104), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n409), .B1(new_n455), .B2(new_n908), .ZN(new_n909));
  AOI211_X1 g0709(.A(KEYINPUT104), .B(new_n417), .C1(new_n424), .C2(new_n432), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n456), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n907), .B1(new_n911), .B2(new_n438), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n913), .B1(new_n460), .B2(new_n467), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT105), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n457), .A2(new_n464), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n435), .A2(KEYINPUT104), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n455), .A2(new_n908), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n918), .A2(new_n409), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n453), .B1(new_n920), .B2(new_n456), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n917), .B1(new_n921), .B2(new_n907), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n458), .B1(new_n911), .B2(new_n438), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n916), .B(KEYINPUT37), .C1(new_n922), .C2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n439), .A2(new_n451), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n439), .A2(new_n707), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n925), .A2(new_n926), .A3(new_n917), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n927), .A2(KEYINPUT37), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n924), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n911), .A2(new_n438), .ZN(new_n930));
  AOI22_X1  g0730(.A1(new_n930), .A2(new_n707), .B1(new_n457), .B2(new_n464), .ZN(new_n931));
  INV_X1    g0731(.A(new_n923), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n916), .B1(new_n933), .B2(KEYINPUT37), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n915), .B1(new_n929), .B2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT38), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OAI211_X1 g0737(.A(KEYINPUT38), .B(new_n915), .C1(new_n929), .C2(new_n934), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n906), .A2(new_n939), .B1(new_n670), .B2(new_n907), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n927), .B(KEYINPUT37), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n460), .A2(new_n467), .ZN(new_n942));
  INV_X1    g0742(.A(new_n926), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n936), .ZN(new_n946));
  AOI21_X1  g0746(.A(KEYINPUT39), .B1(new_n938), .B2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n937), .A2(KEYINPUT39), .A3(new_n938), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT103), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n407), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n406), .A2(KEYINPUT103), .A3(new_n368), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n709), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n948), .A2(new_n949), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n940), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n770), .A2(new_n469), .A3(new_n777), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(new_n673), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n955), .B(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n759), .A2(new_n878), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n896), .B1(new_n394), .B2(new_n395), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n951), .A2(new_n952), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n396), .A2(new_n903), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n896), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n959), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(KEYINPUT40), .B1(new_n939), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n938), .A2(new_n946), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n874), .B1(new_n736), .B2(new_n758), .ZN(new_n967));
  OAI211_X1 g0767(.A(KEYINPUT40), .B(new_n967), .C1(new_n902), .C2(new_n904), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n965), .B1(new_n966), .B2(new_n969), .ZN(new_n970));
  AND2_X1   g0770(.A1(new_n469), .A2(new_n759), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n763), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n970), .B2(new_n971), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n889), .B1(new_n958), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(new_n958), .B2(new_n973), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n608), .A2(new_n609), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT35), .ZN(new_n977));
  OAI211_X1 g0777(.A(G116), .B(new_n217), .C1(new_n976), .C2(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n978), .B1(new_n977), .B2(new_n976), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT36), .Z(new_n980));
  NOR3_X1   g0780(.A1(new_n218), .A2(new_n228), .A3(new_n414), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n201), .A2(new_n222), .ZN(new_n982));
  OAI211_X1 g0782(.A(G1), .B(new_n300), .C1(new_n981), .C2(new_n982), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n975), .A2(new_n980), .A3(new_n983), .ZN(G367));
  NAND2_X1  g0784(.A1(new_n492), .A2(new_n507), .ZN(new_n985));
  AND2_X1   g0785(.A1(new_n709), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n695), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n683), .B2(new_n986), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT106), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT43), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n989), .A2(new_n990), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n697), .B1(new_n620), .B2(new_n712), .ZN(new_n993));
  AND2_X1   g0793(.A1(new_n993), .A2(KEYINPUT107), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n993), .A2(KEYINPUT107), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n994), .A2(new_n995), .B1(new_n689), .B2(new_n712), .ZN(new_n996));
  AND2_X1   g0796(.A1(new_n996), .A2(KEYINPUT108), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n996), .A2(KEYINPUT108), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n716), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT42), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1000), .A2(new_n717), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n709), .B1(new_n1003), .B2(new_n617), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n991), .B(new_n992), .C1(new_n1002), .C2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n999), .A2(new_n725), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1001), .B(KEYINPUT42), .Z(new_n1007));
  INV_X1    g0807(.A(new_n1004), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1007), .A2(new_n990), .A3(new_n989), .A4(new_n1008), .ZN(new_n1009));
  AND3_X1   g0809(.A1(new_n1005), .A2(new_n1006), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1006), .B1(new_n1009), .B2(new_n1005), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n728), .B(KEYINPUT41), .Z(new_n1013));
  INV_X1    g0813(.A(new_n718), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n999), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT44), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1015), .B(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1000), .A2(KEYINPUT45), .A3(new_n718), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT45), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n1014), .B2(new_n999), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n725), .B1(new_n1017), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n711), .A2(new_n714), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1024), .B(new_n715), .C1(new_n724), .C2(KEYINPUT109), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n724), .A2(KEYINPUT109), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1025), .B(new_n1026), .Z(new_n1027));
  NAND3_X1  g0827(.A1(new_n1017), .A2(new_n725), .A3(new_n1021), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1023), .A2(new_n778), .A3(new_n1027), .A4(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1013), .B1(new_n1029), .B2(new_n778), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1012), .B1(new_n782), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n989), .A2(new_n797), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n799), .B1(new_n210), .B2(new_n338), .C1(new_n791), .C2(new_n242), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(new_n783), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT110), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n808), .A2(G159), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n825), .A2(G143), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n262), .B1(new_n817), .B2(new_n286), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(new_n829), .B2(G137), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n823), .A2(new_n228), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n201), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n821), .A2(new_n1041), .B1(new_n802), .B2(new_n222), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n1040), .B(new_n1042), .C1(G150), .C2(new_n819), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1036), .A2(new_n1037), .A3(new_n1039), .A4(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n829), .A2(G317), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1045), .B1(new_n328), .B2(new_n802), .C1(new_n823), .C2(new_n605), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n865), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT46), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(new_n817), .B2(new_n637), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1047), .B(new_n1049), .C1(new_n821), .C2(new_n831), .ZN(new_n1050));
  NOR3_X1   g0850(.A1(new_n1046), .A2(new_n789), .A3(new_n1050), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(KEYINPUT111), .B(G311), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n825), .A2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n827), .B2(new_n849), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(KEYINPUT112), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1051), .B(new_n1055), .C1(new_n531), .C2(new_n854), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1054), .A2(KEYINPUT112), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1044), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT47), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n798), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1032), .B(new_n1035), .C1(new_n1060), .C2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1031), .A2(new_n1063), .ZN(G387));
  INV_X1    g0864(.A(new_n728), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(new_n778), .B2(new_n1027), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(new_n778), .B2(new_n1027), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n714), .A2(new_n841), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n239), .A2(new_n269), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n1069), .A2(new_n790), .B1(new_n729), .B2(new_n787), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n340), .ZN(new_n1071));
  INV_X1    g0871(.A(G50), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT50), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n269), .B1(new_n222), .B2(new_n228), .ZN(new_n1075));
  NOR3_X1   g0875(.A1(new_n1074), .A2(new_n729), .A3(new_n1075), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n1070), .A2(new_n1076), .B1(G107), .B2(new_n210), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n799), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n783), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n849), .A2(new_n1072), .B1(new_n291), .B2(new_n812), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n865), .A2(G77), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n789), .B(new_n1081), .C1(new_n823), .C2(new_n605), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n802), .A2(new_n338), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n821), .A2(new_n222), .ZN(new_n1084));
  NOR4_X1   g0884(.A1(new_n1080), .A2(new_n1082), .A3(new_n1083), .A4(new_n1084), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n1085), .B1(new_n854), .B2(new_n290), .C1(new_n813), .C2(new_n855), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT113), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n789), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(G116), .A2(new_n822), .B1(new_n829), .B2(G326), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n802), .A2(new_n831), .B1(new_n531), .B2(new_n817), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n808), .A2(new_n1052), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n825), .A2(G322), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n857), .A2(G303), .B1(new_n819), .B2(G317), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT48), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1090), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(new_n1095), .B2(new_n1094), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT49), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1088), .B(new_n1089), .C1(new_n1097), .C2(new_n1098), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1087), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n1068), .B(new_n1079), .C1(new_n1101), .C2(new_n798), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(new_n1027), .B2(new_n782), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1067), .A2(new_n1103), .ZN(G393));
  NAND2_X1  g0904(.A1(new_n778), .A2(new_n1027), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1028), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1105), .B1(new_n1106), .B2(new_n1022), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1029), .A2(new_n1107), .A3(new_n728), .ZN(new_n1108));
  AND2_X1   g0908(.A1(new_n790), .A2(new_n246), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n799), .B1(new_n605), .B2(new_n210), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n808), .A2(new_n201), .B1(new_n1071), .B2(new_n857), .ZN(new_n1111));
  AND2_X1   g0911(.A1(new_n1111), .A2(KEYINPUT114), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1111), .A2(KEYINPUT114), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n802), .A2(new_n228), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(G143), .B2(new_n829), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n822), .A2(G87), .B1(G68), .B2(new_n865), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1115), .A2(new_n789), .A3(new_n1116), .ZN(new_n1117));
  NOR3_X1   g0917(.A1(new_n1112), .A2(new_n1113), .A3(new_n1117), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n825), .A2(G150), .B1(G159), .B2(new_n819), .ZN(new_n1119));
  XOR2_X1   g0919(.A(new_n1119), .B(KEYINPUT51), .Z(new_n1120));
  AOI22_X1  g0920(.A1(new_n825), .A2(G317), .B1(G311), .B2(new_n819), .ZN(new_n1121));
  XOR2_X1   g0921(.A(new_n1121), .B(KEYINPUT52), .Z(new_n1122));
  OAI221_X1 g0922(.A(new_n264), .B1(new_n817), .B2(new_n831), .C1(new_n823), .C2(new_n230), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n864), .A2(G116), .B1(new_n829), .B2(G322), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n531), .B2(new_n821), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n1123), .B(new_n1125), .C1(new_n808), .C2(G303), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n1118), .A2(new_n1120), .B1(new_n1122), .B2(new_n1126), .ZN(new_n1127));
  OAI221_X1 g0927(.A(new_n783), .B1(new_n1109), .B2(new_n1110), .C1(new_n1127), .C2(new_n838), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(new_n999), .B2(new_n797), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1106), .A2(new_n1022), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1129), .B1(new_n1130), .B2(new_n782), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1108), .A2(new_n1131), .ZN(G390));
  NAND3_X1  g0932(.A1(new_n776), .A2(new_n712), .A3(new_n872), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n873), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT115), .ZN(new_n1135));
  AND3_X1   g0935(.A1(new_n961), .A2(new_n963), .A3(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1135), .B1(new_n961), .B2(new_n963), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1134), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n953), .B1(new_n938), .B2(new_n946), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n927), .A2(KEYINPUT37), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT37), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(new_n931), .B2(new_n932), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1141), .B1(new_n1143), .B2(new_n916), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n464), .A2(new_n436), .A3(new_n438), .ZN(new_n1145));
  NOR3_X1   g0945(.A1(new_n912), .A2(new_n923), .A3(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(KEYINPUT105), .B1(new_n1146), .B2(new_n1142), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n936), .B(new_n914), .C1(new_n1144), .C2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1147), .A2(new_n928), .A3(new_n924), .ZN(new_n1149));
  AOI21_X1  g0949(.A(KEYINPUT38), .B1(new_n1149), .B2(new_n915), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n947), .B1(new_n1151), .B2(KEYINPUT39), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n879), .A2(new_n873), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n961), .A2(new_n963), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n953), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1140), .B1(new_n1152), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n967), .A2(G330), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n905), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n762), .A2(new_n765), .A3(new_n878), .A4(new_n1154), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1140), .B(new_n1160), .C1(new_n1152), .C2(new_n1155), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1159), .A2(new_n782), .A3(new_n1161), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n802), .A2(new_n813), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n865), .A2(G150), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1164), .B(KEYINPUT53), .ZN(new_n1165));
  AOI211_X1 g0965(.A(new_n1163), .B(new_n1165), .C1(G125), .C2(new_n829), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n264), .B1(new_n819), .B2(G132), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(KEYINPUT54), .B(G143), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n857), .A2(new_n1169), .B1(new_n201), .B2(new_n822), .ZN(new_n1170));
  AND3_X1   g0970(.A1(new_n1166), .A2(new_n1167), .A3(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(G128), .ZN(new_n1172));
  OAI221_X1 g0972(.A(new_n1171), .B1(new_n1172), .B2(new_n855), .C1(new_n859), .C2(new_n854), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n849), .A2(new_n637), .B1(new_n802), .B2(new_n228), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n821), .A2(new_n605), .B1(new_n531), .B2(new_n812), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n264), .B1(new_n817), .B2(new_n224), .ZN(new_n1176));
  NOR4_X1   g0976(.A1(new_n1174), .A2(new_n1175), .A3(new_n862), .A4(new_n1176), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n1177), .B1(new_n854), .B2(new_n328), .C1(new_n831), .C2(new_n855), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n838), .B1(new_n1173), .B2(new_n1178), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n786), .B(new_n1179), .C1(new_n290), .C2(new_n846), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n1152), .B2(new_n796), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1162), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n948), .A2(new_n949), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n953), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1185), .B1(new_n892), .B2(new_n905), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n1184), .A2(new_n1186), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1158), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1161), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1137), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n961), .A2(new_n963), .A3(new_n1135), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1190), .A2(new_n1191), .A3(new_n1157), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1134), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1192), .A2(new_n1160), .A3(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n762), .A2(new_n765), .A3(new_n878), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1158), .B1(new_n1195), .B2(new_n905), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1194), .B1(new_n1196), .B2(new_n892), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n469), .A2(new_n764), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n956), .A2(new_n673), .A3(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1197), .A2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1065), .B1(new_n1189), .B2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT116), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1159), .A2(new_n1161), .A3(new_n1200), .A4(new_n1197), .ZN(new_n1204));
  AND3_X1   g1004(.A1(new_n1202), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1203), .B1(new_n1202), .B2(new_n1204), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1183), .B1(new_n1205), .B2(new_n1206), .ZN(G378));
  NAND2_X1  g1007(.A1(new_n306), .A2(new_n707), .ZN(new_n1208));
  AND2_X1   g1008(.A1(new_n320), .A2(new_n1208), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n320), .A2(new_n1208), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  OR3_X1    g1012(.A1(new_n1209), .A2(new_n1210), .A3(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1212), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(KEYINPUT38), .B1(new_n941), .B2(new_n944), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n914), .B1(new_n1144), .B2(new_n1147), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1216), .B1(new_n1217), .B2(KEYINPUT38), .ZN(new_n1218));
  OAI21_X1  g1018(.A(G330), .B1(new_n1218), .B2(new_n968), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT40), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1154), .A2(new_n967), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1221), .B1(new_n1151), .B2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1215), .B1(new_n1220), .B2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1215), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(new_n965), .A2(new_n1219), .A3(new_n1225), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n955), .B1(new_n1224), .B2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1220), .A2(new_n1223), .A3(new_n1215), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1225), .B1(new_n965), .B2(new_n1219), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1228), .A2(new_n1229), .A3(new_n954), .A4(new_n940), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1227), .A2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n782), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n786), .B1(new_n1041), .B2(new_n846), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n825), .A2(G125), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n808), .A2(G132), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n864), .A2(G150), .B1(new_n865), .B2(new_n1169), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n857), .A2(G137), .B1(new_n819), .B2(G128), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1234), .A2(new_n1235), .A3(new_n1236), .A4(new_n1237), .ZN(new_n1238));
  OR2_X1    g1038(.A1(new_n1238), .A2(KEYINPUT59), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(KEYINPUT59), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(G33), .A2(G41), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(new_n1241), .B(KEYINPUT117), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n823), .A2(new_n813), .ZN(new_n1243));
  AOI211_X1 g1043(.A(new_n1242), .B(new_n1243), .C1(G124), .C2(new_n829), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1239), .A2(new_n1240), .A3(new_n1244), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n789), .A2(G41), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n822), .A2(G58), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n829), .A2(G283), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1246), .A2(new_n1081), .A3(new_n1247), .A4(new_n1248), .ZN(new_n1249));
  XOR2_X1   g1049(.A(new_n1249), .B(KEYINPUT118), .Z(new_n1250));
  AOI22_X1  g1050(.A1(new_n857), .A2(new_n481), .B1(G68), .B2(new_n864), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1251), .B1(new_n230), .B2(new_n849), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(G97), .B2(new_n808), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n1250), .B(new_n1253), .C1(new_n637), .C2(new_n855), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT58), .ZN(new_n1255));
  OR2_X1    g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1072), .B(new_n1242), .C1(new_n789), .C2(G41), .ZN(new_n1258));
  AND4_X1   g1058(.A1(new_n1245), .A2(new_n1256), .A3(new_n1257), .A4(new_n1258), .ZN(new_n1259));
  OAI221_X1 g1059(.A(new_n1233), .B1(new_n838), .B2(new_n1259), .C1(new_n1215), .C2(new_n796), .ZN(new_n1260));
  AND2_X1   g1060(.A1(new_n1232), .A2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT57), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1262), .B1(new_n1227), .B2(new_n1230), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1200), .B1(new_n1189), .B2(new_n1201), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n728), .ZN(new_n1266));
  AOI21_X1  g1066(.A(KEYINPUT57), .B1(new_n1264), .B2(new_n1231), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1261), .B1(new_n1266), .B2(new_n1267), .ZN(G375));
  NAND2_X1  g1068(.A1(new_n1197), .A2(new_n782), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1190), .A2(new_n795), .A3(new_n1191), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n783), .B1(G68), .B2(new_n847), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1083), .B1(G303), .B2(new_n829), .ZN(new_n1272));
  OAI221_X1 g1072(.A(new_n1272), .B1(new_n831), .B2(new_n849), .C1(new_n328), .C2(new_n821), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n264), .B1(new_n817), .B2(new_n605), .ZN(new_n1274));
  NOR3_X1   g1074(.A1(new_n1273), .A2(new_n1040), .A3(new_n1274), .ZN(new_n1275));
  OAI221_X1 g1075(.A(new_n1275), .B1(new_n637), .B2(new_n854), .C1(new_n531), .C2(new_n855), .ZN(new_n1276));
  XNOR2_X1  g1076(.A(new_n1276), .B(KEYINPUT119), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n825), .A2(G132), .ZN(new_n1278));
  OAI221_X1 g1078(.A(new_n1278), .B1(new_n859), .B2(new_n849), .C1(new_n854), .C2(new_n1168), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT120), .ZN(new_n1280));
  AND2_X1   g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  AOI22_X1  g1081(.A1(new_n857), .A2(G150), .B1(G50), .B2(new_n864), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1282), .B1(new_n1172), .B2(new_n812), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1247), .B1(new_n813), .B2(new_n817), .ZN(new_n1284));
  NOR3_X1   g1084(.A1(new_n1283), .A2(new_n1088), .A3(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1285), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1277), .B1(new_n1281), .B2(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1271), .B1(new_n1287), .B2(new_n798), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1270), .A2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1269), .A2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1013), .ZN(new_n1292));
  OAI211_X1 g1092(.A(new_n1199), .B(new_n1194), .C1(new_n892), .C2(new_n1196), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1201), .A2(new_n1292), .A3(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1291), .A2(new_n1294), .ZN(new_n1295));
  XOR2_X1   g1095(.A(new_n1295), .B(KEYINPUT121), .Z(G381));
  NAND3_X1  g1096(.A1(new_n1067), .A2(new_n844), .A3(new_n1103), .ZN(new_n1297));
  NOR3_X1   g1097(.A1(G390), .A2(G384), .A3(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1182), .B1(new_n1204), .B2(new_n1202), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1298), .A2(new_n1031), .A3(new_n1063), .A4(new_n1299), .ZN(new_n1300));
  XNOR2_X1  g1100(.A(G375), .B(KEYINPUT122), .ZN(new_n1301));
  OR3_X1    g1101(.A1(new_n1300), .A2(new_n1301), .A3(G381), .ZN(G407));
  INV_X1    g1102(.A(G343), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(G213), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1299), .A2(new_n1305), .ZN(new_n1306));
  OAI211_X1 g1106(.A(G407), .B(G213), .C1(new_n1301), .C2(new_n1306), .ZN(G409));
  NAND2_X1  g1107(.A1(new_n1264), .A2(new_n1231), .ZN(new_n1308));
  OAI211_X1 g1108(.A(new_n1232), .B(new_n1260), .C1(new_n1308), .C2(new_n1013), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(new_n1299), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1189), .A2(new_n1201), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1311), .A2(new_n1204), .A3(new_n728), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(KEYINPUT116), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1202), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1182), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT123), .ZN(new_n1316));
  NOR3_X1   g1116(.A1(G375), .A2(new_n1315), .A3(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1232), .A2(new_n1260), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1308), .A2(new_n1262), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1065), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1318), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1321));
  AOI21_X1  g1121(.A(KEYINPUT123), .B1(new_n1321), .B2(G378), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1310), .B1(new_n1317), .B2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT125), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT60), .ZN(new_n1325));
  OR3_X1    g1125(.A1(new_n1293), .A2(new_n1324), .A3(new_n1325), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1324), .B1(new_n1293), .B2(new_n1325), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  XNOR2_X1  g1128(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1293), .A2(new_n1329), .ZN(new_n1330));
  AND3_X1   g1130(.A1(new_n1330), .A2(new_n728), .A3(new_n1201), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1328), .A2(new_n1331), .ZN(new_n1332));
  AOI21_X1  g1132(.A(G384), .B1(new_n1332), .B2(new_n1291), .ZN(new_n1333));
  AOI211_X1 g1133(.A(new_n1290), .B(new_n887), .C1(new_n1328), .C2(new_n1331), .ZN(new_n1334));
  NOR2_X1   g1134(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1323), .A2(new_n1304), .A3(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1336), .A2(KEYINPUT62), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT61), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT62), .ZN(new_n1339));
  NAND4_X1  g1139(.A1(new_n1323), .A2(new_n1339), .A3(new_n1304), .A4(new_n1335), .ZN(new_n1340));
  INV_X1    g1140(.A(new_n1333), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1332), .A2(G384), .A3(new_n1291), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1305), .A2(G2897), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1341), .A2(new_n1342), .A3(new_n1343), .ZN(new_n1344));
  OAI211_X1 g1144(.A(G2897), .B(new_n1305), .C1(new_n1333), .C2(new_n1334), .ZN(new_n1345));
  INV_X1    g1145(.A(new_n1310), .ZN(new_n1346));
  OAI21_X1  g1146(.A(new_n1316), .B1(G375), .B2(new_n1315), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1321), .A2(G378), .A3(KEYINPUT123), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1346), .B1(new_n1347), .B2(new_n1348), .ZN(new_n1349));
  OAI211_X1 g1149(.A(new_n1344), .B(new_n1345), .C1(new_n1349), .C2(new_n1305), .ZN(new_n1350));
  NAND4_X1  g1150(.A1(new_n1337), .A2(new_n1338), .A3(new_n1340), .A4(new_n1350), .ZN(new_n1351));
  INV_X1    g1151(.A(new_n1297), .ZN(new_n1352));
  AOI21_X1  g1152(.A(new_n844), .B1(new_n1067), .B2(new_n1103), .ZN(new_n1353));
  NOR2_X1   g1153(.A1(new_n1352), .A2(new_n1353), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(G390), .A2(new_n1354), .ZN(new_n1355));
  OAI211_X1 g1155(.A(new_n1108), .B(new_n1131), .C1(new_n1352), .C2(new_n1353), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1355), .A2(new_n1356), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(G387), .A2(new_n1357), .ZN(new_n1358));
  NAND4_X1  g1158(.A1(new_n1031), .A2(new_n1355), .A3(new_n1063), .A4(new_n1356), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1358), .A2(new_n1359), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1351), .A2(new_n1360), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1344), .A2(new_n1345), .ZN(new_n1362));
  AOI21_X1  g1162(.A(new_n1362), .B1(new_n1323), .B2(new_n1304), .ZN(new_n1363));
  NOR3_X1   g1163(.A1(new_n1363), .A2(KEYINPUT61), .A3(new_n1360), .ZN(new_n1364));
  INV_X1    g1164(.A(KEYINPUT126), .ZN(new_n1365));
  INV_X1    g1165(.A(new_n1335), .ZN(new_n1366));
  NOR3_X1   g1166(.A1(new_n1349), .A2(new_n1305), .A3(new_n1366), .ZN(new_n1367));
  OAI21_X1  g1167(.A(new_n1365), .B1(new_n1367), .B2(KEYINPUT63), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1367), .A2(KEYINPUT63), .ZN(new_n1369));
  INV_X1    g1169(.A(KEYINPUT63), .ZN(new_n1370));
  NAND3_X1  g1170(.A1(new_n1336), .A2(KEYINPUT126), .A3(new_n1370), .ZN(new_n1371));
  NAND4_X1  g1171(.A1(new_n1364), .A2(new_n1368), .A3(new_n1369), .A4(new_n1371), .ZN(new_n1372));
  NAND2_X1  g1172(.A1(new_n1361), .A2(new_n1372), .ZN(G405));
  NAND2_X1  g1173(.A1(new_n1347), .A2(new_n1348), .ZN(new_n1374));
  NAND2_X1  g1174(.A1(G375), .A2(new_n1299), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(new_n1374), .A2(new_n1375), .ZN(new_n1376));
  NAND2_X1  g1176(.A1(new_n1376), .A2(KEYINPUT127), .ZN(new_n1377));
  INV_X1    g1177(.A(KEYINPUT127), .ZN(new_n1378));
  NAND3_X1  g1178(.A1(new_n1374), .A2(new_n1378), .A3(new_n1375), .ZN(new_n1379));
  AND3_X1   g1179(.A1(new_n1377), .A2(new_n1366), .A3(new_n1379), .ZN(new_n1380));
  AOI21_X1  g1180(.A(new_n1366), .B1(new_n1377), .B2(new_n1379), .ZN(new_n1381));
  OAI21_X1  g1181(.A(new_n1360), .B1(new_n1380), .B2(new_n1381), .ZN(new_n1382));
  NAND2_X1  g1182(.A1(new_n1377), .A2(new_n1379), .ZN(new_n1383));
  NAND2_X1  g1183(.A1(new_n1383), .A2(new_n1335), .ZN(new_n1384));
  NAND3_X1  g1184(.A1(new_n1377), .A2(new_n1366), .A3(new_n1379), .ZN(new_n1385));
  INV_X1    g1185(.A(new_n1360), .ZN(new_n1386));
  NAND3_X1  g1186(.A1(new_n1384), .A2(new_n1385), .A3(new_n1386), .ZN(new_n1387));
  NAND2_X1  g1187(.A1(new_n1382), .A2(new_n1387), .ZN(G402));
endmodule


